module real_aes_5668_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_537;
wire n_320;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_298;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_960;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_397;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_140;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
NAND2xp5_ASAP7_75t_L g135 ( .A(n_0), .B(n_136), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_1), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_SL g211 ( .A1(n_2), .A2(n_158), .B(n_212), .C(n_214), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g148 ( .A1(n_3), .A2(n_83), .B1(n_143), .B2(n_149), .Y(n_148) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_4), .A2(n_32), .B1(n_598), .B2(n_599), .Y(n_597) );
OAI22xp5_ASAP7_75t_SL g521 ( .A1(n_5), .A2(n_59), .B1(n_522), .B2(n_523), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_5), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_6), .B(n_526), .Y(n_525) );
INVxp67_ASAP7_75t_L g115 ( .A(n_7), .Y(n_115) );
INVx1_ASAP7_75t_L g545 ( .A(n_7), .Y(n_545) );
INVx1_ASAP7_75t_L g938 ( .A(n_7), .Y(n_938) );
BUFx2_ASAP7_75t_L g957 ( .A(n_7), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_8), .A2(n_91), .B1(n_666), .B2(n_667), .Y(n_665) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_9), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_10), .A2(n_69), .B1(n_149), .B2(n_203), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_11), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_12), .A2(n_33), .B1(n_567), .B2(n_581), .Y(n_580) );
XOR2x2_ASAP7_75t_L g122 ( .A(n_13), .B(n_75), .Y(n_122) );
INVx2_ASAP7_75t_L g640 ( .A(n_13), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_14), .A2(n_61), .B1(n_143), .B2(n_164), .Y(n_201) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_15), .A2(n_68), .B(n_139), .Y(n_138) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_15), .A2(n_68), .B(n_139), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_16), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g638 ( .A(n_17), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_18), .B(n_167), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_19), .Y(n_182) );
BUFx3_ASAP7_75t_L g109 ( .A(n_20), .Y(n_109) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_21), .A2(n_150), .B(n_219), .C(n_220), .Y(n_218) );
OAI22xp33_ASAP7_75t_SL g142 ( .A1(n_22), .A2(n_47), .B1(n_143), .B2(n_144), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_23), .A2(n_31), .B1(n_144), .B2(n_189), .Y(n_264) );
O2A1O1Ixp5_ASAP7_75t_L g687 ( .A1(n_24), .A2(n_584), .B(n_688), .C(n_691), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_25), .B(n_562), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g945 ( .A(n_26), .Y(n_945) );
O2A1O1Ixp5_ASAP7_75t_L g301 ( .A1(n_27), .A2(n_158), .B(n_302), .C(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g120 ( .A(n_28), .Y(n_120) );
INVx1_ASAP7_75t_SL g696 ( .A(n_29), .Y(n_696) );
OAI21xp33_ASAP7_75t_SL g180 ( .A1(n_30), .A2(n_143), .B(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g958 ( .A(n_34), .B(n_959), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_35), .B(n_228), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_36), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_37), .A2(n_41), .B1(n_602), .B2(n_603), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_38), .A2(n_67), .B1(n_603), .B2(n_616), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_39), .B(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g624 ( .A(n_40), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_42), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_43), .B(n_325), .Y(n_672) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_44), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_45), .A2(n_150), .B(n_636), .C(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g658 ( .A(n_46), .Y(n_658) );
INVx2_ASAP7_75t_L g697 ( .A(n_48), .Y(n_697) );
INVx1_ASAP7_75t_L g139 ( .A(n_49), .Y(n_139) );
AND2x4_ASAP7_75t_L g152 ( .A(n_50), .B(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g176 ( .A(n_50), .B(n_153), .Y(n_176) );
INVx2_ASAP7_75t_L g617 ( .A(n_51), .Y(n_617) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_52), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_53), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_54), .A2(n_158), .B(n_186), .C(n_188), .Y(n_185) );
INVx2_ASAP7_75t_L g238 ( .A(n_55), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_56), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_57), .Y(n_160) );
INVx1_ASAP7_75t_SL g692 ( .A(n_58), .Y(n_692) );
INVx1_ASAP7_75t_L g523 ( .A(n_59), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_60), .B(n_167), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_62), .A2(n_79), .B1(n_213), .B2(n_266), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_63), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_64), .A2(n_105), .B1(n_949), .B2(n_960), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_65), .Y(n_165) );
NAND2xp33_ASAP7_75t_R g206 ( .A(n_66), .B(n_178), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_66), .A2(n_103), .B1(n_228), .B2(n_276), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_70), .A2(n_535), .B1(n_536), .B2(n_539), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_70), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_71), .A2(n_150), .B(n_598), .C(n_620), .Y(n_619) );
OR2x6_ASAP7_75t_L g117 ( .A(n_72), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g955 ( .A(n_72), .Y(n_955) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_73), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g644 ( .A(n_74), .Y(n_644) );
INVx1_ASAP7_75t_L g654 ( .A(n_76), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_77), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_78), .B(n_567), .Y(n_566) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_80), .B(n_302), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_81), .A2(n_158), .B(n_613), .C(n_615), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g734 ( .A1(n_81), .A2(n_158), .B(n_613), .C(n_615), .Y(n_734) );
INVx1_ASAP7_75t_L g119 ( .A(n_82), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_82), .B(n_120), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_84), .A2(n_95), .B1(n_586), .B2(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g959 ( .A(n_85), .Y(n_959) );
BUFx5_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_86), .Y(n_145) );
INVx1_ASAP7_75t_L g190 ( .A(n_86), .Y(n_190) );
INVx2_ASAP7_75t_L g225 ( .A(n_87), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_88), .B(n_649), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_89), .A2(n_102), .B1(n_537), .B2(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_89), .Y(n_537) );
INVx2_ASAP7_75t_L g193 ( .A(n_90), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_92), .Y(n_221) );
INVx2_ASAP7_75t_SL g153 ( .A(n_93), .Y(n_153) );
INVx1_ASAP7_75t_L g308 ( .A(n_94), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_96), .B(n_178), .Y(n_655) );
INVx1_ASAP7_75t_SL g607 ( .A(n_97), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_98), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g312 ( .A(n_99), .Y(n_312) );
AND2x2_ASAP7_75t_L g590 ( .A(n_100), .B(n_251), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_101), .A2(n_532), .B1(n_533), .B2(n_534), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_101), .Y(n_532) );
INVx1_ASAP7_75t_L g538 ( .A(n_102), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_103), .B(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_SL g254 ( .A(n_103), .Y(n_254) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_110), .B(n_528), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_109), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_121), .B(n_525), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
BUFx8_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx12f_ASAP7_75t_L g527 ( .A(n_113), .Y(n_527) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OR2x6_ASAP7_75t_L g937 ( .A(n_116), .B(n_938), .Y(n_937) );
INVx8_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g544 ( .A(n_117), .B(n_545), .Y(n_544) );
OR2x6_ASAP7_75t_L g947 ( .A(n_117), .B(n_545), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
XOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
AOI22x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_521), .B2(n_524), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g546 ( .A(n_125), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_125), .A2(n_548), .B1(n_937), .B2(n_941), .Y(n_940) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_435), .Y(n_125) );
NAND4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_332), .C(n_387), .D(n_416), .Y(n_126) );
NOR2xp67_ASAP7_75t_L g127 ( .A(n_128), .B(n_241), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_194), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI221xp5_ASAP7_75t_SL g333 ( .A1(n_130), .A2(n_334), .B1(n_340), .B2(n_342), .C(n_345), .Y(n_333) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_169), .Y(n_130) );
INVx1_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g417 ( .A(n_132), .B(n_418), .Y(n_417) );
OAI21xp33_ASAP7_75t_L g517 ( .A1(n_132), .A2(n_518), .B(n_520), .Y(n_517) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_154), .Y(n_132) );
AND2x2_ASAP7_75t_L g319 ( .A(n_133), .B(n_173), .Y(n_319) );
INVx1_ASAP7_75t_L g412 ( .A(n_133), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_133), .B(n_297), .Y(n_454) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_134), .Y(n_280) );
INVx2_ASAP7_75t_L g291 ( .A(n_134), .Y(n_291) );
NAND2xp33_ASAP7_75t_R g350 ( .A(n_134), .B(n_173), .Y(n_350) );
INVx1_ASAP7_75t_L g373 ( .A(n_134), .Y(n_373) );
AND2x2_ASAP7_75t_L g380 ( .A(n_134), .B(n_154), .Y(n_380) );
AND2x2_ASAP7_75t_L g392 ( .A(n_134), .B(n_173), .Y(n_392) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
INVx2_ASAP7_75t_L g156 ( .A(n_136), .Y(n_156) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_136), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_137), .B(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_137), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g228 ( .A(n_137), .Y(n_228) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
BUFx3_ASAP7_75t_L g325 ( .A(n_138), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_147), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_142), .B(n_146), .Y(n_141) );
AOI22xp33_ASAP7_75t_SL g159 ( .A1(n_143), .A2(n_144), .B1(n_160), .B2(n_161), .Y(n_159) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_143), .A2(n_163), .B1(n_164), .B2(n_165), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_143), .B(n_182), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_143), .A2(n_144), .B1(n_233), .B2(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_143), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_143), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g562 ( .A(n_143), .Y(n_562) );
INVx2_ASAP7_75t_L g567 ( .A(n_143), .Y(n_567) );
INVx2_ASAP7_75t_L g588 ( .A(n_143), .Y(n_588) );
INVx1_ASAP7_75t_L g614 ( .A(n_143), .Y(n_614) );
NAND2xp33_ASAP7_75t_L g631 ( .A(n_143), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g666 ( .A(n_143), .Y(n_666) );
INVx2_ASAP7_75t_L g215 ( .A(n_144), .Y(n_215) );
INVx2_ASAP7_75t_SL g266 ( .A(n_144), .Y(n_266) );
INVx1_ASAP7_75t_L g565 ( .A(n_144), .Y(n_565) );
INVx1_ASAP7_75t_L g647 ( .A(n_144), .Y(n_647) );
INVx2_ASAP7_75t_L g690 ( .A(n_144), .Y(n_690) );
INVx6_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g149 ( .A(n_145), .Y(n_149) );
INVx2_ASAP7_75t_L g164 ( .A(n_145), .Y(n_164) );
INVx3_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx3_ASAP7_75t_L g150 ( .A(n_146), .Y(n_150) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_146), .Y(n_158) );
INVx4_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_146), .Y(n_263) );
INVx1_ASAP7_75t_L g267 ( .A(n_146), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_146), .B(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_L g669 ( .A(n_146), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_150), .B(n_151), .Y(n_147) );
INVx2_ASAP7_75t_L g616 ( .A(n_149), .Y(n_616) );
INVx1_ASAP7_75t_L g649 ( .A(n_149), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g157 ( .A1(n_150), .A2(n_152), .B1(n_158), .B2(n_159), .C(n_162), .Y(n_157) );
INVx3_ASAP7_75t_L g582 ( .A(n_150), .Y(n_582) );
INVx1_ASAP7_75t_L g205 ( .A(n_152), .Y(n_205) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_152), .Y(n_249) );
INVx3_ASAP7_75t_L g570 ( .A(n_152), .Y(n_570) );
AND2x2_ASAP7_75t_L g589 ( .A(n_152), .B(n_324), .Y(n_589) );
AND2x2_ASAP7_75t_L g258 ( .A(n_154), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g321 ( .A(n_154), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g360 ( .A(n_154), .B(n_361), .Y(n_360) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_166), .Y(n_154) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_155), .A2(n_157), .B(n_166), .Y(n_283) );
NOR2x1_ASAP7_75t_SL g628 ( .A(n_155), .B(n_223), .Y(n_628) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OR2x2_ASAP7_75t_L g253 ( .A(n_156), .B(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_158), .A2(n_184), .B1(n_201), .B2(n_202), .Y(n_200) );
INVx1_ASAP7_75t_L g239 ( .A(n_158), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g252 ( .A1(n_158), .A2(n_184), .B1(n_232), .B2(n_236), .Y(n_252) );
INVx1_ASAP7_75t_L g568 ( .A(n_158), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_158), .B(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_158), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_SL g671 ( .A(n_158), .Y(n_671) );
INVx1_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_164), .A2(n_189), .B1(n_237), .B2(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g581 ( .A(n_164), .Y(n_581) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_164), .Y(n_636) );
NOR2xp67_ASAP7_75t_L g204 ( .A(n_167), .B(n_205), .Y(n_204) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_168), .B(n_193), .Y(n_192) );
BUFx3_ASAP7_75t_L g240 ( .A(n_168), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_168), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g414 ( .A(n_169), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_170), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_170), .B(n_341), .Y(n_424) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g270 ( .A(n_172), .Y(n_270) );
AND2x2_ASAP7_75t_L g495 ( .A(n_172), .B(n_380), .Y(n_495) );
AND2x2_ASAP7_75t_L g518 ( .A(n_172), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g284 ( .A(n_173), .Y(n_284) );
INVx2_ASAP7_75t_L g297 ( .A(n_173), .Y(n_297) );
OR2x2_ASAP7_75t_L g385 ( .A(n_173), .B(n_291), .Y(n_385) );
AND2x2_ASAP7_75t_L g432 ( .A(n_173), .B(n_282), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_173), .B(n_283), .Y(n_450) );
BUFx2_ASAP7_75t_L g482 ( .A(n_173), .Y(n_482) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI21x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_179), .B(n_192), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
INVx4_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_176), .B(n_250), .Y(n_261) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx3_ASAP7_75t_L g251 ( .A(n_178), .Y(n_251) );
INVx2_ASAP7_75t_L g277 ( .A(n_178), .Y(n_277) );
INVx1_ASAP7_75t_L g313 ( .A(n_178), .Y(n_313) );
INVx1_ASAP7_75t_L g556 ( .A(n_178), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_183), .B(n_185), .Y(n_179) );
AOI221xp5_ASAP7_75t_L g230 ( .A1(n_183), .A2(n_223), .B1(n_231), .B2(n_235), .C(n_239), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_183), .A2(n_559), .B(n_561), .Y(n_558) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_184), .A2(n_306), .B1(n_307), .B2(n_309), .Y(n_305) );
O2A1O1Ixp5_ASAP7_75t_SL g643 ( .A1(n_184), .A2(n_644), .B(n_645), .C(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g302 ( .A(n_187), .Y(n_302) );
INVx1_ASAP7_75t_L g306 ( .A(n_187), .Y(n_306) );
INVx2_ASAP7_75t_L g560 ( .A(n_187), .Y(n_560) );
INVx2_ASAP7_75t_L g667 ( .A(n_187), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_189), .B(n_191), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_189), .B(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g587 ( .A(n_189), .Y(n_587) );
INVx2_ASAP7_75t_L g603 ( .A(n_189), .Y(n_603) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g203 ( .A(n_190), .Y(n_203) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_194), .A2(n_417), .B1(n_419), .B2(n_422), .C(n_425), .Y(n_416) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_207), .Y(n_195) );
OR2x2_ASAP7_75t_L g244 ( .A(n_196), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_196), .B(n_246), .Y(n_444) );
OR2x2_ASAP7_75t_L g477 ( .A(n_196), .B(n_352), .Y(n_477) );
INVx2_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g288 ( .A(n_198), .B(n_247), .Y(n_288) );
INVx2_ASAP7_75t_L g339 ( .A(n_198), .Y(n_339) );
AND2x2_ASAP7_75t_L g383 ( .A(n_198), .B(n_344), .Y(n_383) );
INVx1_ASAP7_75t_L g397 ( .A(n_198), .Y(n_397) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_206), .Y(n_198) );
AND2x2_ASAP7_75t_L g274 ( .A(n_199), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_204), .Y(n_199) );
INVx2_ASAP7_75t_L g213 ( .A(n_203), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_205), .B(n_325), .Y(n_698) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_207), .Y(n_440) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g434 ( .A(n_208), .B(n_338), .Y(n_434) );
AND2x2_ASAP7_75t_L g507 ( .A(n_208), .B(n_396), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_208), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_226), .Y(n_208) );
AND2x4_ASAP7_75t_L g246 ( .A(n_209), .B(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g287 ( .A(n_209), .Y(n_287) );
INVx1_ASAP7_75t_L g337 ( .A(n_209), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_209), .B(n_299), .Y(n_348) );
INVx2_ASAP7_75t_L g354 ( .A(n_209), .Y(n_354) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_209), .Y(n_400) );
OR2x2_ASAP7_75t_L g421 ( .A(n_209), .B(n_226), .Y(n_421) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_209), .Y(n_515) );
AO31x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_217), .A3(n_222), .B(n_224), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g598 ( .A(n_213), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_215), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_219), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_223), .B(n_301), .C(n_305), .Y(n_300) );
NOR4xp25_ASAP7_75t_L g733 ( .A(n_223), .B(n_619), .C(n_700), .D(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g315 ( .A(n_226), .B(n_287), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_226), .B(n_298), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_226), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
INVx2_ASAP7_75t_L g605 ( .A(n_228), .Y(n_605) );
AND2x2_ASAP7_75t_L g273 ( .A(n_229), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_230), .B(n_240), .Y(n_229) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_240), .A2(n_300), .B(n_311), .Y(n_299) );
INVx2_ASAP7_75t_L g660 ( .A(n_240), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_293), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_255), .B(n_271), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OAI21xp33_ASAP7_75t_L g401 ( .A1(n_246), .A2(n_402), .B(n_404), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_246), .B(n_396), .Y(n_404) );
AND2x2_ASAP7_75t_L g496 ( .A(n_246), .B(n_338), .Y(n_496) );
AND2x2_ASAP7_75t_L g520 ( .A(n_246), .B(n_383), .Y(n_520) );
INVx1_ASAP7_75t_L g328 ( .A(n_247), .Y(n_328) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_252), .B(n_253), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_249), .B(n_324), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_249), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_269), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_258), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_258), .B(n_368), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_258), .A2(n_384), .B(n_430), .Y(n_471) );
INVx1_ASAP7_75t_L g361 ( .A(n_259), .Y(n_361) );
INVx3_ASAP7_75t_L g379 ( .A(n_259), .Y(n_379) );
AND2x2_ASAP7_75t_L g519 ( .A(n_259), .B(n_291), .Y(n_519) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g375 ( .A(n_260), .Y(n_375) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_268), .Y(n_260) );
INVx1_ASAP7_75t_L g323 ( .A(n_262), .Y(n_323) );
OA22x2_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B1(n_265), .B2(n_267), .Y(n_262) );
INVx4_ASAP7_75t_L g584 ( .A(n_263), .Y(n_584) );
INVx1_ASAP7_75t_L g326 ( .A(n_268), .Y(n_326) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_270), .B(n_417), .Y(n_499) );
OAI22x1_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_278), .B1(n_285), .B2(n_289), .Y(n_271) );
OR2x2_ASAP7_75t_L g342 ( .A(n_272), .B(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g409 ( .A(n_272), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g464 ( .A(n_272), .B(n_348), .Y(n_464) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g386 ( .A(n_273), .B(n_344), .Y(n_386) );
INVx1_ASAP7_75t_L g514 ( .A(n_273), .Y(n_514) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_277), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g700 ( .A(n_277), .Y(n_700) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_280), .B(n_375), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g292 ( .A(n_283), .Y(n_292) );
INVx1_ASAP7_75t_L g358 ( .A(n_284), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g458 ( .A1(n_285), .A2(n_389), .B1(n_404), .B2(n_459), .C(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x4_ASAP7_75t_L g346 ( .A(n_288), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g370 ( .A(n_288), .B(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g390 ( .A(n_290), .B(n_374), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_290), .B(n_482), .Y(n_505) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x4_ASAP7_75t_L g393 ( .A(n_292), .B(n_322), .Y(n_393) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_314), .B(n_316), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
BUFx2_ASAP7_75t_L g368 ( .A(n_297), .Y(n_368) );
AND2x4_ASAP7_75t_L g338 ( .A(n_298), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_299), .Y(n_331) );
INVx2_ASAP7_75t_L g344 ( .A(n_299), .Y(n_344) );
AND2x2_ASAP7_75t_L g371 ( .A(n_299), .B(n_354), .Y(n_371) );
AND2x2_ASAP7_75t_L g396 ( .A(n_299), .B(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_R g511 ( .A(n_299), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_315), .B(n_396), .Y(n_426) );
NAND4xp75_ASAP7_75t_L g316 ( .A(n_317), .B(n_320), .C(n_327), .D(n_329), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g340 ( .A(n_318), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_319), .B(n_379), .Y(n_460) );
OAI32xp33_ASAP7_75t_L g408 ( .A1(n_320), .A2(n_409), .A3(n_411), .B1(n_413), .B2(n_414), .Y(n_408) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g341 ( .A(n_321), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B(n_326), .Y(n_322) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND3x1_ASAP7_75t_L g456 ( .A(n_330), .B(n_439), .C(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_362), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g490 ( .A(n_337), .Y(n_490) );
AND2x2_ASAP7_75t_L g438 ( .A(n_338), .B(n_358), .Y(n_438) );
AND2x2_ASAP7_75t_L g365 ( .A(n_339), .B(n_354), .Y(n_365) );
INVx1_ASAP7_75t_L g493 ( .A(n_339), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_341), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g446 ( .A(n_341), .B(n_412), .Y(n_446) );
AND2x2_ASAP7_75t_L g488 ( .A(n_341), .B(n_384), .Y(n_488) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g470 ( .A(n_344), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_349), .B1(n_351), .B2(n_356), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g413 ( .A(n_351), .Y(n_413) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g366 ( .A(n_355), .Y(n_366) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g406 ( .A(n_358), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_358), .B(n_359), .Y(n_466) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_359), .Y(n_462) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g457 ( .A(n_360), .B(n_368), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g479 ( .A(n_360), .B(n_475), .C(n_480), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_369), .B2(n_372), .C(n_376), .Y(n_362) );
INVxp67_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x2_ASAP7_75t_L g468 ( .A(n_365), .B(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_369), .A2(n_466), .B1(n_467), .B2(n_471), .Y(n_465) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g410 ( .A(n_371), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g431 ( .A(n_373), .Y(n_431) );
NOR2xp67_ASAP7_75t_L g449 ( .A(n_373), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_374), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_384), .B2(n_386), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx3_ASAP7_75t_L g418 ( .A(n_379), .Y(n_418) );
AND2x2_ASAP7_75t_L g502 ( .A(n_379), .B(n_495), .Y(n_502) );
AND2x2_ASAP7_75t_L g516 ( .A(n_379), .B(n_392), .Y(n_516) );
AND2x2_ASAP7_75t_L g428 ( .A(n_380), .B(n_418), .Y(n_428) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OR2x2_ASAP7_75t_L g484 ( .A(n_382), .B(n_395), .Y(n_484) );
BUFx2_ASAP7_75t_L g403 ( .A(n_383), .Y(n_403) );
AND2x2_ASAP7_75t_L g486 ( .A(n_384), .B(n_393), .Y(n_486) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_394), .B1(n_401), .B2(n_405), .C(n_408), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx2_ASAP7_75t_L g407 ( .A(n_393), .Y(n_407) );
INVx2_ASAP7_75t_SL g476 ( .A(n_393), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_398), .Y(n_394) );
OR2x2_ASAP7_75t_L g451 ( .A(n_395), .B(n_398), .Y(n_451) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g419 ( .A(n_396), .B(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_413), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g437 ( .A(n_418), .B(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_418), .B(n_481), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_419), .A2(n_434), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_429), .B2(n_433), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g435 ( .A(n_436), .B(n_455), .C(n_472), .D(n_497), .Y(n_435) );
AOI221x1_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_441), .B2(n_445), .C(n_447), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .B(n_452), .Y(n_447) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_458), .C(n_465), .Y(n_455) );
BUFx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI21xp33_ASAP7_75t_SL g473 ( .A1(n_467), .A2(n_474), .B(n_477), .Y(n_473) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_469), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_470), .B(n_493), .Y(n_492) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_478), .B(n_483), .Y(n_472) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_487), .B2(n_489), .C(n_494), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
O2A1O1Ixp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_500), .B(n_503), .C(n_504), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI211xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_508), .C(n_517), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_512), .B(n_516), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g524 ( .A(n_521), .Y(n_524) );
INVx1_ASAP7_75t_L g943 ( .A(n_525), .Y(n_943) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_939), .B(n_948), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_540), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI211xp5_ASAP7_75t_L g939 ( .A1(n_531), .A2(n_940), .B(n_943), .C(n_944), .Y(n_939) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2x1p5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_547), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx8_ASAP7_75t_L g942 ( .A(n_544), .Y(n_942) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_548), .B(n_933), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_549), .B(n_814), .Y(n_548) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_748), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_710), .Y(n_550) );
OAI21xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_572), .B(n_673), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g926 ( .A(n_552), .B(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g725 ( .A(n_554), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g809 ( .A(n_554), .B(n_642), .Y(n_809) );
AND2x2_ASAP7_75t_L g834 ( .A(n_554), .B(n_806), .Y(n_834) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_557), .B(n_571), .Y(n_554) );
OA21x2_ASAP7_75t_L g662 ( .A1(n_555), .A2(n_663), .B(n_672), .Y(n_662) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_556), .B(n_624), .Y(n_623) );
OAI21x1_ASAP7_75t_L g681 ( .A1(n_557), .A2(n_571), .B(n_660), .Y(n_681) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_563), .B(n_569), .Y(n_557) );
INVx1_ASAP7_75t_L g599 ( .A(n_560), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_562), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B(n_568), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_568), .A2(n_630), .B(n_633), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_569), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI21x1_ASAP7_75t_L g659 ( .A1(n_570), .A2(n_655), .B(n_660), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_625), .C(n_661), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g879 ( .A1(n_573), .A2(n_757), .B1(n_880), .B2(n_882), .C1(n_884), .C2(n_887), .Y(n_879) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_591), .Y(n_574) );
OR2x2_ASAP7_75t_L g836 ( .A(n_575), .B(n_837), .Y(n_836) );
AND2x2_ASAP7_75t_L g844 ( .A(n_575), .B(n_774), .Y(n_844) );
BUFx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_576), .B(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g731 ( .A(n_576), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g751 ( .A(n_576), .B(n_608), .Y(n_751) );
INVx1_ASAP7_75t_L g855 ( .A(n_576), .Y(n_855) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2x1_ASAP7_75t_L g708 ( .A(n_577), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g738 ( .A(n_578), .Y(n_738) );
AO31x2_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_583), .A3(n_589), .B(n_590), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_582), .A2(n_601), .B(n_604), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_584), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g652 ( .A(n_588), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g817 ( .A1(n_591), .A2(n_818), .B1(n_819), .B2(n_821), .C(n_825), .Y(n_817) );
NOR2x1_ASAP7_75t_L g832 ( .A(n_591), .B(n_833), .Y(n_832) );
OR2x2_ASAP7_75t_L g881 ( .A(n_591), .B(n_716), .Y(n_881) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2x1p5_ASAP7_75t_L g846 ( .A(n_592), .B(n_707), .Y(n_846) );
AND2x4_ASAP7_75t_L g592 ( .A(n_593), .B(n_608), .Y(n_592) );
OR2x2_ASAP7_75t_L g730 ( .A(n_593), .B(n_718), .Y(n_730) );
AND2x2_ASAP7_75t_L g812 ( .A(n_593), .B(n_662), .Y(n_812) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g766 ( .A(n_594), .Y(n_766) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g709 ( .A(n_595), .Y(n_709) );
AOI21x1_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_600), .B(n_606), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_598), .B(n_692), .Y(n_691) );
AOI21x1_ASAP7_75t_L g718 ( .A1(n_605), .A2(n_719), .B(n_720), .Y(n_718) );
NOR2x1_ASAP7_75t_L g721 ( .A(n_608), .B(n_709), .Y(n_721) );
OA21x2_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_622), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_618), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_616), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g695 ( .A(n_616), .Y(n_695) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVxp67_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g732 ( .A(n_623), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_625), .B(n_712), .Y(n_711) );
OAI32xp33_ASAP7_75t_L g792 ( .A1(n_625), .A2(n_793), .A3(n_794), .B1(n_796), .B2(n_799), .Y(n_792) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g676 ( .A(n_626), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g779 ( .A(n_626), .B(n_780), .Y(n_779) );
NOR2xp67_ASAP7_75t_L g841 ( .A(n_626), .B(n_793), .Y(n_841) );
AND2x2_ASAP7_75t_L g864 ( .A(n_626), .B(n_797), .Y(n_864) );
AND2x2_ASAP7_75t_L g893 ( .A(n_626), .B(n_824), .Y(n_893) );
AND2x4_ASAP7_75t_L g626 ( .A(n_627), .B(n_641), .Y(n_626) );
OR2x2_ASAP7_75t_L g701 ( .A(n_627), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g723 ( .A(n_627), .Y(n_723) );
AND2x2_ASAP7_75t_L g757 ( .A(n_627), .B(n_702), .Y(n_757) );
INVx2_ASAP7_75t_L g788 ( .A(n_627), .Y(n_788) );
OR2x2_ASAP7_75t_L g798 ( .A(n_627), .B(n_641), .Y(n_798) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_627), .Y(n_872) );
AO31x2_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .A3(n_634), .B(n_639), .Y(n_627) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g753 ( .A(n_641), .B(n_685), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_641), .B(n_679), .Y(n_919) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g772 ( .A(n_642), .B(n_680), .Y(n_772) );
OAI21x1_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_650), .B(n_659), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_643), .A2(n_650), .B(n_659), .Y(n_702) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_646), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND3x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_655), .C(n_656), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
OAI32xp33_ASAP7_75t_L g755 ( .A1(n_661), .A2(n_756), .A3(n_757), .B1(n_758), .B2(n_759), .Y(n_755) );
INVx1_ASAP7_75t_L g833 ( .A(n_661), .Y(n_833) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_662), .Y(n_707) );
INVx1_ASAP7_75t_L g740 ( .A(n_662), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_662), .B(n_738), .Y(n_763) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_664), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B1(n_670), .B2(n_671), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_668), .A2(n_694), .B(n_698), .Y(n_693) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g720 ( .A(n_672), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_703), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_682), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_675), .A2(n_758), .B1(n_782), .B2(n_785), .Y(n_781) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NAND2x1p5_ASAP7_75t_L g818 ( .A(n_678), .B(n_753), .Y(n_818) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_SL g747 ( .A(n_679), .Y(n_747) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_679), .Y(n_754) );
AND2x2_ASAP7_75t_L g807 ( .A(n_679), .B(n_788), .Y(n_807) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g684 ( .A(n_680), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g824 ( .A(n_680), .B(n_806), .Y(n_824) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_701), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
BUFx2_ASAP7_75t_L g712 ( .A(n_684), .Y(n_712) );
NAND2x1_ASAP7_75t_SL g883 ( .A(n_684), .B(n_872), .Y(n_883) );
INVx2_ASAP7_75t_SL g744 ( .A(n_685), .Y(n_744) );
BUFx2_ASAP7_75t_L g790 ( .A(n_685), .Y(n_790) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g726 ( .A(n_686), .Y(n_726) );
INVx1_ASAP7_75t_L g761 ( .A(n_686), .Y(n_761) );
OA21x2_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_693), .B(n_699), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g856 ( .A(n_701), .B(n_857), .Y(n_856) );
NAND3xp33_ASAP7_75t_L g860 ( .A(n_701), .B(n_756), .C(n_861), .Y(n_860) );
OR2x2_ASAP7_75t_L g909 ( .A(n_701), .B(n_769), .Y(n_909) );
INVx1_ASAP7_75t_L g921 ( .A(n_701), .Y(n_921) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_702), .Y(n_822) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_704), .A2(n_850), .B1(n_854), .B2(n_856), .Y(n_849) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g904 ( .A(n_705), .B(n_867), .Y(n_904) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g866 ( .A(n_706), .B(n_867), .Y(n_866) );
NOR2x1p5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx2_ASAP7_75t_L g802 ( .A(n_707), .Y(n_802) );
INVx2_ASAP7_75t_L g915 ( .A(n_707), .Y(n_915) );
OR2x2_ASAP7_75t_L g888 ( .A(n_708), .B(n_889), .Y(n_888) );
AND2x2_ASAP7_75t_L g774 ( .A(n_709), .B(n_718), .Y(n_774) );
INVx1_ASAP7_75t_L g830 ( .A(n_709), .Y(n_830) );
OAI222xp33_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_713), .B1(n_722), .B2(n_727), .C1(n_735), .C2(n_741), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_721), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g898 ( .A(n_717), .B(n_766), .Y(n_898) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_721), .B(n_737), .Y(n_784) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx2_ASAP7_75t_SL g746 ( .A(n_723), .Y(n_746) );
AND2x4_ASAP7_75t_L g827 ( .A(n_723), .B(n_809), .Y(n_827) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g793 ( .A(n_725), .Y(n_793) );
INVx2_ASAP7_75t_L g806 ( .A(n_726), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_726), .B(n_853), .Y(n_852) );
O2A1O1Ixp33_ASAP7_75t_L g905 ( .A1(n_727), .A2(n_906), .B(n_908), .C(n_909), .Y(n_905) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
AND2x4_ASAP7_75t_L g750 ( .A(n_729), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g854 ( .A(n_730), .B(n_855), .Y(n_854) );
AND2x4_ASAP7_75t_L g773 ( .A(n_731), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_731), .B(n_778), .Y(n_777) );
INVx2_ASAP7_75t_SL g813 ( .A(n_731), .Y(n_813) );
AND2x2_ASAP7_75t_L g900 ( .A(n_731), .B(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g907 ( .A(n_731), .Y(n_907) );
NOR2x1_ASAP7_75t_L g739 ( .A(n_732), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_732), .B(n_765), .Y(n_764) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_732), .Y(n_795) );
INVx1_ASAP7_75t_L g800 ( .A(n_732), .Y(n_800) );
INVx1_ASAP7_75t_L g876 ( .A(n_732), .Y(n_876) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_735), .B(n_777), .Y(n_776) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_735), .A2(n_767), .B1(n_836), .B2(n_838), .Y(n_835) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g859 ( .A(n_736), .B(n_830), .Y(n_859) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_737), .B(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g896 ( .A(n_737), .Y(n_896) );
BUFx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g889 ( .A(n_739), .Y(n_889) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g769 ( .A(n_744), .Y(n_769) );
AND2x2_ASAP7_75t_L g771 ( .A(n_744), .B(n_772), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_744), .B(n_874), .Y(n_873) );
OR2x6_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g780 ( .A(n_747), .Y(n_780) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_775), .C(n_791), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B1(n_755), .B2(n_767), .C(n_770), .Y(n_749) );
INVx1_ASAP7_75t_L g758 ( .A(n_751), .Y(n_758) );
AND2x2_ASAP7_75t_L g820 ( .A(n_751), .B(n_774), .Y(n_820) );
AND2x2_ASAP7_75t_L g828 ( .A(n_751), .B(n_829), .Y(n_828) );
AND2x2_ASAP7_75t_L g914 ( .A(n_751), .B(n_915), .Y(n_914) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g768 ( .A(n_757), .B(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
BUFx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_R g797 ( .A(n_761), .Y(n_797) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx1_ASAP7_75t_L g923 ( .A(n_763), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_764), .Y(n_924) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g778 ( .A(n_766), .Y(n_778) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_766), .Y(n_901) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
AND2x2_ASAP7_75t_L g871 ( .A(n_771), .B(n_872), .Y(n_871) );
INVx2_ASAP7_75t_L g839 ( .A(n_772), .Y(n_839) );
AND2x2_ASAP7_75t_L g903 ( .A(n_772), .B(n_788), .Y(n_903) );
AND2x2_ASAP7_75t_L g789 ( .A(n_774), .B(n_790), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_779), .B(n_781), .Y(n_775) );
OAI221xp5_ASAP7_75t_L g911 ( .A1(n_782), .A2(n_912), .B1(n_913), .B2(n_916), .C(n_920), .Y(n_911) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g932 ( .A(n_784), .Y(n_932) );
NAND2x1_ASAP7_75t_L g785 ( .A(n_786), .B(n_789), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
OR2x2_ASAP7_75t_L g838 ( .A(n_788), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g853 ( .A(n_788), .Y(n_853) );
INVx1_ASAP7_75t_L g885 ( .A(n_790), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_801), .B(n_803), .Y(n_791) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI222xp33_ASAP7_75t_L g891 ( .A1(n_796), .A2(n_892), .B1(n_894), .B2(n_899), .C1(n_902), .C2(n_904), .Y(n_891) );
OR2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
AND2x2_ASAP7_75t_L g826 ( .A(n_797), .B(n_809), .Y(n_826) );
AND2x2_ASAP7_75t_L g917 ( .A(n_797), .B(n_918), .Y(n_917) );
INVx2_ASAP7_75t_L g886 ( .A(n_798), .Y(n_886) );
INVx1_ASAP7_75t_L g930 ( .A(n_798), .Y(n_930) );
INVx1_ASAP7_75t_L g867 ( .A(n_800), .Y(n_867) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g878 ( .A(n_802), .Y(n_878) );
AOI21xp33_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_808), .B(n_810), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
OR2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g837 ( .A(n_812), .Y(n_837) );
INVx1_ASAP7_75t_L g908 ( .A(n_812), .Y(n_908) );
NOR2x1p5_ASAP7_75t_L g814 ( .A(n_815), .B(n_868), .Y(n_814) );
NAND3xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_840), .C(n_858), .Y(n_815) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_831), .C(n_835), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g928 ( .A1(n_818), .A2(n_848), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
AO22x1_ASAP7_75t_L g831 ( .A1(n_820), .A2(n_826), .B1(n_832), .B2(n_834), .Y(n_831) );
OR2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
INVxp67_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g848 ( .A(n_824), .Y(n_848) );
INVx1_ASAP7_75t_L g857 ( .A(n_824), .Y(n_857) );
OAI21xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_827), .B(n_828), .Y(n_825) );
INVx2_ASAP7_75t_L g874 ( .A(n_827), .Y(n_874) );
INVxp67_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g865 ( .A(n_834), .Y(n_865) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_839), .B(n_852), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_845), .B2(n_847), .C(n_849), .Y(n_840) );
INVxp67_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx2_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_852), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B1(n_862), .B2(n_866), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_863), .B(n_865), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NAND4xp75_ASAP7_75t_L g868 ( .A(n_869), .B(n_890), .C(n_910), .D(n_925), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_870), .B(n_879), .Y(n_869) );
OAI21xp33_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_873), .B(n_875), .Y(n_870) );
INVx1_ASAP7_75t_L g927 ( .A(n_872), .Y(n_927) );
NOR2xp33_ASAP7_75t_SL g875 ( .A(n_876), .B(n_877), .Y(n_875) );
AND2x4_ASAP7_75t_L g931 ( .A(n_877), .B(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_SL g882 ( .A(n_883), .Y(n_882) );
BUFx2_ASAP7_75t_L g912 ( .A(n_883), .Y(n_912) );
AND2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NOR2x1_ASAP7_75t_L g890 ( .A(n_891), .B(n_905), .Y(n_890) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
OR2x2_ASAP7_75t_L g894 ( .A(n_895), .B(n_897), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
AND2x2_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
OAI21xp5_ASAP7_75t_L g925 ( .A1(n_926), .A2(n_928), .B(n_931), .Y(n_925) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
BUFx12f_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
CKINVDCx11_ASAP7_75t_R g935 ( .A(n_936), .Y(n_935) );
INVx2_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx2_ASAP7_75t_SL g941 ( .A(n_942), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
BUFx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
BUFx2_ASAP7_75t_SL g949 ( .A(n_950), .Y(n_949) );
BUFx8_ASAP7_75t_L g961 ( .A(n_950), .Y(n_961) );
AND2x4_ASAP7_75t_L g950 ( .A(n_951), .B(n_953), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
NAND3xp33_ASAP7_75t_L g954 ( .A(n_955), .B(n_956), .C(n_958), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_957), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_961), .Y(n_960) );
endmodule