module fake_jpeg_25541_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_19),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_59),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_52),
.B1(n_67),
.B2(n_55),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_80),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_67),
.B1(n_52),
.B2(n_68),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_58),
.B1(n_66),
.B2(n_64),
.Y(n_87)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_95),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_99),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_65),
.B1(n_61),
.B2(n_50),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_97),
.B1(n_62),
.B2(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_46),
.B1(n_56),
.B2(n_57),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx11_ASAP7_75t_SL g114 ( 
.A(n_100),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_102),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_60),
.C(n_68),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_106),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_62),
.C(n_49),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_1),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_100),
.B(n_45),
.CI(n_2),
.CON(n_112),
.SN(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_54),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_123),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_91),
.B1(n_88),
.B2(n_96),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_120),
.B1(n_125),
.B2(n_104),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_45),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_6),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_88),
.B1(n_48),
.B2(n_54),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_3),
.B(n_5),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_5),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_140)
);

AOI21x1_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_112),
.B(n_105),
.Y(n_127)
);

AOI221xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_133),
.B1(n_137),
.B2(n_8),
.C(n_10),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_130),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_115),
.B(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_138),
.B(n_7),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_24),
.B1(n_43),
.B2(n_42),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_28),
.B1(n_41),
.B2(n_13),
.Y(n_145)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_135),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_6),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_140),
.B(n_143),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_134),
.C(n_12),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_131),
.B1(n_130),
.B2(n_138),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_149),
.B(n_139),
.C(n_146),
.Y(n_150)
);

OAI21x1_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_143),
.B(n_148),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_141),
.C(n_142),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_145),
.B(n_29),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_25),
.B(n_40),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_22),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_21),
.B(n_35),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_15),
.C(n_18),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);


endmodule