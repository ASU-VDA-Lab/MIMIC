module real_aes_8848_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_769;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_756;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_0), .Y(n_460) );
INVx1_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
INVx1_ASAP7_75t_L g488 ( .A(n_2), .Y(n_488) );
INVx1_ASAP7_75t_L g199 ( .A(n_3), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_4), .A2(n_39), .B1(n_160), .B2(n_518), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_5), .A2(n_102), .B1(n_114), .B2(n_777), .Y(n_101) );
AOI21xp33_ASAP7_75t_L g167 ( .A1(n_6), .A2(n_141), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_7), .B(n_134), .Y(n_501) );
AND2x6_ASAP7_75t_L g146 ( .A(n_8), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_9), .A2(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_10), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_10), .B(n_40), .Y(n_457) );
INVx1_ASAP7_75t_L g174 ( .A(n_11), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_12), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g139 ( .A(n_13), .Y(n_139) );
INVx1_ASAP7_75t_L g482 ( .A(n_14), .Y(n_482) );
INVx1_ASAP7_75t_L g255 ( .A(n_15), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_16), .B(n_182), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_17), .B(n_135), .Y(n_559) );
AO32x2_ASAP7_75t_L g531 ( .A1(n_18), .A2(n_134), .A3(n_179), .B1(n_510), .B2(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_19), .A2(n_63), .B1(n_123), .B2(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_19), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_20), .B(n_160), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_21), .B(n_155), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_22), .B(n_135), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_23), .A2(n_51), .B1(n_160), .B2(n_518), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_24), .B(n_141), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_25), .A2(n_77), .B1(n_160), .B2(n_182), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_26), .B(n_160), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_27), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_28), .A2(n_253), .B(n_254), .C(n_256), .Y(n_252) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_29), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_30), .B(n_176), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_31), .B(n_172), .Y(n_201) );
INVx1_ASAP7_75t_L g188 ( .A(n_32), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_33), .B(n_176), .Y(n_548) );
INVx2_ASAP7_75t_L g144 ( .A(n_34), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_35), .B(n_160), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_36), .B(n_176), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_37), .Y(n_774) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_38), .A2(n_146), .B(n_150), .C(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
INVx1_ASAP7_75t_L g186 ( .A(n_41), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_42), .B(n_172), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_43), .B(n_160), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_44), .A2(n_87), .B1(n_218), .B2(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_45), .B(n_160), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_46), .B(n_160), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_47), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_48), .A2(n_70), .B1(n_762), .B2(n_763), .Y(n_761) );
CKINVDCx16_ASAP7_75t_R g763 ( .A(n_48), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_49), .B(n_487), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_50), .B(n_141), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_52), .A2(n_61), .B1(n_160), .B2(n_182), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_53), .A2(n_150), .B1(n_182), .B2(n_184), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_54), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_55), .B(n_160), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_56), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_57), .B(n_160), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_58), .A2(n_159), .B(n_171), .C(n_173), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_59), .Y(n_231) );
INVx1_ASAP7_75t_L g169 ( .A(n_60), .Y(n_169) );
INVx1_ASAP7_75t_L g147 ( .A(n_62), .Y(n_147) );
INVx1_ASAP7_75t_L g123 ( .A(n_63), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_64), .B(n_160), .Y(n_489) );
INVx1_ASAP7_75t_L g138 ( .A(n_65), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
AO32x2_ASAP7_75t_L g515 ( .A1(n_67), .A2(n_134), .A3(n_235), .B1(n_510), .B2(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g508 ( .A(n_68), .Y(n_508) );
INVx1_ASAP7_75t_L g543 ( .A(n_69), .Y(n_543) );
INVx1_ASAP7_75t_L g762 ( .A(n_70), .Y(n_762) );
A2O1A1Ixp33_ASAP7_75t_SL g154 ( .A1(n_71), .A2(n_155), .B(n_156), .C(n_159), .Y(n_154) );
INVxp67_ASAP7_75t_L g157 ( .A(n_72), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_73), .B(n_182), .Y(n_544) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_75), .Y(n_192) );
INVx1_ASAP7_75t_L g224 ( .A(n_76), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_78), .A2(n_146), .B(n_150), .C(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_79), .B(n_518), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_80), .B(n_182), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_81), .B(n_200), .Y(n_214) );
INVx2_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_83), .B(n_155), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_84), .B(n_182), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_85), .A2(n_146), .B(n_150), .C(n_198), .Y(n_197) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_86), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g454 ( .A(n_86), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g465 ( .A(n_86), .B(n_456), .Y(n_465) );
INVx2_ASAP7_75t_L g469 ( .A(n_86), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_88), .A2(n_100), .B1(n_182), .B2(n_183), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_89), .B(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_90), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_91), .A2(n_146), .B(n_150), .C(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_92), .Y(n_245) );
INVx1_ASAP7_75t_L g153 ( .A(n_93), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_94), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_95), .B(n_200), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_96), .B(n_182), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_97), .B(n_134), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_99), .A2(n_141), .B(n_148), .Y(n_140) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_SL g779 ( .A(n_104), .Y(n_779) );
AND2x2_ASAP7_75t_SL g104 ( .A(n_105), .B(n_111), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g456 ( .A(n_107), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_461), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g776 ( .A(n_117), .Y(n_776) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_451), .B(n_458), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_125), .B2(n_450), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g450 ( .A(n_125), .Y(n_450) );
INVx1_ASAP7_75t_SL g466 ( .A(n_125), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_125), .A2(n_765), .B1(n_767), .B2(n_768), .Y(n_764) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND4x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_368), .C(n_415), .D(n_435), .Y(n_126) );
NOR3xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_298), .C(n_323), .Y(n_127) );
OAI211xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_206), .B(n_258), .C(n_288), .Y(n_128) );
INVxp67_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_177), .Y(n_130) );
INVx3_ASAP7_75t_SL g340 ( .A(n_131), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_131), .B(n_271), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_131), .B(n_193), .Y(n_421) );
AND2x2_ASAP7_75t_L g444 ( .A(n_131), .B(n_310), .Y(n_444) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_165), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g262 ( .A(n_133), .B(n_166), .Y(n_262) );
INVx3_ASAP7_75t_L g275 ( .A(n_133), .Y(n_275) );
AND2x2_ASAP7_75t_L g280 ( .A(n_133), .B(n_165), .Y(n_280) );
OR2x2_ASAP7_75t_L g331 ( .A(n_133), .B(n_272), .Y(n_331) );
BUFx2_ASAP7_75t_L g351 ( .A(n_133), .Y(n_351) );
AND2x2_ASAP7_75t_L g361 ( .A(n_133), .B(n_272), .Y(n_361) );
AND2x2_ASAP7_75t_L g367 ( .A(n_133), .B(n_178), .Y(n_367) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_162), .Y(n_133) );
INVx4_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_134), .A2(n_494), .B(n_501), .Y(n_493) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_136), .B(n_137), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx2_ASAP7_75t_L g249 ( .A(n_141), .Y(n_249) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_142), .B(n_146), .Y(n_190) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g487 ( .A(n_143), .Y(n_487) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
INVx1_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
INVx1_ASAP7_75t_L g152 ( .A(n_145), .Y(n_152) );
INVx1_ASAP7_75t_L g155 ( .A(n_145), .Y(n_155) );
INVx3_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_145), .Y(n_185) );
INVx4_ASAP7_75t_SL g161 ( .A(n_146), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_146), .A2(n_481), .B(n_485), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_146), .A2(n_495), .B(n_498), .Y(n_494) );
BUFx3_ASAP7_75t_L g510 ( .A(n_146), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_146), .A2(n_523), .B(n_527), .Y(n_522) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_146), .A2(n_542), .B(n_545), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_153), .B(n_154), .C(n_161), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_149), .A2(n_161), .B(n_169), .C(n_170), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_149), .A2(n_161), .B(n_251), .C(n_252), .Y(n_250) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
BUFx3_ASAP7_75t_L g218 ( .A(n_151), .Y(n_218) );
INVx1_ASAP7_75t_L g518 ( .A(n_151), .Y(n_518) );
INVx1_ASAP7_75t_L g526 ( .A(n_155), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_158), .B(n_174), .Y(n_173) );
INVx5_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g516 ( .A1(n_158), .A2(n_172), .B1(n_517), .B2(n_519), .Y(n_516) );
O2A1O1Ixp5_ASAP7_75t_SL g542 ( .A1(n_159), .A2(n_200), .B(n_543), .C(n_544), .Y(n_542) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_160), .Y(n_242) );
OAI22xp33_ASAP7_75t_L g180 ( .A1(n_161), .A2(n_181), .B1(n_189), .B2(n_190), .Y(n_180) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_163), .A2(n_167), .B(n_175), .Y(n_166) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_SL g220 ( .A(n_164), .B(n_221), .Y(n_220) );
AO21x1_ASAP7_75t_L g554 ( .A1(n_164), .A2(n_555), .B(n_558), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_164), .B(n_510), .C(n_555), .Y(n_573) );
INVx1_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_166), .B(n_272), .Y(n_286) );
INVx2_ASAP7_75t_L g296 ( .A(n_166), .Y(n_296) );
AND2x2_ASAP7_75t_L g309 ( .A(n_166), .B(n_275), .Y(n_309) );
OR2x2_ASAP7_75t_L g320 ( .A(n_166), .B(n_272), .Y(n_320) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_166), .B(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g378 ( .A(n_166), .Y(n_378) );
AND2x2_ASAP7_75t_L g424 ( .A(n_166), .B(n_178), .Y(n_424) );
O2A1O1Ixp5_ASAP7_75t_L g507 ( .A1(n_171), .A2(n_486), .B(n_508), .C(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_171), .A2(n_528), .B(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g241 ( .A(n_172), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_172), .A2(n_490), .B1(n_533), .B2(n_534), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_172), .A2(n_490), .B1(n_556), .B2(n_557), .Y(n_555) );
INVx1_ASAP7_75t_L g205 ( .A(n_176), .Y(n_205) );
INVx2_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_176), .A2(n_248), .B(n_257), .Y(n_247) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_176), .A2(n_522), .B(n_530), .Y(n_521) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_176), .A2(n_541), .B(n_548), .Y(n_540) );
INVx3_ASAP7_75t_SL g297 ( .A(n_177), .Y(n_297) );
OR2x2_ASAP7_75t_L g350 ( .A(n_177), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
INVx3_ASAP7_75t_L g272 ( .A(n_178), .Y(n_272) );
AND2x2_ASAP7_75t_L g339 ( .A(n_178), .B(n_194), .Y(n_339) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_178), .Y(n_407) );
AOI33xp33_ASAP7_75t_L g411 ( .A1(n_178), .A2(n_340), .A3(n_347), .B1(n_356), .B2(n_412), .B3(n_413), .Y(n_411) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_191), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_179), .B(n_192), .Y(n_191) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_179), .A2(n_195), .B(n_203), .Y(n_194) );
INVx2_ASAP7_75t_L g219 ( .A(n_179), .Y(n_219) );
INVx2_ASAP7_75t_L g202 ( .A(n_182), .Y(n_202) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g184 ( .A1(n_185), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_184) );
INVx2_ASAP7_75t_L g187 ( .A(n_185), .Y(n_187) );
INVx4_ASAP7_75t_L g253 ( .A(n_185), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_190), .A2(n_196), .B(n_197), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_190), .A2(n_224), .B(n_225), .Y(n_223) );
INVx1_ASAP7_75t_L g260 ( .A(n_193), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_193), .B(n_275), .Y(n_274) );
NOR3xp33_ASAP7_75t_L g334 ( .A(n_193), .B(n_335), .C(n_337), .Y(n_334) );
AND2x2_ASAP7_75t_L g360 ( .A(n_193), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_193), .B(n_367), .Y(n_370) );
AND2x2_ASAP7_75t_L g423 ( .A(n_193), .B(n_424), .Y(n_423) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g279 ( .A(n_194), .Y(n_279) );
OR2x2_ASAP7_75t_L g373 ( .A(n_194), .B(n_272), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .C(n_202), .Y(n_198) );
INVx2_ASAP7_75t_L g490 ( .A(n_200), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_200), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_200), .A2(n_505), .B(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_202), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_205), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_205), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_232), .Y(n_206) );
AOI32xp33_ASAP7_75t_L g324 ( .A1(n_207), .A2(n_325), .A3(n_327), .B1(n_329), .B2(n_332), .Y(n_324) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_207), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g427 ( .A(n_207), .Y(n_427) );
INVx4_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g359 ( .A(n_208), .B(n_343), .Y(n_359) );
AND2x2_ASAP7_75t_L g379 ( .A(n_208), .B(n_305), .Y(n_379) );
AND2x2_ASAP7_75t_L g447 ( .A(n_208), .B(n_365), .Y(n_447) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_222), .Y(n_208) );
INVx3_ASAP7_75t_L g268 ( .A(n_209), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_209), .B(n_266), .Y(n_282) );
OR2x2_ASAP7_75t_L g287 ( .A(n_209), .B(n_265), .Y(n_287) );
INVx1_ASAP7_75t_L g294 ( .A(n_209), .Y(n_294) );
AND2x2_ASAP7_75t_L g302 ( .A(n_209), .B(n_276), .Y(n_302) );
AND2x2_ASAP7_75t_L g304 ( .A(n_209), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_209), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g357 ( .A(n_209), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_209), .B(n_442), .Y(n_441) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_220), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_212), .B(n_219), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_216), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g256 ( .A(n_218), .Y(n_256) );
INVx1_ASAP7_75t_L g229 ( .A(n_219), .Y(n_229) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_219), .A2(n_480), .B(n_491), .Y(n_479) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_219), .A2(n_503), .B(n_511), .Y(n_502) );
INVx2_ASAP7_75t_L g266 ( .A(n_222), .Y(n_266) );
AND2x2_ASAP7_75t_L g312 ( .A(n_222), .B(n_233), .Y(n_312) );
AND2x2_ASAP7_75t_L g322 ( .A(n_222), .B(n_247), .Y(n_322) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_230), .Y(n_222) );
INVx2_ASAP7_75t_L g442 ( .A(n_232), .Y(n_442) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_246), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_233), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g283 ( .A(n_233), .Y(n_283) );
AND2x2_ASAP7_75t_L g327 ( .A(n_233), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g343 ( .A(n_233), .B(n_306), .Y(n_343) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g291 ( .A(n_234), .Y(n_291) );
AND2x2_ASAP7_75t_L g305 ( .A(n_234), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g356 ( .A(n_234), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_234), .B(n_266), .Y(n_388) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_244), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_242), .Y(n_238) );
AND2x2_ASAP7_75t_L g267 ( .A(n_246), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g328 ( .A(n_246), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_246), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g365 ( .A(n_246), .Y(n_365) );
INVx1_ASAP7_75t_L g398 ( .A(n_246), .Y(n_398) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g276 ( .A(n_247), .B(n_266), .Y(n_276) );
INVx1_ASAP7_75t_L g306 ( .A(n_247), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_253), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g484 ( .A(n_253), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_253), .A2(n_546), .B(n_547), .Y(n_545) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_263), .B1(n_269), .B2(n_276), .C(n_277), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_260), .B(n_280), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_260), .B(n_343), .Y(n_420) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_262), .B(n_310), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_262), .B(n_271), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_262), .B(n_285), .Y(n_414) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g336 ( .A(n_266), .Y(n_336) );
AND2x2_ASAP7_75t_L g311 ( .A(n_267), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g389 ( .A(n_267), .Y(n_389) );
AND2x2_ASAP7_75t_L g321 ( .A(n_268), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_268), .B(n_291), .Y(n_337) );
AND2x2_ASAP7_75t_L g401 ( .A(n_268), .B(n_327), .Y(n_401) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g310 ( .A(n_272), .B(n_279), .Y(n_310) );
AND2x2_ASAP7_75t_L g406 ( .A(n_273), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_275), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_276), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_276), .B(n_283), .Y(n_371) );
AND2x2_ASAP7_75t_L g391 ( .A(n_276), .B(n_291), .Y(n_391) );
AND2x2_ASAP7_75t_L g412 ( .A(n_276), .B(n_356), .Y(n_412) );
OAI32xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .A3(n_283), .B1(n_284), .B2(n_287), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_SL g285 ( .A(n_279), .Y(n_285) );
NAND2x1_ASAP7_75t_L g326 ( .A(n_279), .B(n_309), .Y(n_326) );
OR2x2_ASAP7_75t_L g330 ( .A(n_279), .B(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_279), .B(n_378), .Y(n_431) );
INVx1_ASAP7_75t_L g299 ( .A(n_280), .Y(n_299) );
OAI221xp5_ASAP7_75t_SL g417 ( .A1(n_281), .A2(n_372), .B1(n_418), .B2(n_421), .C(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g289 ( .A(n_282), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g332 ( .A(n_282), .B(n_305), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_282), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g410 ( .A(n_282), .B(n_343), .Y(n_410) );
INVxp67_ASAP7_75t_L g346 ( .A(n_283), .Y(n_346) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g416 ( .A(n_285), .B(n_403), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_285), .B(n_366), .Y(n_439) );
INVx1_ASAP7_75t_L g314 ( .A(n_287), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_287), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g432 ( .A(n_287), .B(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_292), .B(n_295), .Y(n_288) );
AND2x2_ASAP7_75t_L g301 ( .A(n_290), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g385 ( .A(n_294), .B(n_305), .Y(n_385) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x2_ASAP7_75t_L g403 ( .A(n_296), .B(n_361), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_296), .B(n_360), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_297), .B(n_309), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_303), .C(n_313), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g333 ( .A1(n_299), .A2(n_334), .B1(n_338), .B2(n_341), .C(n_344), .Y(n_333) );
AOI31xp33_ASAP7_75t_L g428 ( .A1(n_299), .A2(n_429), .A3(n_430), .B(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .B1(n_309), .B2(n_311), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g429 ( .A(n_309), .Y(n_429) );
INVx1_ASAP7_75t_L g392 ( .A(n_310), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g435 ( .A1(n_312), .A2(n_436), .B(n_438), .C(n_440), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_317), .B2(n_321), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_318), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_320), .A2(n_354), .B1(n_373), .B2(n_409), .C(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g404 ( .A(n_321), .Y(n_404) );
INVx1_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
NAND3xp33_ASAP7_75t_SL g323 ( .A(n_324), .B(n_333), .C(n_348), .Y(n_323) );
OAI21xp33_ASAP7_75t_L g374 ( .A1(n_325), .A2(n_375), .B(n_379), .Y(n_374) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_327), .B(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g434 ( .A(n_328), .Y(n_434) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g372 ( .A(n_335), .B(n_355), .Y(n_372) );
INVx1_ASAP7_75t_L g347 ( .A(n_336), .Y(n_347) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g345 ( .A(n_339), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_339), .B(n_377), .Y(n_376) );
NOR4xp25_ASAP7_75t_L g344 ( .A(n_340), .B(n_345), .C(n_346), .D(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI222xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B1(n_359), .B2(n_360), .C1(n_362), .C2(n_366), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_350), .B(n_352), .Y(n_349) );
INVx1_ASAP7_75t_L g446 ( .A(n_350), .Y(n_446) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_362), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_367), .A2(n_423), .B(n_425), .Y(n_422) );
NOR4xp25_ASAP7_75t_L g368 ( .A(n_369), .B(n_380), .C(n_393), .D(n_408), .Y(n_368) );
OAI221xp5_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_371), .B1(n_372), .B2(n_373), .C(n_374), .Y(n_369) );
INVx1_ASAP7_75t_L g449 ( .A(n_370), .Y(n_449) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_377), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
OAI222xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B1(n_386), .B2(n_387), .C1(n_390), .C2(n_392), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI211xp5_ASAP7_75t_L g415 ( .A1(n_385), .A2(n_416), .B(n_417), .C(n_428), .Y(n_415) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
OAI222xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_399), .B1(n_400), .B2(n_402), .C1(n_404), .C2(n_405), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_410), .A2(n_413), .B1(n_446), .B2(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_443), .B(n_445), .C(n_448), .Y(n_440) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g459 ( .A(n_454), .Y(n_459) );
NOR2x2_ASAP7_75t_L g773 ( .A(n_455), .B(n_469), .Y(n_773) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g468 ( .A(n_456), .B(n_469), .Y(n_468) );
OAI21xp5_ASAP7_75t_SL g461 ( .A1(n_458), .A2(n_462), .B(n_775), .Y(n_461) );
NOR2xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_460), .Y(n_458) );
OAI222xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_761), .B1(n_764), .B2(n_769), .C1(n_770), .C2(n_774), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_466), .B1(n_467), .B2(n_470), .Y(n_463) );
INVx2_ASAP7_75t_L g766 ( .A(n_464), .Y(n_766) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx6_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g767 ( .A(n_468), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_470), .Y(n_768) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_471), .B(n_727), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_631), .C(n_715), .Y(n_471) );
NAND4xp25_ASAP7_75t_L g472 ( .A(n_473), .B(n_574), .C(n_596), .D(n_612), .Y(n_472) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_512), .B1(n_535), .B2(n_553), .C(n_560), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_492), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_476), .B(n_553), .Y(n_586) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_476), .B(n_614), .C(n_627), .D(n_629), .Y(n_626) );
INVxp67_ASAP7_75t_L g743 ( .A(n_476), .Y(n_743) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g625 ( .A(n_477), .B(n_563), .Y(n_625) );
AND2x2_ASAP7_75t_L g649 ( .A(n_477), .B(n_492), .Y(n_649) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g616 ( .A(n_478), .B(n_552), .Y(n_616) );
AND2x2_ASAP7_75t_L g656 ( .A(n_478), .B(n_637), .Y(n_656) );
AND2x2_ASAP7_75t_L g673 ( .A(n_478), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_478), .B(n_493), .Y(n_697) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g551 ( .A(n_479), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g568 ( .A(n_479), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g580 ( .A(n_479), .B(n_493), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_479), .B(n_502), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_488), .B(n_489), .C(n_490), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_490), .A2(n_499), .B(n_500), .Y(n_498) );
AND2x2_ASAP7_75t_L g583 ( .A(n_492), .B(n_584), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_492), .A2(n_633), .B1(n_636), .B2(n_638), .C(n_642), .Y(n_632) );
AND2x2_ASAP7_75t_L g691 ( .A(n_492), .B(n_656), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_492), .B(n_673), .Y(n_725) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
INVx3_ASAP7_75t_L g552 ( .A(n_493), .Y(n_552) );
AND2x2_ASAP7_75t_L g600 ( .A(n_493), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g654 ( .A(n_493), .B(n_569), .Y(n_654) );
AND2x2_ASAP7_75t_L g712 ( .A(n_493), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g553 ( .A(n_502), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g569 ( .A(n_502), .Y(n_569) );
INVx1_ASAP7_75t_L g624 ( .A(n_502), .Y(n_624) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_502), .Y(n_630) );
AND2x2_ASAP7_75t_L g675 ( .A(n_502), .B(n_552), .Y(n_675) );
OR2x2_ASAP7_75t_L g714 ( .A(n_502), .B(n_554), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_507), .B(n_510), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_512), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
AND2x2_ASAP7_75t_L g710 ( .A(n_513), .B(n_707), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_513), .B(n_692), .Y(n_742) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g641 ( .A(n_514), .B(n_565), .Y(n_641) );
AND2x2_ASAP7_75t_L g690 ( .A(n_514), .B(n_538), .Y(n_690) );
INVx1_ASAP7_75t_L g736 ( .A(n_514), .Y(n_736) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_515), .Y(n_550) );
AND2x2_ASAP7_75t_L g591 ( .A(n_515), .B(n_565), .Y(n_591) );
INVx1_ASAP7_75t_L g608 ( .A(n_515), .Y(n_608) );
AND2x2_ASAP7_75t_L g614 ( .A(n_515), .B(n_531), .Y(n_614) );
AND2x2_ASAP7_75t_L g682 ( .A(n_520), .B(n_590), .Y(n_682) );
INVx2_ASAP7_75t_L g747 ( .A(n_520), .Y(n_747) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_531), .Y(n_520) );
AND2x2_ASAP7_75t_L g564 ( .A(n_521), .B(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g577 ( .A(n_521), .B(n_539), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_521), .B(n_538), .Y(n_605) );
INVx1_ASAP7_75t_L g611 ( .A(n_521), .Y(n_611) );
INVx1_ASAP7_75t_L g628 ( .A(n_521), .Y(n_628) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_521), .Y(n_640) );
INVx2_ASAP7_75t_L g708 ( .A(n_521), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_526), .Y(n_523) );
INVx2_ASAP7_75t_L g565 ( .A(n_531), .Y(n_565) );
BUFx2_ASAP7_75t_L g662 ( .A(n_531), .Y(n_662) );
AND2x2_ASAP7_75t_L g707 ( .A(n_531), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_549), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_537), .B(n_644), .Y(n_643) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_537), .A2(n_706), .B(n_720), .Y(n_730) );
AND2x2_ASAP7_75t_L g755 ( .A(n_537), .B(n_641), .Y(n_755) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g677 ( .A(n_539), .Y(n_677) );
AND2x2_ASAP7_75t_L g706 ( .A(n_539), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_540), .Y(n_590) );
INVx2_ASAP7_75t_L g609 ( .A(n_540), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_540), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx2_ASAP7_75t_L g563 ( .A(n_550), .Y(n_563) );
OR2x2_ASAP7_75t_L g576 ( .A(n_550), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g644 ( .A(n_550), .B(n_640), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_550), .B(n_740), .Y(n_739) );
OR2x2_ASAP7_75t_L g745 ( .A(n_550), .B(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_550), .B(n_682), .Y(n_757) );
AND2x2_ASAP7_75t_L g636 ( .A(n_551), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g659 ( .A(n_551), .B(n_553), .Y(n_659) );
INVx2_ASAP7_75t_L g571 ( .A(n_552), .Y(n_571) );
AND2x2_ASAP7_75t_L g599 ( .A(n_552), .B(n_572), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_552), .B(n_624), .Y(n_680) );
AND2x2_ASAP7_75t_L g594 ( .A(n_553), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g741 ( .A(n_553), .Y(n_741) );
AND2x2_ASAP7_75t_L g753 ( .A(n_553), .B(n_616), .Y(n_753) );
AND2x2_ASAP7_75t_L g579 ( .A(n_554), .B(n_569), .Y(n_579) );
INVx1_ASAP7_75t_L g674 ( .A(n_554), .Y(n_674) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g572 ( .A(n_559), .B(n_573), .Y(n_572) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_566), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_563), .B(n_610), .Y(n_619) );
OR2x2_ASAP7_75t_L g751 ( .A(n_563), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g668 ( .A(n_564), .B(n_609), .Y(n_668) );
AND2x2_ASAP7_75t_L g676 ( .A(n_564), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g735 ( .A(n_564), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g759 ( .A(n_564), .B(n_606), .Y(n_759) );
NOR2xp67_ASAP7_75t_L g717 ( .A(n_565), .B(n_718), .Y(n_717) );
OR2x2_ASAP7_75t_L g746 ( .A(n_565), .B(n_609), .Y(n_746) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2x1p5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
AND2x2_ASAP7_75t_L g598 ( .A(n_568), .B(n_599), .Y(n_598) );
INVxp67_ASAP7_75t_L g760 ( .A(n_568), .Y(n_760) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g595 ( .A(n_571), .Y(n_595) );
AND2x2_ASAP7_75t_L g646 ( .A(n_571), .B(n_579), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_571), .B(n_714), .Y(n_740) );
INVx2_ASAP7_75t_L g585 ( .A(n_572), .Y(n_585) );
INVx3_ASAP7_75t_L g637 ( .A(n_572), .Y(n_637) );
OR2x2_ASAP7_75t_L g665 ( .A(n_572), .B(n_666), .Y(n_665) );
AOI311xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_578), .A3(n_580), .B(n_581), .C(n_592), .Y(n_574) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_575), .A2(n_613), .B(n_615), .C(n_617), .Y(n_612) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_SL g597 ( .A(n_577), .Y(n_597) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g615 ( .A(n_579), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_579), .B(n_595), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_579), .B(n_580), .Y(n_748) );
AND2x2_ASAP7_75t_L g670 ( .A(n_580), .B(n_584), .Y(n_670) );
AOI21xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_586), .B(n_587), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g728 ( .A(n_584), .B(n_616), .Y(n_728) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_585), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g622 ( .A(n_585), .Y(n_622) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
AND2x2_ASAP7_75t_L g613 ( .A(n_589), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g658 ( .A(n_591), .Y(n_658) );
AND2x4_ASAP7_75t_L g720 ( .A(n_591), .B(n_689), .Y(n_720) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_594), .A2(n_660), .B1(n_672), .B2(n_676), .C1(n_678), .C2(n_682), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_600), .C(n_603), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_597), .B(n_641), .Y(n_664) );
INVx1_ASAP7_75t_L g686 ( .A(n_599), .Y(n_686) );
INVx1_ASAP7_75t_L g620 ( .A(n_601), .Y(n_620) );
OR2x2_ASAP7_75t_L g685 ( .A(n_602), .B(n_686), .Y(n_685) );
OAI21xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_606), .B(n_610), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_604), .B(n_622), .C(n_623), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_604), .A2(n_641), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_608), .Y(n_661) );
AND2x2_ASAP7_75t_SL g627 ( .A(n_609), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g718 ( .A(n_609), .Y(n_718) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_609), .Y(n_734) );
INVx2_ASAP7_75t_L g692 ( .A(n_610), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_614), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g666 ( .A(n_616), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B1(n_621), .B2(n_625), .C(n_626), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_620), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g754 ( .A(n_620), .Y(n_754) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g635 ( .A(n_627), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_627), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g693 ( .A(n_627), .B(n_641), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_627), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g726 ( .A(n_627), .B(n_661), .Y(n_726) );
BUFx3_ASAP7_75t_L g689 ( .A(n_628), .Y(n_689) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND5xp2_ASAP7_75t_L g631 ( .A(n_632), .B(n_650), .C(n_671), .D(n_683), .E(n_698), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI32xp33_ASAP7_75t_L g723 ( .A1(n_635), .A2(n_662), .A3(n_678), .B1(n_724), .B2(n_726), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_637), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_SL g647 ( .A(n_641), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_647), .B2(n_648), .Y(n_642) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_657), .B1(n_659), .B2(n_660), .C(n_663), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g722 ( .A(n_654), .B(n_673), .Y(n_722) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_659), .A2(n_720), .B1(n_738), .B2(n_743), .C(n_744), .Y(n_737) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx2_ASAP7_75t_L g703 ( .A(n_662), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_667), .B2(n_669), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g681 ( .A(n_673), .Y(n_681) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_687), .B1(n_691), .B2(n_692), .C1(n_693), .C2(n_694), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_692), .A2(n_739), .B1(n_741), .B2(n_742), .Y(n_738) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B(n_704), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_709), .B(n_711), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g752 ( .A(n_707), .Y(n_752) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_719), .B(n_721), .C(n_723), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI211xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B(n_731), .C(n_756), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_728), .Y(n_732) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI211xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B(n_737), .C(n_749), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
AOI21xp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_747), .B(n_748), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B(n_760), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g769 ( .A(n_761), .Y(n_769) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
endmodule