module fake_jpeg_2102_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_58),
.B(n_61),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_44),
.B1(n_46),
.B2(n_50),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_69),
.B1(n_2),
.B2(n_4),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_56),
.B1(n_45),
.B2(n_41),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_49),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_50),
.B1(n_46),
.B2(n_56),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_45),
.B1(n_52),
.B2(n_54),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_52),
.B1(n_60),
.B2(n_5),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_54),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_2),
.C(n_5),
.Y(n_86)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_78),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_75),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_42),
.B1(n_51),
.B2(n_53),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_84),
.B1(n_89),
.B2(n_74),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_42),
.Y(n_83)
);

INVxp33_ASAP7_75t_SL g104 ( 
.A(n_83),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_72),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_71),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_101),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_103),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_22),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_9),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_25),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_64),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_64),
.C(n_23),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_16),
.C(n_17),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_117),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_97),
.B1(n_13),
.B2(n_10),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_10),
.B(n_11),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_18),
.B(n_19),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_24),
.B1(n_38),
.B2(n_15),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_111),
.B(n_119),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_20),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_129),
.Y(n_141)
);

OAI322xp33_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_134),
.A3(n_32),
.B1(n_33),
.B2(n_36),
.C1(n_39),
.C2(n_117),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_136),
.B1(n_138),
.B2(n_137),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_21),
.B(n_26),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_116),
.B(n_130),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_30),
.C(n_31),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_136),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_108),
.B1(n_122),
.B2(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_142),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_144),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_136),
.C(n_131),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_127),
.B(n_126),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_149),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_141),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_154),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_149),
.C(n_143),
.Y(n_158)
);

AOI211xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_147),
.B(n_145),
.C(n_141),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_132),
.Y(n_160)
);


endmodule