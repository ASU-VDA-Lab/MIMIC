module fake_jpeg_9902_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_2),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_24),
.Y(n_25)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_12),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_9),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_19),
.B1(n_18),
.B2(n_6),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_19),
.B1(n_6),
.B2(n_18),
.Y(n_29)
);

AOI21x1_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_28),
.B(n_9),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_8),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_27),
.C(n_9),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_34),
.B1(n_31),
.B2(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_32),
.C(n_16),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_16),
.C(n_5),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_5),
.B(n_1),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_2),
.Y(n_41)
);


endmodule