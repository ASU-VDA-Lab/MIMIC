module fake_ibex_1650_n_3214 (n_179, n_564, n_120, n_48, n_560, n_40, n_412, n_536, n_325, n_113, n_290, n_215, n_477, n_388, n_221, n_26, n_567, n_178, n_497, n_282, n_55, n_277, n_424, n_541, n_588, n_170, n_555, n_575, n_454, n_367, n_29, n_2, n_320, n_470, n_533, n_593, n_395, n_262, n_181, n_368, n_483, n_161, n_508, n_415, n_24, n_239, n_585, n_1, n_233, n_500, n_311, n_563, n_291, n_371, n_552, n_100, n_220, n_579, n_110, n_496, n_331, n_279, n_125, n_381, n_231, n_154, n_251, n_206, n_460, n_352, n_343, n_590, n_551, n_436, n_64, n_418, n_445, n_348, n_131, n_527, n_540, n_561, n_545, n_19, n_202, n_535, n_237, n_39, n_130, n_63, n_592, n_189, n_38, n_380, n_576, n_15, n_339, n_84, n_183, n_20, n_335, n_518, n_68, n_80, n_507, n_37, n_75, n_107, n_482, n_119, n_133, n_356, n_333, n_472, n_595, n_387, n_91, n_538, n_187, n_307, n_135, n_317, n_305, n_139, n_390, n_481, n_157, n_410, n_491, n_448, n_582, n_57, n_149, n_253, n_550, n_584, n_342, n_532, n_394, n_163, n_162, n_209, n_401, n_502, n_398, n_442, n_116, n_366, n_534, n_543, n_559, n_515, n_386, n_548, n_95, n_200, n_167, n_396, n_322, n_441, n_529, n_361, n_318, n_456, n_79, n_10, n_152, n_88, n_160, n_433, n_229, n_480, n_138, n_417, n_192, n_420, n_272, n_473, n_164, n_403, n_490, n_241, n_414, n_228, n_504, n_190, n_198, n_169, n_310, n_5, n_122, n_344, n_72, n_558, n_224, n_102, n_243, n_400, n_369, n_62, n_421, n_392, n_197, n_232, n_104, n_213, n_428, n_172, n_194, n_76, n_294, n_587, n_438, n_118, n_166, n_432, n_146, n_247, n_376, n_451, n_411, n_523, n_283, n_83, n_499, n_226, n_45, n_405, n_36, n_365, n_528, n_542, n_359, n_260, n_573, n_128, n_115, n_106, n_327, n_245, n_32, n_556, n_150, n_236, n_4, n_81, n_300, n_16, n_458, n_329, n_6, n_147, n_457, n_93, n_121, n_140, n_338, n_332, n_570, n_142, n_429, n_539, n_49, n_252, n_580, n_255, n_234, n_304, n_488, n_303, n_274, n_7, n_475, n_520, n_256, n_312, n_466, n_461, n_308, n_354, n_464, n_134, n_270, n_212, n_180, n_292, n_553, n_375, n_35, n_184, n_562, n_218, n_316, n_498, n_56, n_397, n_101, n_21, n_379, n_281, n_514, n_219, n_50, n_459, n_416, n_42, n_566, n_112, n_156, n_86, n_382, n_47, n_565, n_67, n_357, n_434, n_216, n_82, n_204, n_223, n_298, n_87, n_492, n_171, n_265, n_439, n_103, n_96, n_27, n_33, n_301, n_309, n_513, n_452, n_468, n_22, n_314, n_501, n_254, n_258, n_196, n_340, n_225, n_266, n_74, n_288, n_173, n_185, n_505, n_467, n_315, n_31, n_516, n_422, n_503, n_153, n_177, n_511, n_509, n_512, n_264, n_151, n_443, n_287, n_246, n_453, n_574, n_129, n_132, n_469, n_90, n_364, n_426, n_276, n_127, n_249, n_521, n_519, n_52, n_399, n_547, n_273, n_111, n_319, n_321, n_244, n_524, n_360, n_44, n_94, n_168, n_589, n_60, n_182, n_549, n_280, n_358, n_370, n_78, n_69, n_97, n_261, n_355, n_437, n_571, n_510, n_544, n_284, n_143, n_413, n_51, n_208, n_402, n_449, n_594, n_455, n_423, n_569, n_350, n_341, n_73, n_17, n_210, n_175, n_485, n_92, n_336, n_278, n_230, n_3, n_108, n_440, n_419, n_65, n_85, n_377, n_145, n_478, n_257, n_248, n_61, n_450, n_144, n_53, n_383, n_30, n_238, n_12, n_89, n_54, n_158, n_517, n_546, n_8, n_324, n_299, n_374, n_526, n_578, n_302, n_109, n_525, n_296, n_583, n_59, n_46, n_123, n_11, n_572, n_188, n_347, n_363, n_201, n_462, n_275, n_330, n_444, n_323, n_407, n_117, n_242, n_447, n_34, n_293, n_203, n_522, n_25, n_99, n_227, n_431, n_124, n_425, n_136, n_530, n_554, n_577, n_66, n_28, n_77, n_408, n_176, n_126, n_471, n_465, n_71, n_313, n_148, n_353, n_537, n_385, n_285, n_435, n_141, n_586, n_191, n_207, n_268, n_326, n_155, n_493, n_222, n_41, n_351, n_0, n_476, n_174, n_531, n_235, n_479, n_474, n_557, n_58, n_263, n_486, n_463, n_487, n_214, n_345, n_193, n_391, n_337, n_18, n_211, n_306, n_240, n_205, n_373, n_114, n_267, n_427, n_297, n_409, n_70, n_289, n_195, n_384, n_98, n_259, n_269, n_349, n_159, n_43, n_14, n_165, n_372, n_13, n_430, n_9, n_217, n_484, n_489, n_495, n_137, n_346, n_286, n_378, n_186, n_271, n_199, n_334, n_250, n_446, n_494, n_591, n_506, n_568, n_406, n_105, n_404, n_362, n_23, n_389, n_295, n_581, n_393, n_328, n_3214);

input n_179;
input n_564;
input n_120;
input n_48;
input n_560;
input n_40;
input n_412;
input n_536;
input n_325;
input n_113;
input n_290;
input n_215;
input n_477;
input n_388;
input n_221;
input n_26;
input n_567;
input n_178;
input n_497;
input n_282;
input n_55;
input n_277;
input n_424;
input n_541;
input n_588;
input n_170;
input n_555;
input n_575;
input n_454;
input n_367;
input n_29;
input n_2;
input n_320;
input n_470;
input n_533;
input n_593;
input n_395;
input n_262;
input n_181;
input n_368;
input n_483;
input n_161;
input n_508;
input n_415;
input n_24;
input n_239;
input n_585;
input n_1;
input n_233;
input n_500;
input n_311;
input n_563;
input n_291;
input n_371;
input n_552;
input n_100;
input n_220;
input n_579;
input n_110;
input n_496;
input n_331;
input n_279;
input n_125;
input n_381;
input n_231;
input n_154;
input n_251;
input n_206;
input n_460;
input n_352;
input n_343;
input n_590;
input n_551;
input n_436;
input n_64;
input n_418;
input n_445;
input n_348;
input n_131;
input n_527;
input n_540;
input n_561;
input n_545;
input n_19;
input n_202;
input n_535;
input n_237;
input n_39;
input n_130;
input n_63;
input n_592;
input n_189;
input n_38;
input n_380;
input n_576;
input n_15;
input n_339;
input n_84;
input n_183;
input n_20;
input n_335;
input n_518;
input n_68;
input n_80;
input n_507;
input n_37;
input n_75;
input n_107;
input n_482;
input n_119;
input n_133;
input n_356;
input n_333;
input n_472;
input n_595;
input n_387;
input n_91;
input n_538;
input n_187;
input n_307;
input n_135;
input n_317;
input n_305;
input n_139;
input n_390;
input n_481;
input n_157;
input n_410;
input n_491;
input n_448;
input n_582;
input n_57;
input n_149;
input n_253;
input n_550;
input n_584;
input n_342;
input n_532;
input n_394;
input n_163;
input n_162;
input n_209;
input n_401;
input n_502;
input n_398;
input n_442;
input n_116;
input n_366;
input n_534;
input n_543;
input n_559;
input n_515;
input n_386;
input n_548;
input n_95;
input n_200;
input n_167;
input n_396;
input n_322;
input n_441;
input n_529;
input n_361;
input n_318;
input n_456;
input n_79;
input n_10;
input n_152;
input n_88;
input n_160;
input n_433;
input n_229;
input n_480;
input n_138;
input n_417;
input n_192;
input n_420;
input n_272;
input n_473;
input n_164;
input n_403;
input n_490;
input n_241;
input n_414;
input n_228;
input n_504;
input n_190;
input n_198;
input n_169;
input n_310;
input n_5;
input n_122;
input n_344;
input n_72;
input n_558;
input n_224;
input n_102;
input n_243;
input n_400;
input n_369;
input n_62;
input n_421;
input n_392;
input n_197;
input n_232;
input n_104;
input n_213;
input n_428;
input n_172;
input n_194;
input n_76;
input n_294;
input n_587;
input n_438;
input n_118;
input n_166;
input n_432;
input n_146;
input n_247;
input n_376;
input n_451;
input n_411;
input n_523;
input n_283;
input n_83;
input n_499;
input n_226;
input n_45;
input n_405;
input n_36;
input n_365;
input n_528;
input n_542;
input n_359;
input n_260;
input n_573;
input n_128;
input n_115;
input n_106;
input n_327;
input n_245;
input n_32;
input n_556;
input n_150;
input n_236;
input n_4;
input n_81;
input n_300;
input n_16;
input n_458;
input n_329;
input n_6;
input n_147;
input n_457;
input n_93;
input n_121;
input n_140;
input n_338;
input n_332;
input n_570;
input n_142;
input n_429;
input n_539;
input n_49;
input n_252;
input n_580;
input n_255;
input n_234;
input n_304;
input n_488;
input n_303;
input n_274;
input n_7;
input n_475;
input n_520;
input n_256;
input n_312;
input n_466;
input n_461;
input n_308;
input n_354;
input n_464;
input n_134;
input n_270;
input n_212;
input n_180;
input n_292;
input n_553;
input n_375;
input n_35;
input n_184;
input n_562;
input n_218;
input n_316;
input n_498;
input n_56;
input n_397;
input n_101;
input n_21;
input n_379;
input n_281;
input n_514;
input n_219;
input n_50;
input n_459;
input n_416;
input n_42;
input n_566;
input n_112;
input n_156;
input n_86;
input n_382;
input n_47;
input n_565;
input n_67;
input n_357;
input n_434;
input n_216;
input n_82;
input n_204;
input n_223;
input n_298;
input n_87;
input n_492;
input n_171;
input n_265;
input n_439;
input n_103;
input n_96;
input n_27;
input n_33;
input n_301;
input n_309;
input n_513;
input n_452;
input n_468;
input n_22;
input n_314;
input n_501;
input n_254;
input n_258;
input n_196;
input n_340;
input n_225;
input n_266;
input n_74;
input n_288;
input n_173;
input n_185;
input n_505;
input n_467;
input n_315;
input n_31;
input n_516;
input n_422;
input n_503;
input n_153;
input n_177;
input n_511;
input n_509;
input n_512;
input n_264;
input n_151;
input n_443;
input n_287;
input n_246;
input n_453;
input n_574;
input n_129;
input n_132;
input n_469;
input n_90;
input n_364;
input n_426;
input n_276;
input n_127;
input n_249;
input n_521;
input n_519;
input n_52;
input n_399;
input n_547;
input n_273;
input n_111;
input n_319;
input n_321;
input n_244;
input n_524;
input n_360;
input n_44;
input n_94;
input n_168;
input n_589;
input n_60;
input n_182;
input n_549;
input n_280;
input n_358;
input n_370;
input n_78;
input n_69;
input n_97;
input n_261;
input n_355;
input n_437;
input n_571;
input n_510;
input n_544;
input n_284;
input n_143;
input n_413;
input n_51;
input n_208;
input n_402;
input n_449;
input n_594;
input n_455;
input n_423;
input n_569;
input n_350;
input n_341;
input n_73;
input n_17;
input n_210;
input n_175;
input n_485;
input n_92;
input n_336;
input n_278;
input n_230;
input n_3;
input n_108;
input n_440;
input n_419;
input n_65;
input n_85;
input n_377;
input n_145;
input n_478;
input n_257;
input n_248;
input n_61;
input n_450;
input n_144;
input n_53;
input n_383;
input n_30;
input n_238;
input n_12;
input n_89;
input n_54;
input n_158;
input n_517;
input n_546;
input n_8;
input n_324;
input n_299;
input n_374;
input n_526;
input n_578;
input n_302;
input n_109;
input n_525;
input n_296;
input n_583;
input n_59;
input n_46;
input n_123;
input n_11;
input n_572;
input n_188;
input n_347;
input n_363;
input n_201;
input n_462;
input n_275;
input n_330;
input n_444;
input n_323;
input n_407;
input n_117;
input n_242;
input n_447;
input n_34;
input n_293;
input n_203;
input n_522;
input n_25;
input n_99;
input n_227;
input n_431;
input n_124;
input n_425;
input n_136;
input n_530;
input n_554;
input n_577;
input n_66;
input n_28;
input n_77;
input n_408;
input n_176;
input n_126;
input n_471;
input n_465;
input n_71;
input n_313;
input n_148;
input n_353;
input n_537;
input n_385;
input n_285;
input n_435;
input n_141;
input n_586;
input n_191;
input n_207;
input n_268;
input n_326;
input n_155;
input n_493;
input n_222;
input n_41;
input n_351;
input n_0;
input n_476;
input n_174;
input n_531;
input n_235;
input n_479;
input n_474;
input n_557;
input n_58;
input n_263;
input n_486;
input n_463;
input n_487;
input n_214;
input n_345;
input n_193;
input n_391;
input n_337;
input n_18;
input n_211;
input n_306;
input n_240;
input n_205;
input n_373;
input n_114;
input n_267;
input n_427;
input n_297;
input n_409;
input n_70;
input n_289;
input n_195;
input n_384;
input n_98;
input n_259;
input n_269;
input n_349;
input n_159;
input n_43;
input n_14;
input n_165;
input n_372;
input n_13;
input n_430;
input n_9;
input n_217;
input n_484;
input n_489;
input n_495;
input n_137;
input n_346;
input n_286;
input n_378;
input n_186;
input n_271;
input n_199;
input n_334;
input n_250;
input n_446;
input n_494;
input n_591;
input n_506;
input n_568;
input n_406;
input n_105;
input n_404;
input n_362;
input n_23;
input n_389;
input n_295;
input n_581;
input n_393;
input n_328;

output n_3214;



endmodule