module real_jpeg_27455_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_330, n_12, n_6, n_11, n_14, n_7, n_329, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_330;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_329;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_0),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_48),
.B1(n_49),
.B2(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_63),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_0),
.A2(n_28),
.B1(n_34),
.B2(n_63),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_2),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_153),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_153),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_2),
.A2(n_28),
.B1(n_34),
.B2(n_153),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_3),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_142),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_142),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_3),
.A2(n_28),
.B1(n_34),
.B2(n_142),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_7),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_7),
.A2(n_28),
.B1(n_34),
.B2(n_72),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_72),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_72),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_8),
.A2(n_40),
.B1(n_61),
.B2(n_62),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_8),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_8),
.A2(n_28),
.B1(n_34),
.B2(n_40),
.Y(n_223)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_9),
.A2(n_34),
.A3(n_61),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_85),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_10),
.A2(n_28),
.B1(n_34),
.B2(n_85),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_11),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_11),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_11),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_12),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_103),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_12),
.A2(n_28),
.B1(n_34),
.B2(n_103),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_103),
.Y(n_256)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_14),
.A2(n_48),
.B(n_78),
.C(n_81),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_15),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_15),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_15),
.A2(n_28),
.B1(n_34),
.B2(n_53),
.Y(n_167)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_17),
.A2(n_41),
.B1(n_42),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_17),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_17),
.A2(n_45),
.B(n_49),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_17),
.B(n_47),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_17),
.A2(n_61),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_17),
.B(n_61),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_17),
.B(n_100),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_17),
.A2(n_26),
.B1(n_32),
.B2(n_235),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_17),
.A2(n_48),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_309),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_118),
.A3(n_132),
.B1(n_307),
.B2(n_308),
.C(n_329),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_104),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_21),
.B(n_104),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_90),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_22),
.B(n_75),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_55),
.B1(n_56),
.B2(n_74),
.Y(n_22)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_24),
.A2(n_37),
.B(n_55),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_24),
.A2(n_25),
.B1(n_57),
.B2(n_58),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_25),
.B(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B(n_33),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_26),
.A2(n_30),
.B1(n_33),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_26),
.A2(n_30),
.B1(n_94),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_26),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_26),
.A2(n_30),
.B1(n_229),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_26),
.A2(n_30),
.B1(n_223),
.B2(n_264),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_27),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_27),
.A2(n_31),
.B1(n_158),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_27),
.A2(n_159),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_28),
.A2(n_34),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_28),
.B(n_68),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_28),
.B(n_240),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_30),
.Y(n_159)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_SL g224 ( 
.A(n_31),
.Y(n_224)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_52),
.B2(n_54),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_39),
.A2(n_44),
.B1(n_47),
.B2(n_102),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_41),
.A2(n_51),
.B(n_151),
.C(n_156),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_43),
.A2(n_52),
.B1(n_54),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_43),
.A2(n_54),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_43),
.A2(n_54),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_44),
.A2(n_47),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_44),
.A2(n_47),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_44),
.A2(n_47),
.B1(n_102),
.B2(n_182),
.Y(n_196)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_79),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g260 ( 
.A1(n_48),
.A2(n_62),
.A3(n_79),
.B1(n_253),
.B2(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_49),
.B(n_151),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_70),
.B2(n_73),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_65),
.B1(n_66),
.B2(n_96),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_61),
.B(n_262),
.Y(n_261)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_64),
.A2(n_73),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_64),
.A2(n_73),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_66),
.B1(n_71),
.B2(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_66),
.B(n_88),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_65),
.A2(n_66),
.B1(n_96),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_65),
.A2(n_66),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_65),
.A2(n_66),
.B1(n_209),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_65),
.A2(n_66),
.B1(n_147),
.B2(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_66),
.B(n_151),
.Y(n_236)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_87),
.B(n_89),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_87),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_81),
.B1(n_83),
.B2(n_86),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_77),
.A2(n_81),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_77),
.A2(n_81),
.B1(n_143),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_77),
.A2(n_81),
.B1(n_165),
.B2(n_251),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_77),
.A2(n_81),
.B(n_317),
.Y(n_316)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_79),
.Y(n_262)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_105),
.CI(n_117),
.CON(n_104),
.SN(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_105),
.C(n_117),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_90),
.A2(n_91),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.C(n_101),
.Y(n_91)
);

FAx1_ASAP7_75t_L g290 ( 
.A(n_92),
.B(n_97),
.CI(n_101),
.CON(n_290),
.SN(n_290)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_93),
.B(n_95),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_185),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_100),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_100),
.B1(n_112),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_99),
.A2(n_100),
.B1(n_141),
.B2(n_164),
.Y(n_163)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_104),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_116),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_107),
.B1(n_122),
.B2(n_130),
.Y(n_121)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_110),
.C(n_115),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_107),
.B(n_130),
.C(n_131),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_113),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_115),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_113),
.B(n_123),
.C(n_127),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_119),
.B(n_120),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_131),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_125),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_128),
.Y(n_317)
);

AOI321xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_288),
.A3(n_296),
.B1(n_301),
.B2(n_306),
.C(n_330),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_187),
.C(n_199),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_169),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_135),
.B(n_169),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_154),
.C(n_161),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_136),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_149),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_144),
.B2(n_145),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_145),
.C(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_151),
.B(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_154),
.A2(n_161),
.B1(n_162),
.B2(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_154),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_157),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_163),
.B(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_166),
.B(n_168),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_167),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_176),
.C(n_177),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_174),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_186),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_183),
.C(n_186),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_188),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_189),
.B(n_190),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_198),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_192),
.B(n_193),
.C(n_198),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_194),
.B(n_196),
.C(n_197),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_282),
.B(n_287),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_268),
.B(n_281),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_246),
.B(n_267),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_225),
.B(n_245),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_204),
.B(n_214),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_205),
.A2(n_206),
.B1(n_210),
.B2(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_219),
.C(n_221),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_220),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_244),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_231),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_237),
.B(n_243),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_247),
.B(n_248),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_259),
.B1(n_265),
.B2(n_266),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_254),
.B1(n_257),
.B2(n_258),
.Y(n_249)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_254),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_258),
.C(n_266),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_256),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_259),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_263),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_277),
.C(n_279),
.Y(n_283)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_277),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_293),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_291),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_290),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_324),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_312),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_322),
.B2(n_323),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);


endmodule