module fake_jpeg_24114_n_177 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_26),
.B(n_15),
.Y(n_51)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_24),
.Y(n_38)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_21),
.Y(n_48)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_31),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_24),
.B1(n_14),
.B2(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_35),
.B1(n_27),
.B2(n_34),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_64),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_30),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_61),
.Y(n_84)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_24),
.B1(n_32),
.B2(n_13),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_31),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_32),
.B1(n_13),
.B2(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_35),
.B1(n_40),
.B2(n_27),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

XNOR2x1_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_29),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_50),
.C(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_40),
.B1(n_27),
.B2(n_34),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_47),
.C(n_37),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_83),
.C(n_47),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_80),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_71),
.B(n_62),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_30),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_88),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_76),
.B1(n_77),
.B2(n_29),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_90),
.B(n_94),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_69),
.C(n_79),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_36),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_99),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_95),
.C(n_96),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_107),
.B1(n_97),
.B2(n_96),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_70),
.B1(n_78),
.B2(n_59),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_109),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_99),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_70),
.B(n_55),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_36),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_42),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_42),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_91),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_126),
.C(n_127),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_119),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_102),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_94),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_128),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_103),
.B1(n_100),
.B2(n_23),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_95),
.C(n_94),
.Y(n_127)
);

OAI322xp33_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_85),
.A3(n_60),
.B1(n_61),
.B2(n_9),
.C1(n_11),
.C2(n_12),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_129),
.B(n_101),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_111),
.B(n_115),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_120),
.B(n_124),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_114),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_112),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_126),
.C(n_125),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_103),
.B1(n_100),
.B2(n_23),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_127),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_144),
.B1(n_131),
.B2(n_136),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_133),
.C(n_137),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_133),
.C(n_21),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_10),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_10),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_156),
.C(n_158),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_154),
.B(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_157),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_25),
.C(n_22),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_54),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_20),
.B(n_18),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_149),
.B(n_148),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_161),
.B(n_1),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_143),
.B(n_150),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_54),
.B1(n_12),
.B2(n_9),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_1),
.B(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_21),
.Y(n_168)
);

NOR2x1p5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_1),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_169),
.C1(n_170),
.C2(n_171),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_7),
.B(n_8),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_7),
.Y(n_177)
);


endmodule