module fake_jpeg_22332_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_24),
.Y(n_54)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_60),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_28),
.B1(n_18),
.B2(n_27),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_56),
.B1(n_39),
.B2(n_45),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_57),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_29),
.B1(n_27),
.B2(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_22),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_29),
.B1(n_17),
.B2(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_66),
.B1(n_58),
.B2(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_33),
.B1(n_17),
.B2(n_34),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_73),
.B1(n_39),
.B2(n_36),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_70),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_20),
.B1(n_17),
.B2(n_16),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_67),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_23),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_39),
.A2(n_20),
.B1(n_30),
.B2(n_26),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_75),
.A2(n_108),
.B1(n_69),
.B2(n_51),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_80),
.Y(n_114)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_46),
.B(n_26),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_96),
.C(n_24),
.Y(n_137)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_90),
.Y(n_118)
);

AO22x2_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_46),
.B1(n_36),
.B2(n_39),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_97),
.B1(n_111),
.B2(n_56),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_110),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_46),
.C(n_44),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_45),
.B1(n_44),
.B2(n_40),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_103),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_25),
.Y(n_102)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_106),
.B1(n_50),
.B2(n_47),
.Y(n_131)
);

CKINVDCx9p33_ASAP7_75t_R g105 ( 
.A(n_47),
.Y(n_105)
);

CKINVDCx11_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_14),
.Y(n_107)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_111),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_120),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_84),
.B1(n_103),
.B2(n_80),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_85),
.B1(n_84),
.B2(n_97),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_132),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_110),
.B(n_84),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_91),
.C(n_82),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_31),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_14),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_12),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_100),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_140),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_143),
.A2(n_144),
.B1(n_170),
.B2(n_126),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_84),
.B1(n_96),
.B2(n_108),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_145),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_98),
.B1(n_81),
.B2(n_82),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_148),
.B(n_156),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_98),
.B(n_95),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_164),
.Y(n_179)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_167),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_78),
.C(n_104),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_122),
.C(n_133),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_152),
.B(n_165),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_106),
.B1(n_93),
.B2(n_105),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_130),
.A2(n_93),
.B1(n_78),
.B2(n_83),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_0),
.B(n_1),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_79),
.B1(n_82),
.B2(n_109),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_1),
.B(n_2),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_173),
.B(n_7),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_109),
.B1(n_23),
.B2(n_21),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_161),
.B1(n_171),
.B2(n_117),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_76),
.B1(n_21),
.B2(n_3),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_21),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_114),
.B(n_12),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_1),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_6),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_1),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_76),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_174),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_115),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_4),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_5),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_115),
.B(n_6),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_176),
.B(n_142),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_179),
.C(n_151),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_178),
.B(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_188),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_144),
.B(n_122),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_139),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_193),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_192),
.A2(n_173),
.B(n_166),
.Y(n_231)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_200),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_204),
.B1(n_170),
.B2(n_175),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_143),
.A2(n_119),
.B1(n_141),
.B2(n_124),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_201),
.B1(n_209),
.B2(n_171),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_119),
.C(n_141),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_203),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_147),
.A2(n_149),
.B1(n_145),
.B2(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_208),
.Y(n_219)
);

AOI32xp33_ASAP7_75t_L g203 ( 
.A1(n_147),
.A2(n_121),
.A3(n_124),
.B1(n_123),
.B2(n_135),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_155),
.A2(n_142),
.B1(n_135),
.B2(n_139),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_117),
.B(n_135),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_210),
.B(n_180),
.Y(n_226)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_121),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_126),
.Y(n_224)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_167),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_216),
.C(n_217),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_202),
.B1(n_208),
.B2(n_198),
.Y(n_250)
);

BUFx12f_ASAP7_75t_SL g213 ( 
.A(n_199),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_225),
.B(n_226),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_214),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_146),
.C(n_164),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_146),
.C(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_227),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_224),
.B(n_231),
.Y(n_240)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_237),
.B1(n_238),
.B2(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_182),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_166),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_233),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_173),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_193),
.A2(n_173),
.B1(n_121),
.B2(n_126),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_191),
.A2(n_173),
.B1(n_123),
.B2(n_9),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_251),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_244),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_236),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_213),
.B(n_195),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_182),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_230),
.B1(n_233),
.B2(n_211),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_186),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_258),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_219),
.A2(n_195),
.B1(n_204),
.B2(n_178),
.Y(n_253)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_181),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_259),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_220),
.B(n_183),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_232),
.A2(n_177),
.B1(n_194),
.B2(n_192),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_260),
.A2(n_250),
.B1(n_217),
.B2(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_221),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_223),
.B(n_192),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_229),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_240),
.A3(n_246),
.B1(n_251),
.B2(n_239),
.C1(n_228),
.C2(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_266),
.B(n_279),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_257),
.A2(n_226),
.B(n_222),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_278),
.B(n_248),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_269),
.Y(n_284)
);

BUFx12_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_234),
.B(n_225),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_243),
.B(n_216),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_245),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_286),
.Y(n_310)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_245),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_260),
.B1(n_259),
.B2(n_241),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_276),
.B1(n_268),
.B2(n_275),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_242),
.B(n_221),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_294),
.B(n_295),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_263),
.A2(n_247),
.B(n_255),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_255),
.B(n_262),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_185),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_298),
.C(n_280),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_123),
.C(n_8),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_299),
.B(n_298),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_308),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_281),
.C(n_264),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_302),
.A2(n_303),
.B(n_272),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_285),
.C(n_281),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_309),
.B1(n_287),
.B2(n_271),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_267),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_309),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_269),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_284),
.A2(n_272),
.B1(n_277),
.B2(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_277),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_302),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_315),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_316),
.B1(n_305),
.B2(n_299),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_294),
.B(n_288),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_320),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_321),
.C(n_310),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_269),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_286),
.Y(n_321)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_321),
.A3(n_283),
.B1(n_123),
.B2(n_10),
.C1(n_7),
.C2(n_9),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_315),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_328),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_325),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_311),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_329),
.A2(n_323),
.B(n_326),
.Y(n_333)
);

OAI221xp5_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_123),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_330),
.A2(n_331),
.B1(n_7),
.B2(n_10),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_333),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_332),
.B1(n_334),
.B2(n_322),
.Y(n_337)
);


endmodule