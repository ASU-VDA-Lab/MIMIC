module fake_jpeg_498_n_142 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_54),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_0),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_34),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_47),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_36),
.B1(n_45),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_65),
.B1(n_55),
.B2(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_36),
.B1(n_41),
.B2(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_75),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_77),
.B1(n_73),
.B2(n_60),
.Y(n_92)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_78),
.Y(n_89)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_47),
.B1(n_38),
.B2(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_35),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_38),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_66),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_92),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_68),
.B1(n_72),
.B2(n_76),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_32),
.B(n_17),
.C(n_21),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_94),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_42),
.B1(n_58),
.B2(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_93),
.B1(n_60),
.B2(n_5),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_60),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_2),
.Y(n_94)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_2),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_15),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_101),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_108),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_3),
.B(n_6),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_105),
.C(n_8),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_6),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_18),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g115 ( 
.A(n_109),
.B(n_7),
.CON(n_115),
.SN(n_115)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_7),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_118),
.B1(n_108),
.B2(n_98),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_120),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_12),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_24),
.B(n_28),
.C(n_13),
.D(n_14),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_23),
.B(n_27),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_127),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_103),
.B(n_109),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_129),
.B(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_12),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_123),
.C(n_114),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_116),
.C(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_134),
.B(n_117),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_124),
.B(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_135),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_118),
.B(n_117),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_121),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_115),
.Y(n_142)
);


endmodule