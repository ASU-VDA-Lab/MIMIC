module real_aes_233_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g200 ( .A(n_0), .B(n_147), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_1), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_2), .B(n_131), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_3), .B(n_149), .Y(n_559) );
INVx1_ASAP7_75t_L g138 ( .A(n_4), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_5), .B(n_131), .Y(n_130) );
NAND2xp33_ASAP7_75t_SL g244 ( .A(n_6), .B(n_137), .Y(n_244) );
INVx1_ASAP7_75t_L g236 ( .A(n_7), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_8), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_9), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g125 ( .A(n_10), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g497 ( .A(n_11), .B(n_242), .Y(n_497) );
AND2x2_ASAP7_75t_L g561 ( .A(n_12), .B(n_176), .Y(n_561) );
INVx2_ASAP7_75t_L g127 ( .A(n_13), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_14), .B(n_149), .Y(n_543) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_15), .Y(n_108) );
AOI221x1_ASAP7_75t_L g239 ( .A1(n_16), .A2(n_140), .B1(n_240), .B2(n_242), .C(n_243), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_17), .B(n_131), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_18), .B(n_131), .Y(n_516) );
INVx1_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_20), .A2(n_66), .B1(n_436), .B2(n_437), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_20), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_21), .A2(n_92), .B1(n_131), .B2(n_180), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_22), .A2(n_140), .B(n_145), .Y(n_139) );
AOI221xp5_ASAP7_75t_SL g210 ( .A1(n_23), .A2(n_37), .B1(n_131), .B2(n_140), .C(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_24), .B(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g128 ( .A(n_25), .B(n_90), .Y(n_128) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_25), .A2(n_90), .B(n_127), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_26), .B(n_149), .Y(n_227) );
INVxp67_ASAP7_75t_L g238 ( .A(n_27), .Y(n_238) );
AND2x2_ASAP7_75t_L g171 ( .A(n_28), .B(n_161), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_29), .B(n_780), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_30), .A2(n_140), .B(n_199), .Y(n_198) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_31), .A2(n_242), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_32), .B(n_149), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_33), .A2(n_140), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_34), .B(n_149), .Y(n_532) );
AND2x2_ASAP7_75t_L g137 ( .A(n_35), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g141 ( .A(n_35), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g188 ( .A(n_35), .Y(n_188) );
OR2x6_ASAP7_75t_L g110 ( .A(n_36), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_38), .B(n_131), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_39), .A2(n_83), .B1(n_140), .B2(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_40), .B(n_149), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_41), .B(n_131), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_42), .B(n_147), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_43), .A2(n_140), .B(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_44), .A2(n_51), .B1(n_465), .B2(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_44), .Y(n_466) );
AND2x2_ASAP7_75t_L g203 ( .A(n_45), .B(n_161), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_46), .B(n_147), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_47), .B(n_161), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_48), .B(n_131), .Y(n_540) );
INVx1_ASAP7_75t_L g134 ( .A(n_49), .Y(n_134) );
INVx1_ASAP7_75t_L g144 ( .A(n_49), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g115 ( .A1(n_50), .A2(n_53), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_50), .Y(n_117) );
INVx1_ASAP7_75t_L g465 ( .A(n_51), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_52), .B(n_149), .Y(n_495) );
AOI221xp5_ASAP7_75t_L g103 ( .A1(n_53), .A2(n_104), .B1(n_442), .B2(n_449), .C(n_458), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_53), .Y(n_116) );
AND2x2_ASAP7_75t_L g507 ( .A(n_53), .B(n_161), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_54), .B(n_131), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_55), .B(n_147), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_56), .B(n_147), .Y(n_531) );
AND2x2_ASAP7_75t_L g162 ( .A(n_57), .B(n_161), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_58), .B(n_131), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_59), .B(n_149), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_60), .B(n_131), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_61), .A2(n_140), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_62), .B(n_147), .Y(n_158) );
AND2x2_ASAP7_75t_SL g228 ( .A(n_63), .B(n_126), .Y(n_228) );
AND2x2_ASAP7_75t_L g522 ( .A(n_64), .B(n_126), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_65), .A2(n_140), .B(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_66), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_67), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_68), .B(n_176), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_69), .B(n_147), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_70), .B(n_147), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_71), .A2(n_94), .B1(n_140), .B2(n_186), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_72), .B(n_149), .Y(n_519) );
INVx1_ASAP7_75t_L g136 ( .A(n_73), .Y(n_136) );
INVx1_ASAP7_75t_L g142 ( .A(n_73), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_74), .B(n_147), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_75), .A2(n_140), .B(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_76), .A2(n_140), .B(n_485), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_77), .A2(n_140), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g534 ( .A(n_78), .B(n_126), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_79), .A2(n_462), .B1(n_463), .B2(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_79), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_80), .B(n_161), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_81), .B(n_131), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_82), .A2(n_85), .B1(n_131), .B2(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g113 ( .A(n_84), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_86), .B(n_147), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_87), .B(n_147), .Y(n_213) );
AND2x2_ASAP7_75t_L g488 ( .A(n_88), .B(n_176), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_89), .A2(n_140), .B(n_156), .Y(n_155) );
XNOR2xp5_ASAP7_75t_L g460 ( .A(n_91), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_93), .B(n_149), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_95), .A2(n_140), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_96), .B(n_149), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_97), .B(n_131), .Y(n_202) );
INVxp67_ASAP7_75t_L g241 ( .A(n_98), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_99), .B(n_149), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_100), .A2(n_140), .B(n_225), .Y(n_224) );
BUFx2_ASAP7_75t_L g521 ( .A(n_101), .Y(n_521) );
BUFx2_ASAP7_75t_L g448 ( .A(n_102), .Y(n_448) );
BUFx2_ASAP7_75t_SL g455 ( .A(n_102), .Y(n_455) );
OAI21x1_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_114), .B(n_438), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx2_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g441 ( .A(n_107), .Y(n_441) );
BUFx2_ASAP7_75t_L g457 ( .A(n_107), .Y(n_457) );
BUFx2_ASAP7_75t_L g787 ( .A(n_107), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_108), .Y(n_470) );
OR2x2_ASAP7_75t_L g781 ( .A(n_108), .B(n_110), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_SL g458 ( .A1(n_109), .A2(n_459), .B(n_779), .C(n_782), .Y(n_458) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
XOR2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
XNOR2x1_ASAP7_75t_L g118 ( .A(n_119), .B(n_435), .Y(n_118) );
INVx3_ASAP7_75t_SL g471 ( .A(n_119), .Y(n_471) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_365), .Y(n_119) );
NOR4xp25_ASAP7_75t_SL g120 ( .A(n_121), .B(n_258), .C(n_302), .D(n_329), .Y(n_120) );
OAI221xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_219), .B1(n_229), .B2(n_246), .C(n_248), .Y(n_121) );
AOI32xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_172), .A3(n_192), .B1(n_204), .B2(n_215), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_123), .B(n_401), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_123), .A2(n_371), .B1(n_429), .B2(n_432), .Y(n_428) );
AND2x4_ASAP7_75t_SL g123 ( .A(n_124), .B(n_152), .Y(n_123) );
INVx5_ASAP7_75t_L g218 ( .A(n_124), .Y(n_218) );
OR2x2_ASAP7_75t_L g247 ( .A(n_124), .B(n_217), .Y(n_247) );
AND2x4_ASAP7_75t_L g249 ( .A(n_124), .B(n_164), .Y(n_249) );
INVx2_ASAP7_75t_L g264 ( .A(n_124), .Y(n_264) );
OR2x2_ASAP7_75t_L g276 ( .A(n_124), .B(n_173), .Y(n_276) );
AND2x2_ASAP7_75t_L g283 ( .A(n_124), .B(n_163), .Y(n_283) );
AND2x2_ASAP7_75t_SL g325 ( .A(n_124), .B(n_206), .Y(n_325) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_124), .Y(n_382) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_126), .Y(n_161) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x4_ASAP7_75t_L g151 ( .A(n_127), .B(n_128), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_139), .B(n_151), .Y(n_129) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
INVx1_ASAP7_75t_L g245 ( .A(n_132), .Y(n_245) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
AND2x6_ASAP7_75t_L g147 ( .A(n_133), .B(n_142), .Y(n_147) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g149 ( .A(n_135), .B(n_144), .Y(n_149) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx5_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
AND2x2_ASAP7_75t_L g143 ( .A(n_138), .B(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_138), .Y(n_183) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
BUFx3_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
INVx2_ASAP7_75t_L g190 ( .A(n_142), .Y(n_190) );
AND2x4_ASAP7_75t_L g186 ( .A(n_143), .B(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_148), .B(n_150), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_147), .B(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_150), .A2(n_157), .B(n_158), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_150), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_150), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_150), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_150), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_150), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_150), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_150), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_150), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_150), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_150), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_150), .A2(n_558), .B(n_559), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_151), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_151), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_151), .B(n_241), .Y(n_240) );
NOR3xp33_ASAP7_75t_L g243 ( .A(n_151), .B(n_244), .C(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_151), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_151), .A2(n_540), .B(n_541), .Y(n_539) );
INVx3_ASAP7_75t_SL g277 ( .A(n_152), .Y(n_277) );
AND2x2_ASAP7_75t_L g296 ( .A(n_152), .B(n_218), .Y(n_296) );
AOI32xp33_ASAP7_75t_L g411 ( .A1(n_152), .A2(n_282), .A3(n_312), .B1(n_342), .B2(n_377), .Y(n_411) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_163), .Y(n_152) );
AND2x2_ASAP7_75t_L g251 ( .A(n_153), .B(n_173), .Y(n_251) );
OR2x2_ASAP7_75t_L g267 ( .A(n_153), .B(n_164), .Y(n_267) );
INVx1_ASAP7_75t_L g290 ( .A(n_153), .Y(n_290) );
INVx2_ASAP7_75t_L g306 ( .A(n_153), .Y(n_306) );
AND2x2_ASAP7_75t_L g343 ( .A(n_153), .B(n_206), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_153), .B(n_164), .Y(n_362) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_153), .Y(n_431) );
AO21x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_160), .B(n_162), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_159), .Y(n_154) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_160), .A2(n_165), .B(n_171), .Y(n_164) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_160), .A2(n_165), .B(n_171), .Y(n_217) );
AOI21x1_ASAP7_75t_L g554 ( .A1(n_160), .A2(n_555), .B(n_561), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_161), .Y(n_160) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_161), .A2(n_210), .B(n_214), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_161), .A2(n_483), .B(n_484), .Y(n_482) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_161), .A2(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g398 ( .A(n_164), .B(n_173), .Y(n_398) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_164), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_170), .Y(n_165) );
OR2x2_ASAP7_75t_L g246 ( .A(n_172), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g252 ( .A(n_172), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g265 ( .A(n_172), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g427 ( .A(n_172), .B(n_296), .Y(n_427) );
BUFx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g356 ( .A(n_173), .B(n_306), .Y(n_356) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_174), .Y(n_206) );
AOI21x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_178), .B(n_191), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_176), .A2(n_223), .B(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_176), .A2(n_516), .B(n_517), .Y(n_515) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx3_ASAP7_75t_L g196 ( .A(n_177), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_185), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_180), .A2(n_186), .B1(n_235), .B2(n_237), .Y(n_234) );
AND2x4_ASAP7_75t_L g180 ( .A(n_181), .B(n_184), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2x1p5_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_192), .B(n_323), .Y(n_425) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_193), .B(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g208 ( .A(n_194), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g230 ( .A(n_194), .Y(n_230) );
AND2x2_ASAP7_75t_L g256 ( .A(n_194), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_194), .B(n_232), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_194), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g314 ( .A(n_194), .Y(n_314) );
OR2x2_ASAP7_75t_L g333 ( .A(n_194), .B(n_260), .Y(n_333) );
INVx1_ASAP7_75t_L g340 ( .A(n_194), .Y(n_340) );
NOR2xp33_ASAP7_75t_R g392 ( .A(n_194), .B(n_221), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_194), .B(n_233), .Y(n_396) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21x1_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_203), .Y(n_195) );
INVx4_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_196), .A2(n_491), .B(n_497), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
AOI32xp33_ASAP7_75t_L g419 ( .A1(n_204), .A2(n_255), .A3(n_420), .B1(n_421), .B2(n_422), .Y(n_419) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
INVx2_ASAP7_75t_L g286 ( .A(n_206), .Y(n_286) );
AND2x4_ASAP7_75t_L g305 ( .A(n_206), .B(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_206), .B(n_277), .Y(n_334) );
OR2x2_ASAP7_75t_L g388 ( .A(n_206), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g346 ( .A(n_207), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g404 ( .A(n_207), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_208), .B(n_221), .Y(n_370) );
AND2x2_ASAP7_75t_L g407 ( .A(n_208), .B(n_373), .Y(n_407) );
INVx2_ASAP7_75t_L g257 ( .A(n_209), .Y(n_257) );
INVx2_ASAP7_75t_L g260 ( .A(n_209), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_209), .B(n_221), .Y(n_280) );
INVx1_ASAP7_75t_L g311 ( .A(n_209), .Y(n_311) );
OR2x2_ASAP7_75t_L g337 ( .A(n_209), .B(n_221), .Y(n_337) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_209), .Y(n_389) );
BUFx3_ASAP7_75t_L g418 ( .A(n_209), .Y(n_418) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_216), .B(n_305), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_216), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_217), .B(n_290), .Y(n_289) );
OAI21xp33_ASAP7_75t_L g319 ( .A1(n_217), .A2(n_286), .B(n_304), .Y(n_319) );
OAI32xp33_ASAP7_75t_L g341 ( .A1(n_218), .A2(n_342), .A3(n_344), .B1(n_346), .B2(n_348), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_218), .B(n_305), .Y(n_414) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g347 ( .A(n_220), .Y(n_347) );
NOR2x1p5_ASAP7_75t_L g417 ( .A(n_220), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x4_ASAP7_75t_L g231 ( .A(n_221), .B(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_SL g255 ( .A(n_221), .B(n_233), .Y(n_255) );
OR2x2_ASAP7_75t_L g259 ( .A(n_221), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g294 ( .A(n_221), .Y(n_294) );
AND2x2_ASAP7_75t_L g312 ( .A(n_221), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g323 ( .A(n_221), .B(n_233), .Y(n_323) );
OR2x2_ASAP7_75t_L g385 ( .A(n_221), .B(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g402 ( .A(n_221), .B(n_333), .Y(n_402) );
INVx1_ASAP7_75t_L g434 ( .A(n_221), .Y(n_434) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_228), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_230), .B(n_311), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_231), .B(n_345), .Y(n_344) );
AOI222xp33_ASAP7_75t_L g349 ( .A1(n_231), .A2(n_350), .B1(n_355), .B2(n_357), .C1(n_360), .C2(n_363), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_231), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g377 ( .A(n_231), .B(n_256), .Y(n_377) );
AND2x2_ASAP7_75t_L g339 ( .A(n_232), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g354 ( .A(n_232), .B(n_259), .Y(n_354) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_233), .B(n_260), .Y(n_292) );
AND2x4_ASAP7_75t_L g313 ( .A(n_233), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g373 ( .A(n_233), .B(n_294), .Y(n_373) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_239), .Y(n_233) );
INVx3_ASAP7_75t_L g527 ( .A(n_242), .Y(n_527) );
INVx1_ASAP7_75t_SL g253 ( .A(n_247), .Y(n_253) );
NAND2xp33_ASAP7_75t_SL g422 ( .A(n_247), .B(n_277), .Y(n_422) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_252), .C(n_254), .Y(n_248) );
INVx2_ASAP7_75t_SL g299 ( .A(n_249), .Y(n_299) );
AND2x2_ASAP7_75t_L g303 ( .A(n_250), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_251), .B(n_299), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g324 ( .A1(n_251), .A2(n_289), .B(n_325), .C(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g401 ( .A(n_251), .B(n_382), .Y(n_401) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
AND2x4_ASAP7_75t_L g300 ( .A(n_255), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g405 ( .A(n_255), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_261), .B(n_268), .C(n_295), .Y(n_258) );
INVx2_ASAP7_75t_L g270 ( .A(n_259), .Y(n_270) );
OR2x2_ASAP7_75t_L g317 ( .A(n_259), .B(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_260), .Y(n_301) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_263), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g355 ( .A(n_263), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_263), .B(n_343), .Y(n_409) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_265), .A2(n_368), .B1(n_369), .B2(n_371), .C1(n_374), .C2(n_377), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_266), .A2(n_331), .B1(n_334), .B2(n_335), .C(n_341), .Y(n_330) );
AND2x2_ASAP7_75t_L g368 ( .A(n_266), .B(n_325), .Y(n_368) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp33_ASAP7_75t_SL g281 ( .A(n_267), .B(n_282), .Y(n_281) );
AOI221x1_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .B1(n_278), .B2(n_281), .C(n_284), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
AND2x2_ASAP7_75t_L g421 ( .A(n_271), .B(n_359), .Y(n_421) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g279 ( .A(n_272), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
OAI32xp33_ASAP7_75t_L g387 ( .A1(n_277), .A2(n_318), .A3(n_388), .B1(n_390), .B2(n_394), .Y(n_387) );
OAI21xp33_ASAP7_75t_SL g406 ( .A1(n_278), .A2(n_407), .B(n_408), .Y(n_406) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI21xp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .B(n_291), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
OR2x2_ASAP7_75t_L g288 ( .A(n_286), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g361 ( .A(n_286), .B(n_362), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_290), .A2(n_316), .B1(n_319), .B2(n_320), .C(n_324), .Y(n_315) );
INVx1_ASAP7_75t_L g391 ( .A(n_290), .Y(n_391) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_290), .Y(n_397) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OAI21xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_297), .B(n_300), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_299), .B(n_364), .Y(n_363) );
OAI21xp5_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_307), .B(n_315), .Y(n_302) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_306), .Y(n_376) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_309), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g328 ( .A(n_311), .Y(n_328) );
INVx1_ASAP7_75t_L g318 ( .A(n_313), .Y(n_318) );
AND2x2_ASAP7_75t_SL g327 ( .A(n_313), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_313), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_313), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g332 ( .A(n_323), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_328), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_330), .B(n_349), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g345 ( .A(n_333), .Y(n_345) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_SL g359 ( .A(n_337), .Y(n_359) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_339), .B(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_340), .Y(n_353) );
BUFx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_351), .B(n_354), .Y(n_350) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g364 ( .A(n_356), .Y(n_364) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g383 ( .A(n_362), .Y(n_383) );
NOR4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_399), .C(n_410), .D(n_423), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_378), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_368), .A2(n_379), .B(n_384), .C(n_387), .Y(n_378) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g390 ( .A1(n_381), .A2(n_391), .B(n_392), .C(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
OAI21xp33_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_397), .B(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_398), .B(n_430), .Y(n_429) );
OAI221xp5_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_402), .B1(n_403), .B2(n_404), .C(n_406), .Y(n_399) );
INVx1_ASAP7_75t_SL g403 ( .A(n_401), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND3xp33_ASAP7_75t_SL g410 ( .A(n_411), .B(n_412), .C(n_419), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI21xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp33_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
CKINVDCx9p33_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_SL g445 ( .A(n_446), .B(n_448), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_446), .A2(n_453), .B(n_456), .Y(n_452) );
INVx2_ASAP7_75t_L g786 ( .A(n_446), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g785 ( .A(n_448), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
CKINVDCx11_ASAP7_75t_R g453 ( .A(n_454), .Y(n_453) );
CKINVDCx8_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
XNOR2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp33_ASAP7_75t_SL g467 ( .A(n_468), .B(n_472), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_470), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_704), .Y(n_474) );
NOR2xp67_ASAP7_75t_L g475 ( .A(n_476), .B(n_623), .Y(n_475) );
NAND5xp2_ASAP7_75t_L g476 ( .A(n_477), .B(n_567), .C(n_577), .D(n_594), .E(n_610), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_503), .B1(n_545), .B2(n_549), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g551 ( .A(n_481), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g569 ( .A(n_481), .B(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g590 ( .A(n_481), .B(n_591), .Y(n_590) );
INVx4_ASAP7_75t_L g604 ( .A(n_481), .Y(n_604) );
AND2x2_ASAP7_75t_L g613 ( .A(n_481), .B(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_SL g635 ( .A(n_481), .B(n_553), .Y(n_635) );
BUFx2_ASAP7_75t_L g678 ( .A(n_481), .Y(n_678) );
AND2x2_ASAP7_75t_L g693 ( .A(n_481), .B(n_490), .Y(n_693) );
OR2x2_ASAP7_75t_L g725 ( .A(n_481), .B(n_726), .Y(n_725) );
NOR4xp25_ASAP7_75t_L g774 ( .A(n_481), .B(n_775), .C(n_776), .D(n_777), .Y(n_774) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_488), .Y(n_481) );
AOI31xp33_ASAP7_75t_L g642 ( .A1(n_489), .A2(n_643), .A3(n_645), .B(n_647), .Y(n_642) );
INVx2_ASAP7_75t_SL g759 ( .A(n_489), .Y(n_759) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
INVx2_ASAP7_75t_L g566 ( .A(n_490), .Y(n_566) );
AND2x2_ASAP7_75t_L g570 ( .A(n_490), .B(n_554), .Y(n_570) );
INVx2_ASAP7_75t_L g593 ( .A(n_490), .Y(n_593) );
AND2x2_ASAP7_75t_L g612 ( .A(n_490), .B(n_553), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_496), .Y(n_491) );
AND2x2_ASAP7_75t_L g564 ( .A(n_498), .B(n_565), .Y(n_564) );
BUFx3_ASAP7_75t_L g571 ( .A(n_498), .Y(n_571) );
INVx2_ASAP7_75t_L g589 ( .A(n_498), .Y(n_589) );
AND2x2_ASAP7_75t_L g644 ( .A(n_498), .B(n_604), .Y(n_644) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AND2x4_ASAP7_75t_L g615 ( .A(n_499), .B(n_500), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_535), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_523), .Y(n_504) );
OR2x2_ASAP7_75t_L g545 ( .A(n_505), .B(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g696 ( .A(n_505), .Y(n_696) );
OR2x2_ASAP7_75t_L g744 ( .A(n_505), .B(n_745), .Y(n_744) );
NAND2x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
OR2x2_ASAP7_75t_SL g536 ( .A(n_506), .B(n_537), .Y(n_536) );
INVx4_ASAP7_75t_L g574 ( .A(n_506), .Y(n_574) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_506), .Y(n_618) );
INVx2_ASAP7_75t_L g626 ( .A(n_506), .Y(n_626) );
OR2x2_ASAP7_75t_L g661 ( .A(n_506), .B(n_525), .Y(n_661) );
AND2x2_ASAP7_75t_L g773 ( .A(n_506), .B(n_628), .Y(n_773) );
AND2x2_ASAP7_75t_L g778 ( .A(n_506), .B(n_538), .Y(n_778) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
OR2x2_ASAP7_75t_L g537 ( .A(n_514), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g602 ( .A(n_514), .B(n_524), .Y(n_602) );
OR2x2_ASAP7_75t_L g609 ( .A(n_514), .B(n_574), .Y(n_609) );
NOR2x1_ASAP7_75t_SL g628 ( .A(n_514), .B(n_548), .Y(n_628) );
BUFx2_ASAP7_75t_L g660 ( .A(n_514), .Y(n_660) );
AND2x2_ASAP7_75t_L g669 ( .A(n_514), .B(n_574), .Y(n_669) );
AND2x2_ASAP7_75t_L g702 ( .A(n_514), .B(n_622), .Y(n_702) );
INVx2_ASAP7_75t_SL g711 ( .A(n_514), .Y(n_711) );
AND2x2_ASAP7_75t_L g714 ( .A(n_514), .B(n_525), .Y(n_714) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_522), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_523), .B(n_579), .C(n_664), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_523), .B(n_626), .Y(n_729) );
INVxp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_524), .B(n_711), .Y(n_732) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_525), .Y(n_576) );
AND2x2_ASAP7_75t_L g620 ( .A(n_525), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g685 ( .A(n_525), .B(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_534), .Y(n_526) );
AO21x1_ASAP7_75t_SL g548 ( .A1(n_527), .A2(n_528), .B(n_534), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
AND2x4_ASAP7_75t_L g580 ( .A(n_535), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g716 ( .A(n_537), .B(n_661), .Y(n_716) );
AND2x2_ASAP7_75t_L g547 ( .A(n_538), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g584 ( .A(n_538), .Y(n_584) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_538), .Y(n_601) );
INVx2_ASAP7_75t_L g622 ( .A(n_538), .Y(n_622) );
INVx1_ASAP7_75t_L g686 ( .A(n_538), .Y(n_686) );
INVx2_ASAP7_75t_L g768 ( .A(n_545), .Y(n_768) );
OR2x2_ASAP7_75t_L g632 ( .A(n_546), .B(n_609), .Y(n_632) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g772 ( .A(n_547), .B(n_669), .Y(n_772) );
AND2x2_ASAP7_75t_L g665 ( .A(n_548), .B(n_622), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_562), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_551), .A2(n_679), .B1(n_696), .B2(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g592 ( .A(n_553), .Y(n_592) );
AND2x2_ASAP7_75t_L g646 ( .A(n_553), .B(n_566), .Y(n_646) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_553), .Y(n_673) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_554), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_560), .Y(n_555) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_564), .B(n_678), .Y(n_677) );
OAI32xp33_ASAP7_75t_L g694 ( .A1(n_564), .A2(n_695), .A3(n_697), .B1(n_698), .B2(n_700), .Y(n_694) );
BUFx2_ASAP7_75t_L g579 ( .A(n_565), .Y(n_579) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g721 ( .A(n_566), .B(n_615), .Y(n_721) );
OR4x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .C(n_572), .D(n_575), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_568), .A2(n_659), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_569), .Y(n_761) );
AND2x2_ASAP7_75t_L g603 ( .A(n_570), .B(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g683 ( .A(n_570), .Y(n_683) );
INVx1_ASAP7_75t_L g699 ( .A(n_570), .Y(n_699) );
INVx1_ASAP7_75t_L g734 ( .A(n_570), .Y(n_734) );
OR2x2_ASAP7_75t_L g691 ( .A(n_571), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g735 ( .A(n_571), .B(n_736), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_572), .A2(n_609), .B1(n_653), .B2(n_672), .Y(n_674) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g718 ( .A(n_573), .B(n_627), .Y(n_718) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g585 ( .A(n_574), .Y(n_585) );
NOR2xp67_ASAP7_75t_L g600 ( .A(n_574), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g581 ( .A(n_575), .Y(n_581) );
NAND4xp25_ASAP7_75t_L g708 ( .A(n_575), .B(n_579), .C(n_660), .D(n_672), .Y(n_708) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g745 ( .A(n_576), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_580), .B1(n_582), .B2(n_586), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_578), .A2(n_579), .B1(n_729), .B2(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVxp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx3_ASAP7_75t_L g607 ( .A(n_584), .Y(n_607) );
AOI32xp33_ASAP7_75t_L g723 ( .A1(n_584), .A2(n_724), .A3(n_728), .B1(n_733), .B2(n_737), .Y(n_723) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
NOR2xp67_ASAP7_75t_L g629 ( .A(n_587), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g682 ( .A(n_587), .B(n_683), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_587), .A2(n_595), .B1(n_707), .B2(n_712), .C(n_715), .Y(n_706) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g639 ( .A(n_588), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g754 ( .A(n_588), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_589), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g596 ( .A(n_591), .Y(n_596) );
AND2x2_ASAP7_75t_L g614 ( .A(n_591), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_SL g654 ( .A(n_592), .Y(n_654) );
INVx1_ASAP7_75t_L g638 ( .A(n_593), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B1(n_603), .B2(n_605), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g740 ( .A(n_596), .B(n_670), .Y(n_740) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g680 ( .A(n_599), .Y(n_680) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
AND2x2_ASAP7_75t_L g611 ( .A(n_604), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_604), .B(n_641), .Y(n_640) );
NAND2x1p5_ASAP7_75t_L g653 ( .A(n_604), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_604), .B(n_646), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g764 ( .A1(n_605), .A2(n_765), .B1(n_766), .B2(n_768), .Y(n_764) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x2_ASAP7_75t_L g647 ( .A(n_607), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g657 ( .A(n_607), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_607), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_607), .B(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_SL g712 ( .A(n_607), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g688 ( .A(n_609), .B(n_689), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B(n_616), .Y(n_610) );
INVx1_ASAP7_75t_L g630 ( .A(n_612), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_613), .A2(n_650), .B1(n_657), .B2(n_662), .Y(n_649) );
INVx3_ASAP7_75t_L g652 ( .A(n_615), .Y(n_652) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
OAI32xp33_ASAP7_75t_SL g707 ( .A1(n_618), .A2(n_678), .A3(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g627 ( .A(n_621), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND4xp25_ASAP7_75t_SL g623 ( .A(n_624), .B(n_649), .C(n_666), .D(n_681), .Y(n_623) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_629), .B1(n_631), .B2(n_633), .C(n_642), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx2_ASAP7_75t_L g664 ( .A(n_626), .Y(n_664) );
AND2x2_ASAP7_75t_L g713 ( .A(n_626), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_626), .B(n_665), .Y(n_751) );
AND2x2_ASAP7_75t_L g762 ( .A(n_626), .B(n_685), .Y(n_762) );
INVx2_ASAP7_75t_L g648 ( .A(n_628), .Y(n_648) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_639), .Y(n_633) );
AND2x2_ASAP7_75t_L g765 ( .A(n_634), .B(n_636), .Y(n_765) );
INVx2_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_635), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g742 ( .A(n_640), .Y(n_742) );
INVx1_ASAP7_75t_L g727 ( .A(n_641), .Y(n_727) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_644), .B(n_699), .Y(n_698) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_645), .B(n_652), .Y(n_656) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g755 ( .A(n_646), .Y(n_755) );
INVx1_ASAP7_75t_L g737 ( .A(n_648), .Y(n_737) );
OR2x2_ASAP7_75t_L g753 ( .A(n_648), .B(n_664), .Y(n_753) );
NAND2xp33_ASAP7_75t_SL g650 ( .A(n_651), .B(n_655), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx2_ASAP7_75t_L g670 ( .A(n_652), .Y(n_670) );
AND2x2_ASAP7_75t_L g675 ( .A(n_652), .B(n_665), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_652), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g749 ( .A(n_653), .Y(n_749) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_658), .A2(n_739), .B1(n_741), .B2(n_743), .Y(n_738) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g703 ( .A(n_661), .Y(n_703) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g689 ( .A(n_665), .Y(n_689) );
AOI322xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .A3(n_671), .B1(n_674), .B2(n_675), .C1(n_676), .C2(n_679), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g717 ( .A1(n_667), .A2(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g684 ( .A(n_669), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g741 ( .A(n_670), .B(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_677), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g697 ( .A(n_678), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_678), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_687), .B2(n_690), .C(n_694), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g769 ( .A1(n_683), .A2(n_770), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_685), .B(n_696), .Y(n_695) );
BUFx2_ASAP7_75t_L g736 ( .A(n_686), .Y(n_736) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI21xp5_ASAP7_75t_L g760 ( .A1(n_690), .A2(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp33_ASAP7_75t_SL g770 ( .A(n_699), .B(n_771), .Y(n_770) );
INVx3_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
NOR4xp75_ASAP7_75t_L g704 ( .A(n_705), .B(n_722), .C(n_746), .D(n_763), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_717), .Y(n_705) );
INVx1_ASAP7_75t_L g776 ( .A(n_714), .Y(n_776) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g748 ( .A(n_721), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g775 ( .A(n_721), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_723), .B(n_738), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_SL g771 ( .A(n_742), .Y(n_771) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NAND3x1_ASAP7_75t_L g746 ( .A(n_747), .B(n_756), .C(n_760), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_750), .B(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_769), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_787), .Y(n_783) );
INVxp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
endmodule