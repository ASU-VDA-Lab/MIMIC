module fake_jpeg_2307_n_663 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_663);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_663;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_483;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_540;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_554;
wire n_280;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_419;
wire n_378;
wire n_133;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_12),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_12),
.B(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx8_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_58),
.B(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_61),
.B(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g203 ( 
.A(n_63),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_70),
.B(n_14),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_71),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_74),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_75),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_15),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_77),
.Y(n_196)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_83),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_84),
.B(n_99),
.Y(n_211)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_85),
.Y(n_195)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_92),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_95),
.Y(n_218)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_36),
.B(n_17),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_98),
.B(n_111),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_40),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_100),
.Y(n_192)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_101),
.Y(n_207)
);

INVx2_ASAP7_75t_R g102 ( 
.A(n_56),
.Y(n_102)
);

NAND2x1_ASAP7_75t_SL g161 ( 
.A(n_102),
.B(n_52),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_105),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_22),
.Y(n_110)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_40),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_40),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_116),
.Y(n_169)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_114),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_44),
.B(n_17),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_122),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_23),
.Y(n_121)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_41),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_41),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_123),
.B(n_127),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_125),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_23),
.Y(n_128)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_41),
.B(n_17),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_50),
.Y(n_181)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_91),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_139),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_143),
.B(n_185),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_76),
.A2(n_129),
.B1(n_46),
.B2(n_44),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_147),
.B(n_229),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_148),
.B(n_149),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_83),
.B(n_50),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_81),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_153),
.B(n_183),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_38),
.Y(n_157)
);

NAND2xp33_ASAP7_75t_SL g295 ( 
.A(n_157),
.B(n_1),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_161),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_165),
.Y(n_283)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_168),
.Y(n_248)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_172),
.Y(n_280)
);

BUFx12_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g297 ( 
.A(n_176),
.Y(n_297)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

NOR2x1_ASAP7_75t_R g273 ( 
.A(n_181),
.B(n_53),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_109),
.B(n_51),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_82),
.B(n_38),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_64),
.B(n_27),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_187),
.B(n_188),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_90),
.B(n_43),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_85),
.B(n_52),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_191),
.B(n_193),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_59),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_92),
.B(n_31),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_217),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_97),
.B(n_51),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_200),
.B(n_204),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_106),
.B(n_47),
.Y(n_204)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_60),
.Y(n_214)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_214),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_62),
.B(n_34),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_216),
.B(n_228),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_67),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

BUFx4f_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_69),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_74),
.Y(n_224)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_114),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

BUFx12_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

INVx13_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_75),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_35),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_106),
.B(n_47),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_77),
.B(n_43),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_167),
.A2(n_126),
.B1(n_124),
.B2(n_117),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g320 ( 
.A1(n_232),
.A2(n_281),
.B1(n_305),
.B2(n_207),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_140),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_233),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_157),
.B(n_115),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_235),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_194),
.A2(n_22),
.B1(n_78),
.B2(n_34),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_238),
.B(n_246),
.Y(n_333)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_164),
.Y(n_239)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_239),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_241),
.Y(n_350)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_242),
.Y(n_359)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_243),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_197),
.A2(n_191),
.B(n_185),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_244),
.A2(n_207),
.B(n_151),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_175),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_181),
.A2(n_103),
.B1(n_89),
.B2(n_107),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_247),
.A2(n_265),
.B1(n_306),
.B2(n_200),
.Y(n_321)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_250),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_154),
.A2(n_105),
.B1(n_104),
.B2(n_125),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_251),
.A2(n_182),
.B1(n_180),
.B2(n_196),
.Y(n_341)
);

CKINVDCx12_ASAP7_75t_R g253 ( 
.A(n_177),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_253),
.Y(n_358)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_255),
.Y(n_347)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_140),
.Y(n_256)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_132),
.Y(n_257)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_257),
.Y(n_373)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_134),
.A2(n_39),
.B(n_13),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_259),
.B(n_267),
.Y(n_327)
);

AO22x1_ASAP7_75t_SL g260 ( 
.A1(n_138),
.A2(n_115),
.B1(n_39),
.B2(n_53),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_260),
.B(n_295),
.Y(n_362)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_144),
.Y(n_261)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_154),
.A2(n_35),
.B1(n_27),
.B2(n_39),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

CKINVDCx12_ASAP7_75t_R g267 ( 
.A(n_177),
.Y(n_267)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_137),
.Y(n_269)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_269),
.Y(n_340)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_141),
.Y(n_270)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_271),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_198),
.B(n_0),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_272),
.B(n_287),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_273),
.B(n_294),
.Y(n_353)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_150),
.Y(n_276)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_276),
.Y(n_357)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_192),
.Y(n_277)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_277),
.Y(n_360)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_166),
.Y(n_279)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_279),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_213),
.A2(n_223),
.B1(n_187),
.B2(n_161),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_160),
.Y(n_284)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_284),
.Y(n_367)
);

CKINVDCx12_ASAP7_75t_R g285 ( 
.A(n_177),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_144),
.Y(n_286)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_169),
.B(n_0),
.Y(n_287)
);

INVx13_ASAP7_75t_L g288 ( 
.A(n_176),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_288),
.Y(n_335)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_178),
.Y(n_289)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_289),
.Y(n_370)
);

INVx6_ASAP7_75t_SL g290 ( 
.A(n_135),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_290),
.Y(n_363)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_146),
.Y(n_293)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_293),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_134),
.B(n_0),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_211),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_300),
.Y(n_346)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_169),
.A2(n_53),
.B(n_2),
.C(n_3),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_298),
.A2(n_219),
.B(n_6),
.C(n_7),
.Y(n_334)
);

INVx11_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_309),
.Y(n_317)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_220),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_146),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_301),
.B(n_302),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_192),
.B(n_173),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_152),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_310),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_183),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_202),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_173),
.B(n_3),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_308),
.A2(n_189),
.B1(n_163),
.B2(n_215),
.Y(n_351)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_145),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_152),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_315),
.Y(n_319)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_171),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_320),
.B(n_321),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_158),
.C(n_156),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g405 ( 
.A(n_322),
.B(n_331),
.C(n_343),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_228),
.B(n_204),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_326),
.A2(n_276),
.B(n_250),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_329),
.B(n_264),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_155),
.C(n_142),
.Y(n_331)
);

O2A1O1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_334),
.A2(n_352),
.B(n_4),
.C(n_6),
.Y(n_413)
);

NAND2x1_ASAP7_75t_L g338 ( 
.A(n_268),
.B(n_201),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g410 ( 
.A1(n_338),
.A2(n_307),
.B(n_278),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_202),
.B1(n_171),
.B2(n_180),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_339),
.A2(n_261),
.B1(n_293),
.B2(n_286),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_341),
.A2(n_310),
.B1(n_303),
.B2(n_301),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_275),
.B(n_199),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_342),
.B(n_345),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_189),
.C(n_195),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_231),
.B(n_184),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_351),
.Y(n_404)
);

OA22x2_ASAP7_75t_L g352 ( 
.A1(n_260),
.A2(n_232),
.B1(n_305),
.B2(n_237),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_162),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_354),
.B(n_364),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_235),
.B(n_206),
.C(n_182),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_241),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_205),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_245),
.B(n_205),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_234),
.Y(n_418)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

AOI21xp33_ASAP7_75t_L g460 ( 
.A1(n_379),
.A2(n_391),
.B(n_401),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_311),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_380),
.B(n_385),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_364),
.A2(n_252),
.B1(n_258),
.B2(n_212),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_381),
.A2(n_388),
.B1(n_389),
.B2(n_398),
.Y(n_427)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_382),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_383),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_342),
.B(n_252),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_384),
.B(n_387),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_324),
.B(n_243),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_354),
.B(n_230),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_321),
.A2(n_162),
.B1(n_131),
.B2(n_196),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_362),
.A2(n_131),
.B1(n_209),
.B2(n_190),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_390),
.A2(n_316),
.B1(n_376),
.B2(n_368),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_323),
.A2(n_270),
.B(n_248),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_392),
.A2(n_317),
.B(n_359),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_394),
.Y(n_448)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_360),
.Y(n_395)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_395),
.Y(n_441)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_396),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_331),
.B(n_249),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_397),
.B(n_400),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_362),
.A2(n_209),
.B1(n_208),
.B2(n_190),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_323),
.A2(n_309),
.B1(n_263),
.B2(n_240),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_399),
.A2(n_403),
.B1(n_406),
.B2(n_239),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_375),
.B(n_333),
.Y(n_400)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_326),
.B(n_288),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_362),
.A2(n_242),
.B1(n_257),
.B2(n_284),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_407),
.Y(n_453)
);

AND2x6_ASAP7_75t_L g408 ( 
.A(n_345),
.B(n_278),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_409),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_350),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_410),
.A2(n_338),
.B(n_351),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_332),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_415),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_339),
.A2(n_208),
.B1(n_145),
.B2(n_315),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_412),
.A2(n_390),
.B1(n_388),
.B2(n_341),
.Y(n_430)
);

O2A1O1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_413),
.A2(n_347),
.B(n_367),
.C(n_357),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_283),
.Y(n_415)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_356),
.Y(n_417)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_417),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_420),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_337),
.B(n_283),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_419),
.B(n_421),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_322),
.B(n_313),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_355),
.B(n_292),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_330),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_424),
.Y(n_439)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_371),
.B(n_343),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_365),
.C(n_361),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_429),
.B(n_438),
.C(n_443),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_430),
.A2(n_442),
.B1(n_373),
.B2(n_344),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_434),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_365),
.C(n_329),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_440),
.A2(n_450),
.B(n_457),
.Y(n_482)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_378),
.B(n_327),
.C(n_353),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_378),
.B(n_336),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_447),
.B(n_397),
.C(n_420),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_416),
.A2(n_352),
.B1(n_320),
.B2(n_334),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_449),
.A2(n_458),
.B1(n_465),
.B2(n_398),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_404),
.A2(n_320),
.B1(n_352),
.B2(n_335),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_383),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_452),
.B(n_456),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_320),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_391),
.A2(n_317),
.B(n_359),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_457),
.A2(n_410),
.B(n_392),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_416),
.A2(n_352),
.B1(n_318),
.B2(n_256),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_395),
.Y(n_461)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_461),
.Y(n_467)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_396),
.Y(n_462)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

OAI22x1_ASAP7_75t_L g471 ( 
.A1(n_463),
.A2(n_410),
.B1(n_418),
.B2(n_393),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_464),
.A2(n_383),
.B1(n_402),
.B2(n_407),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_416),
.A2(n_369),
.B1(n_233),
.B2(n_349),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_400),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_466),
.B(n_494),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_428),
.B(n_384),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_468),
.B(n_472),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_444),
.B(n_381),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_469),
.B(n_496),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_471),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_425),
.Y(n_472)
);

A2O1A1Ixp33_ASAP7_75t_SL g473 ( 
.A1(n_456),
.A2(n_413),
.B(n_401),
.C(n_414),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_473),
.A2(n_451),
.B(n_453),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_475),
.A2(n_480),
.B1(n_484),
.B2(n_493),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_429),
.B(n_438),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_476),
.B(n_477),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_433),
.B(n_424),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_425),
.Y(n_478)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_478),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_497),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_449),
.A2(n_414),
.B1(n_386),
.B2(n_404),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_455),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_481),
.B(n_498),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_482),
.A2(n_485),
.B(n_487),
.Y(n_515)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_441),
.Y(n_483)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_483),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_458),
.A2(n_435),
.B1(n_431),
.B2(n_436),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_486),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_450),
.A2(n_408),
.B(n_387),
.Y(n_487)
);

BUFx12_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_488),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_443),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_434),
.A2(n_422),
.B(n_347),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_490),
.A2(n_348),
.B(n_394),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_435),
.A2(n_389),
.B1(n_412),
.B2(n_403),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_446),
.B(n_370),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_SL g509 ( 
.A1(n_495),
.A2(n_430),
.B1(n_440),
.B2(n_427),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_444),
.B(n_340),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_426),
.B(n_377),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_439),
.B(n_366),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_439),
.B(n_328),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_500),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_437),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_431),
.A2(n_417),
.B1(n_423),
.B2(n_409),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_501),
.A2(n_452),
.B1(n_432),
.B2(n_427),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g524 ( 
.A1(n_502),
.A2(n_465),
.B1(n_432),
.B2(n_459),
.Y(n_524)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_503),
.Y(n_532)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_445),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_504),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_477),
.B(n_447),
.Y(n_505)
);

XNOR2x1_ASAP7_75t_L g561 ( 
.A(n_505),
.B(n_521),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_484),
.B1(n_475),
.B2(n_480),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_507),
.A2(n_524),
.B1(n_540),
.B2(n_271),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_509),
.A2(n_485),
.B1(n_471),
.B2(n_473),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_512),
.B(n_236),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_470),
.B(n_436),
.Y(n_513)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_513),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_518),
.A2(n_493),
.B1(n_501),
.B2(n_473),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_372),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_519),
.B(n_537),
.Y(n_568)
);

XOR2x1_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_437),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_476),
.B(n_462),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_474),
.Y(n_544)
);

NOR2x1_ASAP7_75t_L g523 ( 
.A(n_470),
.B(n_445),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_523),
.B(n_536),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_482),
.A2(n_460),
.B(n_463),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_525),
.A2(n_538),
.B(n_248),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_504),
.B(n_453),
.Y(n_529)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_529),
.Y(n_557)
);

A2O1A1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_533),
.A2(n_539),
.B(n_488),
.C(n_394),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_503),
.B(n_451),
.Y(n_534)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_534),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_467),
.B(n_483),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_487),
.B(n_373),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_492),
.A2(n_459),
.B(n_454),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_492),
.A2(n_454),
.B1(n_423),
.B2(n_374),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_530),
.Y(n_541)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_541),
.Y(n_578)
);

XNOR2x2_ASAP7_75t_SL g542 ( 
.A(n_533),
.B(n_473),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_542),
.B(n_540),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_474),
.C(n_490),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_543),
.B(n_547),
.C(n_550),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_544),
.B(n_548),
.Y(n_571)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_530),
.Y(n_545)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_545),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_546),
.A2(n_549),
.B1(n_562),
.B2(n_525),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_467),
.C(n_486),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_522),
.B(n_512),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_505),
.B(n_479),
.C(n_478),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_473),
.C(n_348),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_551),
.B(n_552),
.C(n_554),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_531),
.B(n_497),
.C(n_488),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_553),
.A2(n_556),
.B(n_538),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_515),
.B(n_350),
.C(n_377),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_506),
.Y(n_558)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_558),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_510),
.B(n_234),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_559),
.B(n_565),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_560),
.A2(n_514),
.B1(n_518),
.B2(n_528),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_507),
.A2(n_255),
.B1(n_280),
.B2(n_236),
.Y(n_562)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_528),
.Y(n_564)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_564),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_511),
.B(n_297),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_526),
.B(n_297),
.Y(n_566)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_566),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_567),
.B(n_534),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_563),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_570),
.B(n_573),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_568),
.B(n_526),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_574),
.A2(n_587),
.B1(n_527),
.B2(n_508),
.Y(n_612)
);

AO22x2_ASAP7_75t_L g576 ( 
.A1(n_542),
.A2(n_514),
.B1(n_521),
.B2(n_515),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_577),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_545),
.B(n_523),
.Y(n_579)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_579),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_580),
.A2(n_553),
.B1(n_549),
.B2(n_557),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_556),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_582),
.B(n_586),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_584),
.B(n_588),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_547),
.B(n_511),
.Y(n_586)
);

INVxp67_ASAP7_75t_SL g587 ( 
.A(n_555),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_548),
.B(n_544),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_543),
.B(n_506),
.C(n_513),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_589),
.B(n_581),
.C(n_585),
.Y(n_601)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_569),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_592),
.B(n_520),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_SL g595 ( 
.A(n_593),
.B(n_551),
.C(n_561),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_594),
.A2(n_596),
.B1(n_599),
.B2(n_595),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_595),
.B(n_609),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_575),
.A2(n_552),
.B1(n_562),
.B2(n_516),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_574),
.A2(n_517),
.B1(n_561),
.B2(n_536),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_597),
.A2(n_612),
.B1(n_576),
.B2(n_578),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_593),
.A2(n_550),
.B1(n_567),
.B2(n_554),
.Y(n_599)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_600),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_601),
.B(n_603),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_579),
.Y(n_603)
);

INVx11_ASAP7_75t_L g604 ( 
.A(n_590),
.Y(n_604)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_604),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_529),
.C(n_532),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_605),
.B(n_571),
.C(n_299),
.Y(n_627)
);

BUFx12_ASAP7_75t_L g608 ( 
.A(n_584),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_608),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_589),
.B(n_532),
.Y(n_609)
);

AOI31xp33_ASAP7_75t_L g610 ( 
.A1(n_591),
.A2(n_508),
.A3(n_527),
.B(n_236),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_610),
.B(n_578),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_602),
.A2(n_577),
.B1(n_583),
.B2(n_572),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_615),
.B(n_620),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g616 ( 
.A1(n_613),
.A2(n_576),
.B(n_583),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g634 ( 
.A1(n_616),
.A2(n_621),
.B(n_599),
.Y(n_634)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_618),
.Y(n_631)
);

BUFx24_ASAP7_75t_SL g619 ( 
.A(n_611),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_619),
.B(n_604),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_SL g621 ( 
.A1(n_613),
.A2(n_576),
.B(n_588),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_606),
.A2(n_607),
.B(n_594),
.Y(n_624)
);

OAI21xp33_ASAP7_75t_SL g630 ( 
.A1(n_624),
.A2(n_596),
.B(n_609),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_605),
.B(n_571),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_625),
.B(n_626),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_597),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_627),
.B(n_629),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_630),
.A2(n_629),
.B1(n_623),
.B2(n_614),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_622),
.B(n_601),
.C(n_598),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_633),
.A2(n_634),
.B(n_640),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_617),
.B(n_598),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_635),
.Y(n_644)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_638),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_608),
.Y(n_639)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_639),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_SL g640 ( 
.A1(n_616),
.A2(n_608),
.B(n_297),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_624),
.A2(n_133),
.B(n_7),
.Y(n_641)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_641),
.Y(n_645)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_637),
.B(n_623),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_642),
.B(n_647),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_636),
.A2(n_621),
.B(n_618),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_648),
.A2(n_631),
.B1(n_637),
.B2(n_639),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_644),
.B(n_632),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_651),
.A2(n_653),
.B(n_654),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_652),
.B(n_643),
.C(n_646),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_649),
.B(n_614),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_642),
.B(n_627),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_655),
.B(n_657),
.Y(n_658)
);

AOI21x1_ASAP7_75t_L g657 ( 
.A1(n_650),
.A2(n_648),
.B(n_645),
.Y(n_657)
);

AOI21xp33_ASAP7_75t_L g659 ( 
.A1(n_658),
.A2(n_656),
.B(n_7),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_4),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_660),
.B(n_4),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_661),
.B(n_7),
.Y(n_662)
);

AO22x1_ASAP7_75t_L g663 ( 
.A1(n_662),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_663)
);


endmodule