module fake_jpeg_24811_n_253 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_1),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_2),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_20),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_21),
.B(n_29),
.C(n_15),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_25),
.B(n_17),
.Y(n_67)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_20),
.B1(n_22),
.B2(n_21),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_23),
.B1(n_42),
.B2(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_57),
.B(n_63),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_22),
.B1(n_31),
.B2(n_25),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_75),
.B1(n_79),
.B2(n_84),
.Y(n_87)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_49),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_36),
.B1(n_38),
.B2(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

BUFx2_ASAP7_75t_SL g108 ( 
.A(n_76),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_38),
.B1(n_28),
.B2(n_31),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_80),
.B1(n_50),
.B2(n_44),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_31),
.B1(n_28),
.B2(n_19),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_48),
.B1(n_54),
.B2(n_42),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_52),
.B1(n_51),
.B2(n_49),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_59),
.B1(n_64),
.B2(n_56),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_92),
.B1(n_100),
.B2(n_105),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_90),
.B(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_94),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_50),
.B1(n_65),
.B2(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_65),
.B1(n_54),
.B2(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_109),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_71),
.B1(n_78),
.B2(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AO22x1_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_48),
.B1(n_34),
.B2(n_23),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_2),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_66),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_83),
.C(n_66),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_116),
.C(n_106),
.Y(n_149)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_123),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_72),
.Y(n_113)
);

NAND2xp67_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_121),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_126),
.B(n_105),
.C(n_87),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_92),
.C(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_72),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_78),
.B1(n_71),
.B2(n_74),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_109),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_78),
.B1(n_71),
.B2(n_74),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_94),
.B1(n_98),
.B2(n_76),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_34),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_133),
.Y(n_167)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_145),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_144),
.B1(n_150),
.B2(n_152),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_107),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_87),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_147),
.A2(n_143),
.B(n_141),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_154),
.C(n_155),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_3),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_129),
.B(n_127),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_4),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_5),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_116),
.B1(n_118),
.B2(n_131),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_173),
.A2(n_147),
.B1(n_113),
.B2(n_148),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_127),
.C(n_111),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_176),
.C(n_155),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_128),
.C(n_113),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_137),
.B1(n_153),
.B2(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_179),
.C(n_183),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_143),
.C(n_148),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_194),
.B1(n_160),
.B2(n_9),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_154),
.C(n_147),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_114),
.C(n_126),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_176),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_121),
.B(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_190),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_161),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_125),
.B1(n_121),
.B2(n_8),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_173),
.B1(n_169),
.B2(n_157),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_125),
.B1(n_7),
.B2(n_8),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_186),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_197),
.B(n_189),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_204),
.B1(n_205),
.B2(n_209),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_178),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_159),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_9),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_182),
.A2(n_163),
.B1(n_167),
.B2(n_166),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_164),
.B1(n_170),
.B2(n_168),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_208),
.B1(n_192),
.B2(n_194),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_160),
.B(n_9),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_187),
.B1(n_191),
.B2(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_216),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_179),
.C(n_184),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_215),
.C(n_221),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_200),
.B1(n_198),
.B2(n_204),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_192),
.C(n_180),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_202),
.B(n_188),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_187),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_218),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_5),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_14),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_229),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_221),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_199),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_208),
.B(n_206),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_230),
.A2(n_231),
.B(n_216),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_10),
.C(n_11),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_235),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_238),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_R g236 ( 
.A(n_228),
.B(n_10),
.C(n_11),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_12),
.C(n_13),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_242),
.B(n_225),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_237),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_231),
.C(n_223),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_247),
.B1(n_12),
.B2(n_13),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_13),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_250),
.Y(n_251)
);

OAI21x1_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_249),
.B(n_244),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_14),
.Y(n_253)
);


endmodule