module fake_jpeg_31226_n_212 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_4),
.B(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_10),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_53),
.Y(n_91)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_0),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_57),
.Y(n_92)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_1),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_29),
.B(n_1),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_64),
.Y(n_101)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_3),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_29),
.B(n_9),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_16),
.B(n_4),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_6),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_5),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_28),
.Y(n_79)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_71),
.B1(n_63),
.B2(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_72),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_27),
.B1(n_20),
.B2(n_24),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_34),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_31),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_96),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_38),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_26),
.B1(n_34),
.B2(n_25),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_37),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_7),
.B1(n_100),
.B2(n_86),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_73),
.Y(n_135)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_110),
.Y(n_136)
);

AND2x4_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_116),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_83),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_61),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_72),
.A2(n_50),
.B(n_36),
.C(n_45),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_43),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_125),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_68),
.C(n_50),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_113),
.B(n_121),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_34),
.B1(n_7),
.B2(n_9),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_127),
.B1(n_100),
.B2(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx11_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_76),
.A2(n_6),
.B1(n_7),
.B2(n_95),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_132),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_130),
.Y(n_155)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_98),
.B1(n_102),
.B2(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_135),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_139),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_89),
.B1(n_80),
.B2(n_97),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_154),
.B(n_121),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_107),
.B1(n_93),
.B2(n_102),
.Y(n_144)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_115),
.B(n_91),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_122),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_158),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_154),
.A2(n_112),
.B(n_109),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_168),
.C(n_145),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

AO22x2_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_116),
.B1(n_124),
.B2(n_131),
.Y(n_166)
);

AO22x2_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_109),
.B1(n_139),
.B2(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_152),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_92),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_140),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_141),
.B1(n_137),
.B2(n_138),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_176),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_137),
.B1(n_138),
.B2(n_147),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_151),
.C(n_136),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_166),
.B1(n_144),
.B2(n_156),
.Y(n_178)
);

OAI322xp33_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_159),
.A3(n_109),
.B1(n_162),
.B2(n_151),
.C1(n_168),
.C2(n_136),
.Y(n_183)
);

AOI321xp33_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_172),
.A3(n_177),
.B1(n_166),
.B2(n_181),
.C(n_173),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_163),
.C(n_142),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_185),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_163),
.C(n_142),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_186),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_166),
.C(n_155),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_189),
.C(n_124),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_177),
.B(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

AOI31xp67_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_185),
.A3(n_187),
.B(n_188),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_194),
.B(n_117),
.C(n_82),
.Y(n_204)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_194),
.C(n_153),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_129),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_117),
.A3(n_118),
.B1(n_123),
.B2(n_149),
.C1(n_114),
.C2(n_153),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_207),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_149),
.A3(n_80),
.B1(n_107),
.B2(n_130),
.C1(n_126),
.C2(n_128),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_202),
.B(n_97),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_211),
.Y(n_212)
);


endmodule