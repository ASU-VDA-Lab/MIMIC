module fake_jpeg_15646_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVxp33_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_28),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_46),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_42),
.B1(n_41),
.B2(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_45),
.B1(n_55),
.B2(n_36),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_25),
.B1(n_16),
.B2(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_58),
.Y(n_68)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_16),
.B1(n_20),
.B2(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_17),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_78),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_71),
.B(n_74),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_15),
.B1(n_23),
.B2(n_36),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_76),
.B(n_82),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_48),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_60),
.B1(n_52),
.B2(n_51),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_81),
.B1(n_59),
.B2(n_33),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_36),
.B1(n_15),
.B2(n_39),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_15),
.B(n_38),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_13),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_35),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_54),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_22),
.C(n_35),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_90),
.A2(n_83),
.B1(n_77),
.B2(n_82),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_51),
.B1(n_60),
.B2(n_59),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_106),
.B1(n_77),
.B2(n_83),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_102),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_38),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_68),
.C(n_78),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_38),
.B(n_22),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_115),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_110),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_73),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_75),
.Y(n_141)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_120),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_122),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_70),
.B1(n_77),
.B2(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_137),
.B1(n_131),
.B2(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_65),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_124),
.B1(n_129),
.B2(n_131),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_94),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_138),
.Y(n_153)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_65),
.B1(n_71),
.B2(n_74),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_113),
.B(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_64),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_135),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_137),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_139),
.B1(n_140),
.B2(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_69),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_97),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_22),
.B(n_109),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_115),
.C(n_101),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_153),
.C(n_35),
.Y(n_180)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_89),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_154),
.B(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_152),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_167),
.B(n_22),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_89),
.B(n_113),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_91),
.B1(n_96),
.B2(n_95),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_157),
.B1(n_165),
.B2(n_119),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_95),
.B1(n_93),
.B2(n_92),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_93),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_122),
.Y(n_171)
);

BUFx24_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_164),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_109),
.B1(n_100),
.B2(n_111),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_22),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_147),
.B1(n_134),
.B2(n_151),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_176),
.B1(n_193),
.B2(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_123),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_180),
.C(n_192),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_128),
.B(n_135),
.C(n_130),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_175),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_194),
.B1(n_145),
.B2(n_146),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_133),
.C(n_14),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_183),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_148),
.B(n_30),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_179),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_167),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_184),
.A2(n_183),
.B(n_181),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_124),
.B1(n_100),
.B2(n_111),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_189),
.B1(n_168),
.B2(n_164),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_56),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_190),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_149),
.A2(n_114),
.B1(n_104),
.B2(n_81),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_56),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_35),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_104),
.B1(n_32),
.B2(n_39),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_154),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_207),
.C(n_214),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_177),
.B1(n_182),
.B2(n_188),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_166),
.B1(n_156),
.B2(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_204),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_33),
.B1(n_34),
.B2(n_66),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_161),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_159),
.B1(n_155),
.B2(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_208),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_150),
.B(n_164),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_210),
.A2(n_195),
.B1(n_188),
.B2(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_142),
.C(n_157),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_184),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_142),
.C(n_162),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_164),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_189),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_35),
.C(n_87),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_87),
.C(n_67),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_228),
.B1(n_234),
.B2(n_217),
.Y(n_254)
);

AO22x2_ASAP7_75t_SL g221 ( 
.A1(n_215),
.A2(n_205),
.B1(n_213),
.B2(n_218),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_197),
.B(n_179),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_222),
.B(n_225),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_174),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_185),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_232),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_195),
.B1(n_173),
.B2(n_193),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_67),
.C(n_66),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_240),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_210),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_224),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_211),
.B(n_206),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_245),
.A2(n_255),
.B(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_212),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_250),
.B(n_252),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_207),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_227),
.C(n_223),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_29),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_209),
.B(n_219),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_204),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_230),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_198),
.B1(n_203),
.B2(n_61),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_232),
.B1(n_236),
.B2(n_226),
.Y(n_262)
);

AO221x1_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_61),
.B1(n_84),
.B2(n_29),
.C(n_26),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_61),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_235),
.B(n_220),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_267),
.B1(n_21),
.B2(n_29),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_29),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_268),
.B1(n_255),
.B2(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_241),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_270),
.C(n_243),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_248),
.B(n_230),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_251),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_242),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_84),
.C(n_34),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_10),
.B(n_14),
.Y(n_272)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_245),
.B(n_14),
.Y(n_278)
);

INVx11_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_274),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_247),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_249),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_243),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_283),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_26),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_290),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_261),
.B(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_5),
.Y(n_300)
);

O2A1O1Ixp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_265),
.B(n_26),
.C(n_30),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_293),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_21),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_291),
.B(n_276),
.Y(n_297)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_4),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_6),
.B(n_7),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_304),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_21),
.C(n_30),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_305),
.C(n_5),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_296),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_295),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_306),
.B(n_307),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_6),
.B(n_7),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_312),
.B(n_298),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_8),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_299),
.A2(n_7),
.B(n_8),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_315),
.B(n_310),
.C(n_303),
.Y(n_316)
);

OAI321xp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_314),
.A3(n_311),
.B1(n_310),
.B2(n_9),
.C(n_8),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_8),
.B1(n_9),
.B2(n_309),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_9),
.Y(n_319)
);


endmodule