module real_aes_6175_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_693;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
wire n_237;
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_0), .A2(n_197), .B1(n_404), .B2(n_406), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g407 ( .A1(n_1), .A2(n_88), .B1(n_408), .B2(n_410), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_2), .B(n_275), .Y(n_598) );
AOI22xp5_ASAP7_75t_SL g319 ( .A1(n_3), .A2(n_48), .B1(n_320), .B2(n_323), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_4), .A2(n_21), .B1(n_564), .B2(n_679), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_5), .A2(n_124), .B1(n_280), .B2(n_577), .C(n_637), .Y(n_636) );
XOR2x2_ASAP7_75t_L g421 ( .A(n_6), .B(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_7), .A2(n_105), .B1(n_281), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_8), .A2(n_20), .B1(n_531), .B2(n_533), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_9), .A2(n_153), .B1(n_351), .B2(n_425), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_10), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_11), .A2(n_181), .B1(n_413), .B2(n_414), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_12), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_13), .A2(n_118), .B1(n_453), .B2(n_535), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g605 ( .A1(n_14), .A2(n_97), .B1(n_532), .B2(n_562), .Y(n_605) );
OA22x2_ASAP7_75t_L g509 ( .A1(n_15), .A2(n_510), .B1(n_511), .B2(n_541), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_15), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g602 ( .A1(n_16), .A2(n_159), .B1(n_360), .B2(n_535), .Y(n_602) );
AOI222xp33_ASAP7_75t_L g640 ( .A1(n_17), .A2(n_106), .B1(n_135), .B2(n_500), .C1(n_558), .C2(n_641), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_18), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_19), .A2(n_192), .B1(n_414), .B2(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_22), .A2(n_188), .B1(n_618), .B2(n_670), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_23), .A2(n_211), .B1(n_339), .B2(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_24), .A2(n_150), .B1(n_404), .B2(n_416), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_25), .A2(n_215), .B1(n_287), .B2(n_335), .Y(n_709) );
AOI22xp5_ASAP7_75t_SL g313 ( .A1(n_26), .A2(n_214), .B1(n_314), .B2(n_316), .Y(n_313) );
AO22x2_ASAP7_75t_L g247 ( .A1(n_27), .A2(n_70), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g659 ( .A(n_27), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_28), .A2(n_195), .B1(n_425), .B2(n_481), .C(n_483), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_29), .A2(n_33), .B1(n_268), .B2(n_344), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_30), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_31), .A2(n_196), .B1(n_300), .B2(n_679), .Y(n_703) );
AOI222xp33_ASAP7_75t_L g498 ( .A1(n_32), .A2(n_85), .B1(n_133), .B2(n_384), .C1(n_499), .C2(n_500), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_34), .Y(n_478) );
AOI22xp5_ASAP7_75t_SL g296 ( .A1(n_35), .A2(n_116), .B1(n_297), .B2(n_300), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_36), .Y(n_705) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_37), .A2(n_107), .B1(n_166), .B2(n_681), .C1(n_682), .C2(n_683), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_38), .A2(n_212), .B1(n_288), .B2(n_558), .Y(n_557) );
AO22x2_ASAP7_75t_L g251 ( .A1(n_39), .A2(n_72), .B1(n_248), .B2(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g660 ( .A(n_39), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_40), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_41), .A2(n_53), .B1(n_458), .B2(n_579), .Y(n_578) );
AOI222xp33_ASAP7_75t_L g581 ( .A1(n_42), .A2(n_131), .B1(n_177), .B2(n_441), .C1(n_500), .C2(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_43), .B(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_44), .A2(n_221), .B1(n_420), .B2(n_433), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_45), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_46), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_47), .A2(n_198), .B1(n_300), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_49), .A2(n_119), .B1(n_288), .B2(n_458), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_50), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_51), .A2(n_199), .B1(n_430), .B2(n_431), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_52), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_54), .A2(n_160), .B1(n_360), .B2(n_405), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_55), .B(n_281), .Y(n_460) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_56), .A2(n_120), .B1(n_470), .B2(n_472), .C(n_474), .Y(n_469) );
INVx1_ASAP7_75t_L g442 ( .A(n_57), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_58), .A2(n_122), .B1(n_437), .B2(n_491), .C(n_492), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_59), .A2(n_184), .B1(n_430), .B2(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_SL g286 ( .A1(n_60), .A2(n_203), .B1(n_287), .B2(n_291), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_61), .A2(n_132), .B1(n_452), .B2(n_453), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_62), .A2(n_207), .B1(n_269), .B2(n_385), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_63), .A2(n_611), .B1(n_642), .B2(n_643), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_63), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_64), .A2(n_468), .B1(n_501), .B2(n_502), .Y(n_467) );
INVx1_ASAP7_75t_L g501 ( .A(n_64), .Y(n_501) );
AOI222xp33_ASAP7_75t_L g713 ( .A1(n_65), .A2(n_130), .B1(n_139), .B2(n_291), .C1(n_499), .C2(n_500), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_66), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_67), .A2(n_172), .B1(n_287), .B2(n_292), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_68), .A2(n_104), .B1(n_365), .B2(n_433), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_69), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_71), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_73), .A2(n_174), .B1(n_358), .B2(n_360), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_74), .B(n_280), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_75), .Y(n_616) );
INVx1_ASAP7_75t_L g230 ( .A(n_76), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_77), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_78), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_79), .A2(n_158), .B1(n_452), .B2(n_453), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_80), .A2(n_180), .B1(n_335), .B2(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_81), .A2(n_92), .B1(n_570), .B2(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g228 ( .A(n_82), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_83), .A2(n_146), .B1(n_314), .B2(n_358), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_84), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_86), .A2(n_140), .B1(n_281), .B2(n_346), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_87), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_89), .A2(n_110), .B1(n_343), .B2(n_344), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_90), .A2(n_121), .B1(n_533), .B2(n_564), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_91), .A2(n_109), .B1(n_288), .B2(n_385), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g336 ( .A(n_93), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_94), .A2(n_103), .B1(n_481), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g259 ( .A1(n_95), .A2(n_145), .B1(n_260), .B2(n_268), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_96), .A2(n_101), .B1(n_323), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_98), .A2(n_137), .B1(n_535), .B2(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_99), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_100), .A2(n_179), .B1(n_304), .B2(n_325), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_102), .A2(n_152), .B1(n_362), .B2(n_364), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_108), .A2(n_183), .B1(n_349), .B2(n_350), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_111), .A2(n_178), .B1(n_416), .B2(n_419), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_112), .Y(n_394) );
XNOR2x2_ASAP7_75t_L g566 ( .A(n_113), .B(n_567), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_114), .A2(n_663), .B1(n_664), .B2(n_685), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_114), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_115), .Y(n_258) );
INVx2_ASAP7_75t_L g231 ( .A(n_117), .Y(n_231) );
INVx1_ASAP7_75t_L g607 ( .A(n_123), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_125), .B(n_275), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_126), .B(n_436), .Y(n_555) );
AND2x6_ASAP7_75t_L g227 ( .A(n_127), .B(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_127), .Y(n_653) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_128), .A2(n_187), .B1(n_248), .B2(n_252), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_129), .A2(n_171), .B1(n_425), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_134), .A2(n_205), .B1(n_339), .B2(n_458), .Y(n_553) );
AOI22xp5_ASAP7_75t_SL g302 ( .A1(n_136), .A2(n_186), .B1(n_303), .B2(n_308), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_138), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_141), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_142), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_143), .A2(n_223), .B(n_232), .C(n_661), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_144), .A2(n_176), .B1(n_263), .B2(n_288), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_147), .B(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_148), .A2(n_220), .B1(n_436), .B2(n_437), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_149), .Y(n_475) );
AO22x2_ASAP7_75t_L g257 ( .A1(n_151), .A2(n_200), .B1(n_248), .B2(n_249), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_154), .A2(n_218), .B1(n_405), .B2(n_564), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g620 ( .A(n_155), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_156), .A2(n_185), .B1(n_405), .B2(n_413), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_157), .A2(n_206), .B1(n_308), .B2(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_161), .A2(n_182), .B1(n_323), .B2(n_477), .Y(n_574) );
INVx1_ASAP7_75t_L g326 ( .A(n_162), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_163), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_164), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_165), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_167), .A2(n_170), .B1(n_353), .B2(n_355), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_168), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_169), .A2(n_216), .B1(n_561), .B2(n_562), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_173), .B(n_275), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_175), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_187), .B(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_189), .Y(n_371) );
OA22x2_ASAP7_75t_L g327 ( .A1(n_190), .A2(n_328), .B1(n_329), .B2(n_366), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_190), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_191), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_193), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g464 ( .A1(n_194), .A2(n_219), .B1(n_322), .B2(n_418), .Y(n_464) );
INVx1_ASAP7_75t_L g656 ( .A(n_200), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_201), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_202), .B(n_280), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_204), .Y(n_378) );
INVx1_ASAP7_75t_L g248 ( .A(n_208), .Y(n_248) );
INVx1_ASAP7_75t_L g250 ( .A(n_208), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_209), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_210), .B(n_273), .Y(n_272) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_213), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_217), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_228), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_229), .A2(n_651), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_506), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_232) );
INVx1_ASAP7_75t_L g646 ( .A(n_233), .Y(n_646) );
AOI22xp5_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_235), .B1(n_446), .B2(n_505), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_236), .A2(n_237), .B1(n_368), .B2(n_369), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B1(n_327), .B2(n_367), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
XOR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_326), .Y(n_240) );
NAND3x1_ASAP7_75t_L g241 ( .A(n_242), .B(n_295), .C(n_312), .Y(n_241) );
NOR2x1_ASAP7_75t_L g242 ( .A(n_243), .B(n_271), .Y(n_242) );
OAI21xp5_ASAP7_75t_SL g243 ( .A1(n_244), .A2(n_258), .B(n_259), .Y(n_243) );
BUFx2_ASAP7_75t_L g332 ( .A(n_244), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_244), .A2(n_456), .B(n_457), .Y(n_455) );
INVx4_ASAP7_75t_L g499 ( .A(n_244), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_244), .A2(n_552), .B(n_553), .Y(n_551) );
INVx4_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_SL g387 ( .A(n_245), .Y(n_387) );
BUFx3_ASAP7_75t_L g441 ( .A(n_245), .Y(n_441) );
INVx2_ASAP7_75t_L g519 ( .A(n_245), .Y(n_519) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_245), .Y(n_681) );
AND2x6_ASAP7_75t_L g245 ( .A(n_246), .B(n_253), .Y(n_245) );
AND2x4_ASAP7_75t_L g292 ( .A(n_246), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g398 ( .A(n_246), .Y(n_398) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_251), .Y(n_246) );
AND2x2_ASAP7_75t_L g267 ( .A(n_247), .B(n_255), .Y(n_267) );
INVx2_ASAP7_75t_L g277 ( .A(n_247), .Y(n_277) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g252 ( .A(n_250), .Y(n_252) );
INVx2_ASAP7_75t_L g266 ( .A(n_251), .Y(n_266) );
AND2x2_ASAP7_75t_L g276 ( .A(n_251), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g285 ( .A(n_251), .B(n_277), .Y(n_285) );
INVx1_ASAP7_75t_L g290 ( .A(n_251), .Y(n_290) );
AND2x2_ASAP7_75t_L g298 ( .A(n_253), .B(n_299), .Y(n_298) );
AND2x6_ASAP7_75t_L g322 ( .A(n_253), .B(n_284), .Y(n_322) );
AND2x4_ASAP7_75t_L g325 ( .A(n_253), .B(n_276), .Y(n_325) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
AND2x2_ASAP7_75t_L g278 ( .A(n_254), .B(n_257), .Y(n_278) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g307 ( .A(n_255), .B(n_294), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_255), .B(n_257), .Y(n_311) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g265 ( .A(n_257), .Y(n_265) );
INVx1_ASAP7_75t_L g294 ( .A(n_257), .Y(n_294) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx4_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx2_ASAP7_75t_L g682 ( .A(n_262), .Y(n_682) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_263), .Y(n_385) );
BUFx4f_ASAP7_75t_SL g558 ( .A(n_263), .Y(n_558) );
BUFx2_ASAP7_75t_L g582 ( .A(n_263), .Y(n_582) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g270 ( .A(n_265), .Y(n_270) );
AND2x2_ASAP7_75t_L g299 ( .A(n_266), .B(n_277), .Y(n_299) );
INVx1_ASAP7_75t_L g393 ( .A(n_266), .Y(n_393) );
AND2x4_ASAP7_75t_L g269 ( .A(n_267), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g288 ( .A(n_267), .B(n_289), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_267), .B(n_393), .Y(n_392) );
BUFx4f_ASAP7_75t_SL g500 ( .A(n_268), .Y(n_500) );
INVx2_ASAP7_75t_L g684 ( .A(n_268), .Y(n_684) );
BUFx12f_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_269), .Y(n_339) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_269), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_279), .C(n_286), .Y(n_271) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g577 ( .A(n_274), .Y(n_577) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g346 ( .A(n_275), .Y(n_346) );
BUFx4f_ASAP7_75t_L g437 ( .A(n_275), .Y(n_437) );
AND2x6_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
AND2x2_ASAP7_75t_L g306 ( .A(n_276), .B(n_307), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g380 ( .A(n_276), .B(n_278), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_276), .B(n_307), .Y(n_486) );
AND2x4_ASAP7_75t_L g283 ( .A(n_278), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g301 ( .A(n_278), .B(n_299), .Y(n_301) );
INVx1_ASAP7_75t_L g377 ( .A(n_278), .Y(n_377) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g436 ( .A(n_282), .Y(n_436) );
INVx2_ASAP7_75t_L g597 ( .A(n_282), .Y(n_597) );
INVx2_ASAP7_75t_L g708 ( .A(n_282), .Y(n_708) );
INVx4_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g376 ( .A(n_285), .B(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g343 ( .A(n_288), .Y(n_343) );
INVx1_ASAP7_75t_L g580 ( .A(n_288), .Y(n_580) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x6_ASAP7_75t_L g310 ( .A(n_290), .B(n_311), .Y(n_310) );
BUFx2_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g344 ( .A(n_292), .Y(n_344) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_292), .Y(n_458) );
INVx1_ASAP7_75t_L g399 ( .A(n_293), .Y(n_399) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_302), .Y(n_295) );
BUFx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g363 ( .A(n_298), .Y(n_363) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_298), .Y(n_405) );
BUFx2_ASAP7_75t_SL g430 ( .A(n_298), .Y(n_430) );
AND2x2_ASAP7_75t_L g315 ( .A(n_299), .B(n_307), .Y(n_315) );
AND2x4_ASAP7_75t_L g317 ( .A(n_299), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_299), .B(n_307), .Y(n_635) );
BUFx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx3_ASAP7_75t_L g365 ( .A(n_301), .Y(n_365) );
BUFx3_ASAP7_75t_L g420 ( .A(n_301), .Y(n_420) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_301), .Y(n_452) );
INVx2_ASAP7_75t_L g540 ( .A(n_301), .Y(n_540) );
BUFx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g409 ( .A(n_304), .Y(n_409) );
INVx4_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g354 ( .A(n_305), .Y(n_354) );
INVx2_ASAP7_75t_L g427 ( .A(n_305), .Y(n_427) );
INVx5_ASAP7_75t_L g532 ( .A(n_305), .Y(n_532) );
INVx3_ASAP7_75t_L g564 ( .A(n_305), .Y(n_564) );
BUFx3_ASAP7_75t_L g702 ( .A(n_305), .Y(n_702) );
INVx8_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
BUFx2_ASAP7_75t_L g489 ( .A(n_309), .Y(n_489) );
BUFx2_ASAP7_75t_L g679 ( .A(n_309), .Y(n_679) );
INVx6_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g410 ( .A(n_310), .Y(n_410) );
INVx1_ASAP7_75t_L g533 ( .A(n_310), .Y(n_533) );
INVx1_ASAP7_75t_L g318 ( .A(n_311), .Y(n_318) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_319), .Y(n_312) );
INVx1_ASAP7_75t_L g473 ( .A(n_314), .Y(n_473) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx3_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
BUFx3_ASAP7_75t_L g418 ( .A(n_315), .Y(n_418) );
BUFx3_ASAP7_75t_L g535 ( .A(n_315), .Y(n_535) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx3_ASAP7_75t_L g360 ( .A(n_317), .Y(n_360) );
BUFx2_ASAP7_75t_SL g414 ( .A(n_317), .Y(n_414) );
BUFx3_ASAP7_75t_L g433 ( .A(n_317), .Y(n_433) );
BUFx3_ASAP7_75t_L g570 ( .A(n_317), .Y(n_570) );
BUFx3_ASAP7_75t_L g618 ( .A(n_317), .Y(n_618) );
AND2x2_ASAP7_75t_L g453 ( .A(n_318), .B(n_393), .Y(n_453) );
INVx1_ASAP7_75t_L g626 ( .A(n_320), .Y(n_626) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
INVx4_ASAP7_75t_L g431 ( .A(n_321), .Y(n_431) );
INVx4_ASAP7_75t_L g537 ( .A(n_321), .Y(n_537) );
INVx11_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx11_ASAP7_75t_L g359 ( .A(n_322), .Y(n_359) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g425 ( .A(n_324), .Y(n_425) );
INVx3_ASAP7_75t_L g677 ( .A(n_324), .Y(n_677) );
INVx6_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g349 ( .A(n_325), .Y(n_349) );
BUFx3_ASAP7_75t_L g406 ( .A(n_325), .Y(n_406) );
BUFx3_ASAP7_75t_L g562 ( .A(n_325), .Y(n_562) );
INVx1_ASAP7_75t_L g367 ( .A(n_327), .Y(n_367) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_347), .C(n_356), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_341), .Y(n_330) );
OAI222xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B1(n_334), .B2(n_336), .C1(n_337), .C2(n_340), .Y(n_331) );
INVx1_ASAP7_75t_L g641 ( .A(n_332), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_335), .Y(n_334) );
OAI222xp33_ASAP7_75t_L g382 ( .A1(n_337), .A2(n_383), .B1(n_386), .B2(n_387), .C1(n_388), .C2(n_389), .Y(n_382) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx4f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_352), .Y(n_347) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVxp67_ASAP7_75t_L g622 ( .A(n_355), .Y(n_622) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx5_ASAP7_75t_SL g413 ( .A(n_359), .Y(n_413) );
INVx4_ASAP7_75t_L g477 ( .A(n_359), .Y(n_477) );
INVx2_ASAP7_75t_SL g561 ( .A(n_359), .Y(n_561) );
INVx2_ASAP7_75t_L g668 ( .A(n_359), .Y(n_668) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g670 ( .A(n_363), .Y(n_670) );
INVx1_ASAP7_75t_L g615 ( .A(n_364), .Y(n_615) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_421), .B1(n_444), .B2(n_445), .Y(n_369) );
INVx2_ASAP7_75t_L g444 ( .A(n_370), .Y(n_444) );
XNOR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_401), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_382), .C(n_390), .Y(n_373) );
OAI22xp5_ASAP7_75t_SL g374 ( .A1(n_375), .A2(n_378), .B1(n_379), .B2(n_381), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_375), .A2(n_525), .B1(n_526), .B2(n_527), .Y(n_524) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g528 ( .A(n_380), .Y(n_528) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_394), .B1(n_395), .B2(n_400), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx4_ASAP7_75t_L g495 ( .A(n_392), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_392), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g516 ( .A(n_396), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g396 ( .A(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g497 ( .A(n_397), .Y(n_497) );
OR2x6_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_411), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_407), .Y(n_402) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
INVx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g445 ( .A(n_421), .Y(n_445) );
NOR4xp75_ASAP7_75t_L g422 ( .A(n_423), .B(n_428), .C(n_434), .D(n_439), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_424), .B(n_426), .Y(n_423) );
INVx2_ASAP7_75t_L g628 ( .A(n_425), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_429), .B(n_432), .Y(n_428) );
INVx1_ASAP7_75t_L g631 ( .A(n_430), .Y(n_631) );
INVx1_ASAP7_75t_L g479 ( .A(n_433), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_435), .B(n_438), .Y(n_434) );
BUFx2_ASAP7_75t_L g491 ( .A(n_436), .Y(n_491) );
OAI21xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_442), .B(n_443), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g505 ( .A(n_446), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_467), .B1(n_503), .B2(n_504), .Y(n_446) );
INVx3_ASAP7_75t_L g503 ( .A(n_447), .Y(n_503) );
XOR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_466), .Y(n_447) );
NAND3x1_ASAP7_75t_SL g448 ( .A(n_449), .B(n_454), .C(n_463), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
INVx4_ASAP7_75t_L g482 ( .A(n_452), .Y(n_482) );
NOR2x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_459), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .C(n_462), .Y(n_459) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g504 ( .A(n_467), .Y(n_504) );
INVx1_ASAP7_75t_L g502 ( .A(n_468), .Y(n_502) );
AND4x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_480), .C(n_490), .D(n_498), .Y(n_468) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_478), .B2(n_479), .Y(n_474) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_487), .B2(n_488), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_485), .A2(n_620), .B1(n_621), .B2(n_622), .Y(n_619) );
BUFx2_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_496), .B2(n_497), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_494), .A2(n_497), .B1(n_638), .B2(n_639), .Y(n_637) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g647 ( .A(n_506), .Y(n_647) );
AOI22xp5_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_585), .B1(n_586), .B2(n_645), .Y(n_506) );
INVx1_ASAP7_75t_L g645 ( .A(n_507), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_542), .B2(n_584), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g541 ( .A(n_511), .Y(n_541) );
NAND2x1_ASAP7_75t_L g511 ( .A(n_512), .B(n_529), .Y(n_511) );
NOR3xp33_ASAP7_75t_SL g512 ( .A(n_513), .B(n_517), .C(n_524), .Y(n_512) );
OAI21xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_519), .A2(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OA211x2_ASAP7_75t_L g671 ( .A1(n_527), .A2(n_672), .B(n_673), .C(n_674), .Y(n_671) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_SL g706 ( .A(n_528), .Y(n_706) );
AND4x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .C(n_536), .D(n_538), .Y(n_529) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g584 ( .A(n_542), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_566), .B2(n_583), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
XOR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_565), .Y(n_545) );
NAND3x1_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .C(n_559), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NOR2x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_557), .Y(n_554) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx2_ASAP7_75t_L g583 ( .A(n_566), .Y(n_583) );
NAND4xp75_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .C(n_575), .D(n_581), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_SL g575 ( .A(n_576), .B(n_578), .Y(n_575) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_608), .B1(n_609), .B2(n_644), .Y(n_586) );
INVx1_ASAP7_75t_L g644 ( .A(n_587), .Y(n_644) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
XOR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_607), .Y(n_589) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_591), .B(n_600), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .C(n_599), .Y(n_595) );
NOR2x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g643 ( .A(n_611), .Y(n_643) );
AND4x1_ASAP7_75t_L g611 ( .A(n_612), .B(n_623), .C(n_636), .D(n_640), .Y(n_611) );
NOR2xp33_ASAP7_75t_SL g612 ( .A(n_613), .B(n_619), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_616), .B2(n_617), .Y(n_613) );
INVxp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_629), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_627), .B2(n_628), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_632), .B2(n_633), .Y(n_629) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
NOR2x1_ASAP7_75t_L g649 ( .A(n_650), .B(n_654), .Y(n_649) );
OR2x2_ASAP7_75t_SL g716 ( .A(n_650), .B(n_655), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_651), .Y(n_688) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_652), .B(n_690), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g690 ( .A(n_653), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
OAI322xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_686), .A3(n_689), .B1(n_691), .B2(n_694), .C1(n_695), .C2(n_714), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_664), .Y(n_663) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND4xp75_ASAP7_75t_L g665 ( .A(n_666), .B(n_671), .C(n_675), .D(n_680), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
XOR2x2_ASAP7_75t_L g697 ( .A(n_694), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND4xp75_ASAP7_75t_L g698 ( .A(n_699), .B(n_704), .C(n_710), .D(n_713), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .Y(n_699) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OA211x2_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B(n_707), .C(n_709), .Y(n_704) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_716), .Y(n_715) );
endmodule