module fake_jpeg_19695_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_13),
.B1(n_10),
.B2(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_18),
.B1(n_12),
.B2(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_30),
.Y(n_35)
);

AO22x1_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_11),
.B1(n_9),
.B2(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_24),
.B(n_22),
.C(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_38),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_23),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_42),
.B(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_21),
.Y(n_43)
);

XNOR2x1_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_11),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_17),
.B(n_25),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_32),
.B1(n_29),
.B2(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_55),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_36),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_44),
.B(n_38),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_32),
.B1(n_25),
.B2(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_37),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_59),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_37),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_34),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_58),
.B1(n_60),
.B2(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_50),
.Y(n_67)
);

XOR2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_42),
.Y(n_65)
);

A2O1A1O1Ixp25_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_53),
.B(n_48),
.C(n_45),
.D(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NOR4xp25_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_54),
.C(n_46),
.D(n_49),
.Y(n_68)
);

OA21x2_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_62),
.B(n_59),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_76),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_63),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_6),
.C(n_8),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_61),
.B1(n_57),
.B2(n_55),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_86),
.C(n_70),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_52),
.B(n_11),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_74),
.B(n_31),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_11),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_83),
.Y(n_88)
);

AOI31xp67_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_92),
.A3(n_78),
.B(n_79),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_86),
.B(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_73),
.C(n_31),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_84),
.C(n_85),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_81),
.A3(n_80),
.B1(n_31),
.B2(n_18),
.C1(n_15),
.C2(n_5),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_94),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_6),
.B1(n_8),
.B2(n_7),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_81),
.C(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_18),
.A3(n_15),
.B1(n_2),
.B2(n_3),
.C1(n_1),
.C2(n_0),
.Y(n_104)
);

AOI21x1_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_5),
.B(n_7),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_4),
.A3(n_7),
.B1(n_2),
.B2(n_3),
.C1(n_0),
.C2(n_1),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_104),
.C(n_15),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_4),
.B(n_31),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_99),
.B(n_98),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.B(n_15),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_0),
.Y(n_108)
);


endmodule