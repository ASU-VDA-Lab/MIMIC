module fake_jpeg_17907_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx10_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

OR2x2_ASAP7_75t_SL g18 ( 
.A(n_15),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_3),
.Y(n_23)
);

AND2x4_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_4),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_17),
.B(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_39),
.B1(n_30),
.B2(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_42),
.B1(n_30),
.B2(n_10),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_24),
.B1(n_17),
.B2(n_19),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_47),
.B(n_36),
.C(n_8),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_27),
.B(n_24),
.C(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_45),
.B1(n_8),
.B2(n_5),
.Y(n_51)
);

AO21x2_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_19),
.B(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_49),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_35),
.B1(n_34),
.B2(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_50),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_48),
.B(n_47),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_55),
.B(n_52),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_48),
.B1(n_51),
.B2(n_46),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_8),
.C(n_36),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_8),
.Y(n_59)
);


endmodule