module real_jpeg_31771_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_0),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_40)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_43),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g161 ( 
.A1(n_1),
.A2(n_43),
.B1(n_162),
.B2(n_166),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_1),
.B(n_95),
.Y(n_259)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_1),
.A2(n_278),
.A3(n_283),
.B1(n_286),
.B2(n_294),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_1),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_1),
.B(n_195),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_3),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_3),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_4),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_5),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_6),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_6),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_6),
.Y(n_177)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_8),
.A2(n_31),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

OAI22x1_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_31),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_31),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_10),
.A2(n_228),
.B1(n_229),
.B2(n_231),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_10),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_244),
.Y(n_12)
);

NAND2xp33_ASAP7_75t_R g13 ( 
.A(n_14),
.B(n_243),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_212),
.Y(n_14)
);

INVxp33_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_16),
.B(n_213),
.Y(n_243)
);

OAI21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_143),
.B(n_211),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_18),
.B(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_78),
.Y(n_18)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_19),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_45),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_20),
.B(n_46),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_20),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_20),
.B(n_216),
.C(n_327),
.Y(n_345)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_21),
.B(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_21),
.B(n_340),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B1(n_36),
.B2(n_40),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_22),
.B(n_40),
.Y(n_157)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_22),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_23),
.B(n_221),
.Y(n_301)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_28),
.Y(n_150)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_28),
.Y(n_318)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_29),
.Y(n_263)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_34),
.A2(n_178),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_35),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_35),
.Y(n_323)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_36),
.Y(n_156)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_38),
.Y(n_262)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_40),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_43),
.A2(n_75),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_43),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_43),
.B(n_312),
.Y(n_311)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_43),
.A2(n_175),
.B(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_43),
.B(n_128),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21x1_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_52),
.B(n_64),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_62),
.Y(n_109)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_74),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_104),
.Y(n_78)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_79),
.Y(n_242)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_86),
.B1(n_100),
.B2(n_103),
.Y(n_79)
);

OA21x2_ASAP7_75t_L g209 ( 
.A1(n_80),
.A2(n_103),
.B(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_87),
.B(n_101),
.Y(n_210)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_104),
.B(n_239),
.C(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_104),
.B(n_259),
.C(n_260),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_104),
.A2(n_105),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_113),
.B1(n_128),
.B2(n_138),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22x1_ASAP7_75t_L g205 ( 
.A1(n_107),
.A2(n_114),
.B1(n_139),
.B2(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_113),
.A2(n_128),
.B(n_138),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_128),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_122),
.B2(n_124),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_127),
.Y(n_293)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_136),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_131),
.Y(n_299)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_197),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_144),
.B(n_197),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_144),
.B(n_198),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_158),
.B2(n_196),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_146),
.B(n_158),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_156),
.B(n_157),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_147),
.A2(n_221),
.B1(n_222),
.B2(n_226),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g261 ( 
.A1(n_157),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

OAI211xp5_ASAP7_75t_L g274 ( 
.A1(n_157),
.A2(n_259),
.B(n_262),
.C(n_263),
.Y(n_274)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_158),
.B(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_158),
.A2(n_196),
.B1(n_310),
.B2(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_158),
.A2(n_196),
.B1(n_205),
.B2(n_253),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_158),
.B(n_253),
.C(n_347),
.Y(n_351)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22x1_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_170),
.B1(n_186),
.B2(n_195),
.Y(n_159)
);

AOI22x1_ASAP7_75t_L g217 ( 
.A1(n_160),
.A2(n_170),
.B1(n_195),
.B2(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_165),
.Y(n_285)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_175),
.B(n_180),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_177),
.Y(n_314)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_201),
.C(n_202),
.Y(n_200)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_182),
.Y(n_338)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.C(n_207),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_205),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_209),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_238),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_233),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_271),
.C(n_275),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_216),
.A2(n_217),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_216),
.A2(n_275),
.B1(n_276),
.B2(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_217),
.Y(n_354)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_266),
.B(n_357),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_264),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_248),
.B(n_264),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_255),
.C(n_257),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_249),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_261),
.B(n_274),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_260),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_260),
.B(n_330),
.Y(n_342)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_261),
.B(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21x1_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_305),
.B(n_356),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_302),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_270),
.B(n_302),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_271),
.B(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_300),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_277),
.B(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

BUFx4f_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI21x1_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_350),
.B(n_355),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_344),
.B(n_349),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_328),
.B(n_343),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_324),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_SL g343 ( 
.A(n_309),
.B(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_315),
.B(n_319),
.Y(n_310)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI21x1_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_332),
.B(n_342),
.Y(n_328)
);

AOI21x1_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_339),
.B(n_341),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_345),
.B(n_346),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_352),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);


endmodule