module real_aes_8517_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_0), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g444 ( .A(n_0), .Y(n_444) );
INVx1_ASAP7_75t_L g529 ( .A(n_1), .Y(n_529) );
INVx1_ASAP7_75t_L g193 ( .A(n_2), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_3), .A2(n_38), .B1(n_155), .B2(n_471), .Y(n_488) );
AOI21xp33_ASAP7_75t_L g134 ( .A1(n_4), .A2(n_135), .B(n_142), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_5), .B(n_128), .Y(n_520) );
AND2x6_ASAP7_75t_L g140 ( .A(n_6), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_7), .A2(n_234), .B(n_235), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_8), .B(n_39), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_8), .B(n_39), .Y(n_445) );
INVx1_ASAP7_75t_L g152 ( .A(n_9), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_10), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g133 ( .A(n_11), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_12), .B(n_165), .Y(n_466) );
INVx1_ASAP7_75t_L g240 ( .A(n_13), .Y(n_240) );
INVx1_ASAP7_75t_L g524 ( .A(n_14), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_15), .B(n_129), .Y(n_505) );
AO32x2_ASAP7_75t_L g486 ( .A1(n_16), .A2(n_128), .A3(n_162), .B1(n_487), .B2(n_491), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_17), .B(n_155), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_18), .B(n_181), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_19), .B(n_129), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_20), .A2(n_49), .B1(n_155), .B2(n_471), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_21), .B(n_135), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_22), .A2(n_75), .B1(n_155), .B2(n_165), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_23), .B(n_155), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_24), .B(n_126), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_25), .A2(n_238), .B(n_239), .C(n_241), .Y(n_237) );
OAI222xp33_ASAP7_75t_L g450 ( .A1(n_26), .A2(n_451), .B1(n_738), .B2(n_744), .C1(n_745), .C2(n_747), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_26), .Y(n_744) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_28), .B(n_158), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_29), .B(n_150), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_30), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_31), .Y(n_747) );
INVx1_ASAP7_75t_L g171 ( .A(n_32), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_33), .B(n_158), .Y(n_484) );
INVx2_ASAP7_75t_L g138 ( .A(n_34), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_35), .B(n_155), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_36), .B(n_158), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_37), .A2(n_140), .B(n_145), .C(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g169 ( .A(n_40), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_41), .B(n_150), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_42), .B(n_155), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_43), .A2(n_85), .B1(n_212), .B2(n_471), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_44), .B(n_155), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_45), .B(n_155), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_46), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_47), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_48), .B(n_135), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_50), .A2(n_59), .B1(n_155), .B2(n_165), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_51), .A2(n_145), .B1(n_165), .B2(n_167), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_52), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_53), .B(n_155), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_54), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_55), .B(n_155), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_56), .A2(n_149), .B(n_151), .C(n_154), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_57), .Y(n_258) );
INVx1_ASAP7_75t_L g143 ( .A(n_58), .Y(n_143) );
INVx1_ASAP7_75t_L g141 ( .A(n_60), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_61), .A2(n_116), .B1(n_117), .B2(n_436), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_61), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_62), .B(n_155), .Y(n_530) );
INVx1_ASAP7_75t_L g132 ( .A(n_63), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_64), .Y(n_113) );
AO32x2_ASAP7_75t_L g496 ( .A1(n_65), .A2(n_128), .A3(n_220), .B1(n_491), .B2(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g541 ( .A(n_66), .Y(n_541) );
INVx1_ASAP7_75t_L g479 ( .A(n_67), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_SL g180 ( .A1(n_68), .A2(n_154), .B(n_181), .C(n_182), .Y(n_180) );
INVxp67_ASAP7_75t_L g183 ( .A(n_69), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_70), .B(n_165), .Y(n_480) );
INVx1_ASAP7_75t_L g108 ( .A(n_71), .Y(n_108) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_72), .A2(n_100), .B1(n_109), .B2(n_751), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_73), .Y(n_175) );
INVx1_ASAP7_75t_L g251 ( .A(n_74), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_76), .A2(n_140), .B(n_145), .C(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_77), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_78), .B(n_165), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_79), .B(n_194), .Y(n_208) );
INVx2_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_81), .B(n_181), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_82), .B(n_165), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_83), .A2(n_140), .B(n_145), .C(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g105 ( .A(n_84), .Y(n_105) );
OR2x2_ASAP7_75t_L g441 ( .A(n_84), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g453 ( .A(n_84), .B(n_443), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_86), .A2(n_98), .B1(n_165), .B2(n_166), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_87), .B(n_158), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_88), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_89), .A2(n_140), .B(n_145), .C(n_223), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_90), .Y(n_230) );
INVx1_ASAP7_75t_L g179 ( .A(n_91), .Y(n_179) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_92), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_93), .B(n_194), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_94), .B(n_165), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_95), .B(n_128), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_96), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_97), .A2(n_135), .B(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g752 ( .A(n_101), .Y(n_752) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
OR2x2_ASAP7_75t_L g455 ( .A(n_105), .B(n_443), .Y(n_455) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_105), .B(n_442), .Y(n_746) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OAI21xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_449), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g750 ( .A(n_112), .Y(n_750) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_438), .B(n_446), .Y(n_114) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_119), .A2(n_452), .B1(n_454), .B2(n_456), .Y(n_451) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g437 ( .A(n_120), .Y(n_437) );
AND3x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_358), .C(n_403), .Y(n_120) );
NOR4xp25_ASAP7_75t_L g121 ( .A(n_122), .B(n_281), .C(n_322), .D(n_339), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_185), .B(n_201), .C(n_243), .Y(n_122) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_159), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_124), .B(n_186), .Y(n_185) );
NOR4xp25_ASAP7_75t_L g305 ( .A(n_124), .B(n_299), .C(n_306), .D(n_312), .Y(n_305) );
AND2x2_ASAP7_75t_L g378 ( .A(n_124), .B(n_267), .Y(n_378) );
AND2x2_ASAP7_75t_L g397 ( .A(n_124), .B(n_343), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_124), .B(n_392), .Y(n_406) );
AND2x2_ASAP7_75t_L g419 ( .A(n_124), .B(n_200), .Y(n_419) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g264 ( .A(n_125), .Y(n_264) );
AND2x2_ASAP7_75t_L g271 ( .A(n_125), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g321 ( .A(n_125), .B(n_160), .Y(n_321) );
AND2x2_ASAP7_75t_SL g332 ( .A(n_125), .B(n_267), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_125), .B(n_160), .Y(n_336) );
AND2x2_ASAP7_75t_L g345 ( .A(n_125), .B(n_270), .Y(n_345) );
BUFx2_ASAP7_75t_L g368 ( .A(n_125), .Y(n_368) );
AND2x2_ASAP7_75t_L g372 ( .A(n_125), .B(n_176), .Y(n_372) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_134), .B(n_157), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_127), .B(n_215), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_127), .B(n_491), .C(n_507), .Y(n_506) );
AO21x1_ASAP7_75t_L g544 ( .A1(n_127), .A2(n_507), .B(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_128), .A2(n_177), .B(n_184), .Y(n_176) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_128), .A2(n_512), .B(n_520), .Y(n_511) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_130), .B(n_131), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx2_ASAP7_75t_L g234 ( .A(n_135), .Y(n_234) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_136), .B(n_140), .Y(n_173) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g519 ( .A(n_137), .Y(n_519) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
INVx1_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
INVx1_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_139), .Y(n_153) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx4_ASAP7_75t_SL g156 ( .A(n_140), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_140), .A2(n_464), .B(n_468), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_140), .A2(n_478), .B(n_481), .Y(n_477) );
BUFx3_ASAP7_75t_L g491 ( .A(n_140), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_140), .A2(n_513), .B(n_516), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_140), .A2(n_523), .B(n_527), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_148), .C(n_156), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_144), .A2(n_156), .B(n_179), .C(n_180), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_144), .A2(n_156), .B(n_236), .C(n_237), .Y(n_235) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
BUFx3_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
INVx1_ASAP7_75t_L g471 ( .A(n_146), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_149), .A2(n_469), .B(n_470), .Y(n_468) );
O2A1O1Ixp5_ASAP7_75t_L g540 ( .A1(n_149), .A2(n_528), .B(n_541), .C(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g226 ( .A(n_150), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_150), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_487) );
OAI22xp5_ASAP7_75t_SL g497 ( .A1(n_150), .A2(n_153), .B1(n_498), .B2(n_499), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_150), .A2(n_489), .B1(n_508), .B2(n_509), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_153), .B(n_183), .Y(n_182) );
INVx5_ASAP7_75t_L g194 ( .A(n_153), .Y(n_194) );
O2A1O1Ixp5_ASAP7_75t_SL g478 ( .A1(n_154), .A2(n_194), .B(n_479), .C(n_480), .Y(n_478) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_155), .Y(n_227) );
OAI22xp33_ASAP7_75t_L g163 ( .A1(n_156), .A2(n_164), .B1(n_172), .B2(n_173), .Y(n_163) );
INVx1_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
INVx2_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_158), .A2(n_233), .B(n_242), .Y(n_232) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_158), .A2(n_463), .B(n_472), .Y(n_462) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_158), .A2(n_477), .B(n_484), .Y(n_476) );
OR2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_176), .Y(n_159) );
AND2x2_ASAP7_75t_L g200 ( .A(n_160), .B(n_176), .Y(n_200) );
BUFx2_ASAP7_75t_L g274 ( .A(n_160), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_160), .A2(n_307), .B1(n_309), .B2(n_310), .Y(n_306) );
OR2x2_ASAP7_75t_L g328 ( .A(n_160), .B(n_188), .Y(n_328) );
AND2x2_ASAP7_75t_L g392 ( .A(n_160), .B(n_270), .Y(n_392) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g260 ( .A(n_161), .B(n_188), .Y(n_260) );
AND2x2_ASAP7_75t_L g267 ( .A(n_161), .B(n_176), .Y(n_267) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_161), .Y(n_309) );
OR2x2_ASAP7_75t_L g344 ( .A(n_161), .B(n_187), .Y(n_344) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_174), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_162), .B(n_175), .Y(n_174) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_162), .A2(n_189), .B(n_197), .Y(n_188) );
INVx2_ASAP7_75t_L g213 ( .A(n_162), .Y(n_213) );
INVx2_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_167) );
INVx2_ASAP7_75t_L g170 ( .A(n_168), .Y(n_170) );
INVx4_ASAP7_75t_L g238 ( .A(n_168), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_173), .A2(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_173), .A2(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g263 ( .A(n_176), .Y(n_263) );
INVx3_ASAP7_75t_L g272 ( .A(n_176), .Y(n_272) );
BUFx2_ASAP7_75t_L g296 ( .A(n_176), .Y(n_296) );
AND2x2_ASAP7_75t_L g329 ( .A(n_176), .B(n_264), .Y(n_329) );
INVx1_ASAP7_75t_L g467 ( .A(n_181), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_185), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_414) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_200), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_187), .B(n_272), .Y(n_276) );
INVx1_ASAP7_75t_L g304 ( .A(n_187), .Y(n_304) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g270 ( .A(n_188), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .C(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g489 ( .A(n_194), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_194), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_194), .A2(n_538), .B(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_196), .A2(n_524), .B(n_525), .C(n_526), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_199), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_199), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
NAND2x1_ASAP7_75t_SL g201 ( .A(n_202), .B(n_216), .Y(n_201) );
AND2x2_ASAP7_75t_L g280 ( .A(n_202), .B(n_231), .Y(n_280) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_202), .Y(n_354) );
AND2x2_ASAP7_75t_L g381 ( .A(n_202), .B(n_301), .Y(n_381) );
AND2x2_ASAP7_75t_L g389 ( .A(n_202), .B(n_351), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_202), .B(n_246), .Y(n_416) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g247 ( .A(n_203), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g265 ( .A(n_203), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g286 ( .A(n_203), .Y(n_286) );
INVx1_ASAP7_75t_L g292 ( .A(n_203), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_203), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g325 ( .A(n_203), .B(n_249), .Y(n_325) );
OR2x2_ASAP7_75t_L g363 ( .A(n_203), .B(n_318), .Y(n_363) );
AOI32xp33_ASAP7_75t_L g375 ( .A1(n_203), .A2(n_376), .A3(n_379), .B1(n_380), .B2(n_381), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_203), .B(n_351), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_203), .B(n_311), .Y(n_426) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_206), .B(n_213), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_210), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g241 ( .A(n_212), .Y(n_241) );
INVx1_ASAP7_75t_L g256 ( .A(n_213), .Y(n_256) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_213), .A2(n_522), .B(n_531), .Y(n_521) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_213), .A2(n_536), .B(n_543), .Y(n_535) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g337 ( .A(n_217), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
INVx1_ASAP7_75t_L g299 ( .A(n_218), .Y(n_299) );
AND2x2_ASAP7_75t_L g301 ( .A(n_218), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_218), .B(n_248), .Y(n_318) );
AND2x2_ASAP7_75t_L g351 ( .A(n_218), .B(n_327), .Y(n_351) );
AND2x2_ASAP7_75t_L g388 ( .A(n_218), .B(n_249), .Y(n_388) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g246 ( .A(n_219), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_219), .B(n_248), .Y(n_278) );
AND2x2_ASAP7_75t_L g285 ( .A(n_219), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g326 ( .A(n_219), .B(n_327), .Y(n_326) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_229), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_228), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_227), .Y(n_223) );
INVx2_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_231), .B(n_248), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_231), .B(n_293), .Y(n_374) );
INVx1_ASAP7_75t_L g396 ( .A(n_231), .Y(n_396) );
INVx1_ASAP7_75t_L g413 ( .A(n_231), .Y(n_413) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g266 ( .A(n_232), .B(n_248), .Y(n_266) );
AND2x2_ASAP7_75t_L g288 ( .A(n_232), .B(n_249), .Y(n_288) );
INVx1_ASAP7_75t_L g327 ( .A(n_232), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_238), .B(n_240), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_238), .A2(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g526 ( .A(n_238), .Y(n_526) );
AOI221x1_ASAP7_75t_SL g243 ( .A1(n_244), .A2(n_259), .B1(n_265), .B2(n_267), .C(n_268), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_244), .A2(n_332), .B1(n_399), .B2(n_400), .Y(n_398) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
AND2x2_ASAP7_75t_L g290 ( .A(n_245), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g385 ( .A(n_245), .B(n_265), .Y(n_385) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g341 ( .A(n_246), .B(n_266), .Y(n_341) );
INVx1_ASAP7_75t_L g353 ( .A(n_247), .Y(n_353) );
AND2x2_ASAP7_75t_L g364 ( .A(n_247), .B(n_351), .Y(n_364) );
AND2x2_ASAP7_75t_L g431 ( .A(n_247), .B(n_326), .Y(n_431) );
INVx2_ASAP7_75t_L g293 ( .A(n_248), .Y(n_293) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_256), .B(n_257), .Y(n_249) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_260), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g383 ( .A(n_260), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_261), .B(n_344), .Y(n_347) );
INVx3_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_262), .A2(n_383), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_SL g405 ( .A(n_265), .B(n_291), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_266), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g357 ( .A(n_266), .B(n_285), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_266), .B(n_292), .Y(n_434) );
AND2x2_ASAP7_75t_L g303 ( .A(n_267), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g370 ( .A(n_267), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .B(n_277), .Y(n_268) );
NAND2x1_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_270), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g319 ( .A(n_270), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g331 ( .A(n_270), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_270), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g355 ( .A(n_271), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_271), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_271), .B(n_274), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AOI211xp5_ASAP7_75t_L g342 ( .A1(n_274), .A2(n_313), .B(n_343), .C(n_345), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_274), .A2(n_361), .B1(n_364), .B2(n_365), .C(n_369), .Y(n_360) );
AND2x2_ASAP7_75t_L g356 ( .A(n_275), .B(n_309), .Y(n_356) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g316 ( .A(n_280), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g387 ( .A(n_280), .B(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_289), .C(n_314), .Y(n_281) );
NAND3xp33_ASAP7_75t_SL g400 ( .A(n_282), .B(n_401), .C(n_402), .Y(n_400) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
OR2x2_ASAP7_75t_L g373 ( .A(n_284), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_294), .B1(n_297), .B2(n_303), .C(n_305), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_291), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_291), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_296), .A2(n_353), .B1(n_354), .B2(n_355), .Y(n_352) );
OR2x2_ASAP7_75t_L g433 ( .A(n_296), .B(n_344), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVxp67_ASAP7_75t_L g407 ( .A(n_299), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_301), .B(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g308 ( .A(n_302), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_304), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_304), .B(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_304), .B(n_371), .Y(n_410) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_308), .Y(n_334) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g424 ( .A(n_313), .B(n_344), .Y(n_424) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g402 ( .A(n_319), .Y(n_402) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI322xp33_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_328), .A3(n_329), .B1(n_330), .B2(n_333), .C1(n_335), .C2(n_337), .Y(n_322) );
OAI322xp33_ASAP7_75t_L g404 ( .A1(n_323), .A2(n_405), .A3(n_406), .B1(n_407), .B2(n_408), .C1(n_409), .C2(n_411), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx4_ASAP7_75t_L g338 ( .A(n_325), .Y(n_338) );
AND2x2_ASAP7_75t_L g399 ( .A(n_325), .B(n_351), .Y(n_399) );
AND2x2_ASAP7_75t_L g412 ( .A(n_325), .B(n_413), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_328), .Y(n_423) );
INVx1_ASAP7_75t_L g401 ( .A(n_329), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OR2x2_ASAP7_75t_L g335 ( .A(n_331), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g418 ( .A(n_331), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_331), .B(n_372), .Y(n_429) );
OR2x2_ASAP7_75t_L g362 ( .A(n_334), .B(n_363), .Y(n_362) );
INVxp33_ASAP7_75t_L g379 ( .A(n_334), .Y(n_379) );
OAI221xp5_ASAP7_75t_SL g339 ( .A1(n_338), .A2(n_340), .B1(n_342), .B2(n_346), .C(n_348), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_338), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g422 ( .A(n_338), .Y(n_422) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
INVx3_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AOI322xp5_ASAP7_75t_L g386 ( .A1(n_345), .A2(n_370), .A3(n_387), .B1(n_389), .B2(n_390), .C1(n_393), .C2(n_397), .Y(n_386) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B1(n_356), .B2(n_357), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_382), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_360), .B(n_375), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_363), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_366), .B(n_377), .Y(n_380) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
OAI322xp33_ASAP7_75t_L g420 ( .A1(n_368), .A2(n_421), .A3(n_423), .B1(n_424), .B2(n_425), .C1(n_427), .C2(n_430), .Y(n_420) );
AOI21xp33_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_371), .B(n_373), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_378), .B(n_426), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_384), .B(n_386), .C(n_398), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NOR4xp25_ASAP7_75t_L g403 ( .A(n_404), .B(n_414), .C(n_420), .D(n_432), .Y(n_403) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
CKINVDCx14_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_434), .B(n_435), .Y(n_432) );
BUFx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_437), .A2(n_739), .B1(n_742), .B2(n_743), .Y(n_738) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g447 ( .A(n_441), .Y(n_447) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_446), .A2(n_450), .B(n_748), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g741 ( .A(n_453), .Y(n_741) );
INVx6_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g742 ( .A(n_455), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_456), .Y(n_743) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_660), .Y(n_456) );
NAND5xp2_ASAP7_75t_L g457 ( .A(n_458), .B(n_579), .C(n_594), .D(n_620), .E(n_642), .Y(n_457) );
NOR2xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_559), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_500), .B1(n_532), .B2(n_548), .C(n_549), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_492), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_461), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g736 ( .A(n_461), .Y(n_736) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
INVx1_ASAP7_75t_L g576 ( .A(n_462), .Y(n_576) );
AND2x2_ASAP7_75t_L g578 ( .A(n_462), .B(n_486), .Y(n_578) );
AND2x2_ASAP7_75t_L g588 ( .A(n_462), .B(n_485), .Y(n_588) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_462), .Y(n_606) );
INVx1_ASAP7_75t_L g616 ( .A(n_462), .Y(n_616) );
OR2x2_ASAP7_75t_L g654 ( .A(n_462), .B(n_553), .Y(n_654) );
INVx2_ASAP7_75t_L g704 ( .A(n_462), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_462), .B(n_552), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_467), .Y(n_464) );
NOR2xp67_ASAP7_75t_L g473 ( .A(n_474), .B(n_485), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_475), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_475), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_475), .B(n_576), .Y(n_636) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_476), .Y(n_494) );
INVx2_ASAP7_75t_L g553 ( .A(n_476), .Y(n_553) );
OR2x2_ASAP7_75t_L g615 ( .A(n_476), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g554 ( .A(n_485), .B(n_496), .Y(n_554) );
AND2x2_ASAP7_75t_L g571 ( .A(n_485), .B(n_551), .Y(n_571) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g495 ( .A(n_486), .B(n_496), .Y(n_495) );
BUFx2_ASAP7_75t_L g574 ( .A(n_486), .Y(n_574) );
AND2x2_ASAP7_75t_L g703 ( .A(n_486), .B(n_704), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_489), .A2(n_517), .B(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_489), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_491), .A2(n_537), .B(n_540), .Y(n_536) );
INVx1_ASAP7_75t_L g548 ( .A(n_492), .Y(n_548) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x2_ASAP7_75t_L g666 ( .A(n_493), .B(n_554), .Y(n_666) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g667 ( .A(n_494), .B(n_578), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_495), .A2(n_635), .B(n_637), .C(n_639), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_495), .B(n_635), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_495), .A2(n_565), .B1(n_708), .B2(n_709), .C(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g551 ( .A(n_496), .Y(n_551) );
INVx1_ASAP7_75t_L g587 ( .A(n_496), .Y(n_587) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_496), .Y(n_596) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
AND2x2_ASAP7_75t_L g613 ( .A(n_502), .B(n_558), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_502), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_503), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g705 ( .A(n_503), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g737 ( .A(n_503), .Y(n_737) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g567 ( .A(n_504), .Y(n_567) );
AND2x2_ASAP7_75t_L g593 ( .A(n_504), .B(n_547), .Y(n_593) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_504), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g609 ( .A(n_504), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g545 ( .A(n_505), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_510), .B(n_649), .Y(n_684) );
INVx1_ASAP7_75t_SL g688 ( .A(n_510), .Y(n_688) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
INVx3_ASAP7_75t_L g547 ( .A(n_511), .Y(n_547) );
AND2x2_ASAP7_75t_L g558 ( .A(n_511), .B(n_535), .Y(n_558) );
AND2x2_ASAP7_75t_L g580 ( .A(n_511), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g625 ( .A(n_511), .B(n_619), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_511), .B(n_557), .Y(n_706) );
INVx2_ASAP7_75t_L g528 ( .A(n_519), .Y(n_528) );
AND2x2_ASAP7_75t_L g546 ( .A(n_521), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g557 ( .A(n_521), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_521), .B(n_535), .Y(n_582) );
AND2x2_ASAP7_75t_L g618 ( .A(n_521), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_546), .Y(n_533) );
INVx1_ASAP7_75t_L g598 ( .A(n_534), .Y(n_598) );
AND2x2_ASAP7_75t_L g640 ( .A(n_534), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_534), .B(n_561), .Y(n_646) );
AOI21xp5_ASAP7_75t_SL g720 ( .A1(n_534), .A2(n_552), .B(n_575), .Y(n_720) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
OR2x2_ASAP7_75t_L g563 ( .A(n_535), .B(n_544), .Y(n_563) );
AND2x2_ASAP7_75t_L g610 ( .A(n_535), .B(n_547), .Y(n_610) );
INVx2_ASAP7_75t_L g619 ( .A(n_535), .Y(n_619) );
INVx1_ASAP7_75t_L g725 ( .A(n_535), .Y(n_725) );
AND2x2_ASAP7_75t_L g649 ( .A(n_544), .B(n_619), .Y(n_649) );
INVx1_ASAP7_75t_L g674 ( .A(n_544), .Y(n_674) );
AND2x2_ASAP7_75t_L g583 ( .A(n_546), .B(n_567), .Y(n_583) );
AND2x2_ASAP7_75t_L g595 ( .A(n_546), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_SL g713 ( .A(n_546), .Y(n_713) );
INVx2_ASAP7_75t_L g603 ( .A(n_547), .Y(n_603) );
AND2x2_ASAP7_75t_L g641 ( .A(n_547), .B(n_557), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_547), .B(n_725), .Y(n_724) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_554), .B(n_555), .Y(n_549) );
AND2x2_ASAP7_75t_L g656 ( .A(n_550), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g710 ( .A(n_550), .Y(n_710) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g630 ( .A(n_551), .Y(n_630) );
BUFx2_ASAP7_75t_L g729 ( .A(n_551), .Y(n_729) );
BUFx2_ASAP7_75t_L g600 ( .A(n_552), .Y(n_600) );
AND2x2_ASAP7_75t_L g702 ( .A(n_552), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g685 ( .A(n_553), .Y(n_685) );
AND2x4_ASAP7_75t_L g612 ( .A(n_554), .B(n_575), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_554), .B(n_636), .Y(n_648) );
AOI32xp33_ASAP7_75t_L g572 ( .A1(n_555), .A2(n_573), .A3(n_575), .B1(n_577), .B2(n_578), .Y(n_572) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx3_ASAP7_75t_L g561 ( .A(n_556), .Y(n_561) );
OR2x2_ASAP7_75t_L g697 ( .A(n_556), .B(n_653), .Y(n_697) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g566 ( .A(n_557), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g673 ( .A(n_557), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g565 ( .A(n_558), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g577 ( .A(n_558), .B(n_567), .Y(n_577) );
INVx1_ASAP7_75t_L g698 ( .A(n_558), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_558), .B(n_673), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_564), .B(n_568), .C(n_572), .Y(n_559) );
OAI322xp33_ASAP7_75t_L g668 ( .A1(n_560), .A2(n_605), .A3(n_669), .B1(n_671), .B2(n_675), .C1(n_676), .C2(n_680), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVxp67_ASAP7_75t_L g633 ( .A(n_561), .Y(n_633) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g687 ( .A(n_563), .B(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_563), .B(n_603), .Y(n_734) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g626 ( .A(n_566), .Y(n_626) );
OR2x2_ASAP7_75t_L g712 ( .A(n_567), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_570), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g621 ( .A(n_571), .B(n_600), .Y(n_621) );
AND2x2_ASAP7_75t_L g692 ( .A(n_571), .B(n_605), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_571), .B(n_679), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_573), .A2(n_580), .B1(n_583), .B2(n_584), .C(n_589), .Y(n_579) );
OR2x2_ASAP7_75t_L g590 ( .A(n_573), .B(n_586), .Y(n_590) );
AND2x2_ASAP7_75t_L g678 ( .A(n_573), .B(n_679), .Y(n_678) );
AOI32xp33_ASAP7_75t_L g717 ( .A1(n_573), .A2(n_603), .A3(n_718), .B1(n_719), .B2(n_722), .Y(n_717) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_574), .B(n_610), .C(n_633), .Y(n_651) );
AND2x2_ASAP7_75t_L g677 ( .A(n_574), .B(n_670), .Y(n_677) );
INVxp67_ASAP7_75t_L g657 ( .A(n_575), .Y(n_657) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_578), .B(n_630), .Y(n_686) );
INVx2_ASAP7_75t_L g696 ( .A(n_578), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_578), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g665 ( .A(n_581), .Y(n_665) );
OR2x2_ASAP7_75t_L g591 ( .A(n_582), .B(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_584), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_587), .Y(n_670) );
AND2x2_ASAP7_75t_L g629 ( .A(n_588), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g675 ( .A(n_588), .Y(n_675) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_588), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AOI21xp33_ASAP7_75t_SL g614 ( .A1(n_590), .A2(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g708 ( .A(n_593), .B(n_618), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B(n_607), .C(n_614), .Y(n_594) );
AND2x2_ASAP7_75t_L g638 ( .A(n_596), .B(n_606), .Y(n_638) );
INVx2_ASAP7_75t_L g653 ( .A(n_596), .Y(n_653) );
OR2x2_ASAP7_75t_L g691 ( .A(n_596), .B(n_654), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_596), .B(n_734), .Y(n_733) );
AOI211xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_599), .B(n_601), .C(n_604), .Y(n_597) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_600), .B(n_638), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g719 ( .A1(n_601), .A2(n_696), .B(n_720), .C(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_602), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g659 ( .A(n_603), .B(n_649), .Y(n_659) );
INVx1_ASAP7_75t_L g664 ( .A(n_603), .Y(n_664) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_611), .Y(n_607) );
INVxp33_ASAP7_75t_L g715 ( .A(n_609), .Y(n_715) );
AND2x2_ASAP7_75t_L g694 ( .A(n_610), .B(n_673), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_615), .A2(n_677), .B(n_678), .Y(n_676) );
OAI322xp33_ASAP7_75t_L g695 ( .A1(n_617), .A2(n_696), .A3(n_697), .B1(n_698), .B2(n_699), .C1(n_701), .C2(n_705), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_627), .B2(n_631), .C(n_634), .Y(n_620) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g672 ( .A(n_625), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g716 ( .A(n_629), .Y(n_716) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_632), .B(n_652), .Y(n_718) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g681 ( .A(n_641), .B(n_649), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_647), .B2(n_649), .C(n_650), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_645), .A2(n_662), .B1(n_666), .B2(n_667), .C(n_668), .Y(n_661) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_649), .B(n_664), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_655), .B2(n_658), .Y(n_650) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx2_ASAP7_75t_SL g679 ( .A(n_654), .Y(n_679) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND5xp2_ASAP7_75t_L g660 ( .A(n_661), .B(n_682), .C(n_707), .D(n_717), .E(n_727), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_665), .Y(n_662) );
NOR4xp25_ASAP7_75t_L g735 ( .A(n_664), .B(n_670), .C(n_736), .D(n_737), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_667), .A2(n_728), .B1(n_730), .B2(n_732), .C(n_735), .Y(n_727) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g726 ( .A(n_673), .Y(n_726) );
OAI322xp33_ASAP7_75t_L g683 ( .A1(n_677), .A2(n_684), .A3(n_685), .B1(n_686), .B2(n_687), .C1(n_689), .C2(n_693), .Y(n_683) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_695), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g728 ( .A(n_703), .B(n_729), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_711) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVxp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
endmodule