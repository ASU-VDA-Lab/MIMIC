module fake_jpeg_18197_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_12),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_33),
.B1(n_23),
.B2(n_25),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_38),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_40),
.B1(n_17),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_59),
.B1(n_35),
.B2(n_43),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_23),
.B1(n_34),
.B2(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_18),
.B1(n_30),
.B2(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_36),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_23),
.B1(n_32),
.B2(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_66),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_37),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_70),
.B(n_75),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_77),
.Y(n_130)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_37),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_42),
.B1(n_35),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_96),
.B1(n_51),
.B2(n_49),
.Y(n_116)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_37),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_20),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_31),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_42),
.B1(n_31),
.B2(n_32),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_94),
.B1(n_43),
.B2(n_17),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_28),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_28),
.B1(n_27),
.B2(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_97),
.B(n_99),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_43),
.B1(n_26),
.B2(n_19),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_44),
.B(n_27),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_44),
.A2(n_19),
.B(n_26),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_70),
.B(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_49),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_16),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_112),
.C(n_41),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_108),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_41),
.C(n_36),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_63),
.B(n_16),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_51),
.B1(n_49),
.B2(n_43),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_41),
.C(n_36),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_36),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_51),
.B1(n_49),
.B2(n_41),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_133),
.B(n_141),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_125),
.B(n_130),
.C(n_124),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_145),
.B(n_160),
.Y(n_167)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_87),
.B1(n_78),
.B2(n_61),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_142),
.B1(n_151),
.B2(n_118),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_78),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_117),
.A2(n_92),
.B1(n_100),
.B2(n_51),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_109),
.B(n_26),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_0),
.B(n_1),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_128),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_60),
.B1(n_93),
.B2(n_80),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_153),
.B1(n_128),
.B2(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_109),
.B(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_149),
.B(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_152),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_80),
.B1(n_60),
.B2(n_68),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_65),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_90),
.B1(n_69),
.B2(n_74),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_97),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_134),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_157),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_161),
.Y(n_163)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_122),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_97),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_107),
.C(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_170),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_165),
.A2(n_173),
.B1(n_183),
.B2(n_184),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_133),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_123),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_160),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_129),
.B(n_123),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_185),
.B(n_189),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_106),
.B1(n_126),
.B2(n_113),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_140),
.B(n_145),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_174),
.A2(n_182),
.B(n_30),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_108),
.C(n_110),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_192),
.C(n_157),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_115),
.B1(n_110),
.B2(n_102),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_105),
.B(n_120),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_132),
.B1(n_72),
.B2(n_43),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_132),
.B1(n_41),
.B2(n_67),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_22),
.B(n_16),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_67),
.B1(n_11),
.B2(n_12),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_22),
.B(n_1),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_36),
.B1(n_15),
.B2(n_14),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_191),
.A2(n_193),
.B1(n_0),
.B2(n_2),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_137),
.C(n_147),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_13),
.B1(n_11),
.B2(n_2),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_160),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_221),
.B(n_166),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_197),
.B(n_217),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_206),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_211),
.C(n_215),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_154),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_204),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_138),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_202),
.B(n_208),
.Y(n_231)
);

AOI21x1_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_159),
.B(n_138),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_207),
.B(n_219),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_171),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_190),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_167),
.C(n_194),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_30),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_192),
.C(n_169),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_216),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_30),
.C(n_21),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_21),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_21),
.C(n_18),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_18),
.C(n_1),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_3),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_185),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_162),
.B(n_0),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_164),
.B1(n_177),
.B2(n_180),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_182),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_223),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_179),
.B1(n_195),
.B2(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_170),
.B1(n_184),
.B2(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_243),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_165),
.B1(n_173),
.B2(n_180),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_241),
.B1(n_214),
.B2(n_222),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_214),
.A2(n_162),
.B1(n_183),
.B2(n_166),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_189),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_196),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_205),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_260),
.Y(n_270)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_239),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_204),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_231),
.B(n_211),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_200),
.C(n_201),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_261),
.C(n_238),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_197),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_176),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_257),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

AO221x1_ASAP7_75t_L g268 ( 
.A1(n_258),
.A2(n_228),
.B1(n_235),
.B2(n_233),
.C(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_240),
.B1(n_241),
.B2(n_237),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_227),
.B(n_215),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_205),
.C(n_217),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_264),
.B1(n_233),
.B2(n_236),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_224),
.B(n_167),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_262),
.B1(n_249),
.B2(n_265),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_272),
.C(n_279),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_247),
.B1(n_249),
.B2(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_238),
.C(n_243),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_245),
.C(n_232),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_212),
.B(n_219),
.C(n_193),
.D(n_6),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_277),
.A2(n_278),
.B1(n_281),
.B2(n_6),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_256),
.B(n_9),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_3),
.C(n_4),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_3),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_258),
.C(n_5),
.Y(n_287)
);

XOR2x1_ASAP7_75t_SL g281 ( 
.A(n_246),
.B(n_4),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_263),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_285),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_293),
.B1(n_277),
.B2(n_279),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_289),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_280),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_4),
.C(n_5),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_292),
.C(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_4),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_290),
.B(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_6),
.C(n_7),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_294),
.B(n_296),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_273),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_298),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_276),
.B(n_273),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_302),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_9),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_282),
.B(n_292),
.Y(n_304)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_288),
.C(n_287),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_308),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_299),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_307),
.C(n_294),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_301),
.B(n_296),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_312),
.B(n_305),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_314),
.B(n_310),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_309),
.B1(n_311),
.B2(n_306),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_7),
.B(n_8),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_8),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_8),
.Y(n_319)
);


endmodule