module fake_jpeg_8951_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_40),
.B(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_31),
.B(n_44),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_62),
.B(n_40),
.C(n_21),
.Y(n_79)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_22),
.B1(n_20),
.B2(n_26),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_65),
.B1(n_38),
.B2(n_33),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_64),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_22),
.B1(n_24),
.B2(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_24),
.C(n_32),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_64),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g107 ( 
.A(n_70),
.B(n_86),
.CON(n_107),
.SN(n_107)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_74),
.B1(n_23),
.B2(n_34),
.Y(n_110)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_75),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_45),
.B1(n_43),
.B2(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_20),
.B1(n_35),
.B2(n_33),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_35),
.B1(n_29),
.B2(n_26),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_79),
.B(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_83),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_88),
.B1(n_34),
.B2(n_61),
.Y(n_105)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_33),
.B(n_25),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_25),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_26),
.B1(n_35),
.B2(n_29),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_29),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_70),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_95),
.Y(n_117)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_102),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_116),
.B1(n_100),
.B2(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_108),
.B1(n_32),
.B2(n_18),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_46),
.B1(n_61),
.B2(n_17),
.Y(n_108)
);

NOR2x1p5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_120),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_94),
.B1(n_83),
.B2(n_73),
.Y(n_132)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_50),
.Y(n_114)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_23),
.B(n_90),
.C(n_36),
.D(n_32),
.Y(n_138)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_124),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_23),
.B1(n_50),
.B2(n_30),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_120),
.B(n_74),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_0),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_39),
.C(n_44),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_36),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_28),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_135),
.Y(n_163)
);

BUFx8_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_128),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_132),
.B1(n_136),
.B2(n_139),
.Y(n_156)
);

XOR2x1_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_114),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_81),
.B1(n_90),
.B2(n_95),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_140),
.B1(n_152),
.B2(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_85),
.B1(n_80),
.B2(n_87),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_113),
.B(n_18),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_32),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_87),
.B1(n_85),
.B2(n_80),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_96),
.B1(n_97),
.B2(n_75),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_147),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_149),
.B1(n_151),
.B2(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_109),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_28),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_154),
.B(n_119),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_109),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_170),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_158),
.B(n_167),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_160),
.A2(n_164),
.B(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_165),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_107),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_175),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_109),
.B(n_120),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_122),
.C(n_102),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_120),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_181),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_152),
.B1(n_132),
.B2(n_130),
.Y(n_197)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_125),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_71),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_30),
.B(n_19),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_145),
.C(n_138),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_181),
.Y(n_215)
);

AOI21x1_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_138),
.B(n_137),
.Y(n_189)
);

AOI21x1_ASAP7_75t_L g235 ( 
.A1(n_189),
.A2(n_32),
.B(n_28),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_192),
.Y(n_240)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_203),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_130),
.B1(n_135),
.B2(n_144),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_210),
.B1(n_211),
.B2(n_176),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_172),
.B(n_154),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_160),
.A2(n_144),
.B1(n_147),
.B2(n_143),
.Y(n_204)
);

OAI31xp33_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_142),
.A3(n_149),
.B(n_32),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_0),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_106),
.B1(n_125),
.B2(n_121),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_167),
.A2(n_106),
.B1(n_121),
.B2(n_89),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_184),
.A2(n_106),
.B1(n_118),
.B2(n_112),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_158),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_213),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_171),
.B1(n_165),
.B2(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_215),
.A2(n_218),
.B(n_223),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_162),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_236),
.C(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_169),
.B1(n_163),
.B2(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_202),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_198),
.A2(n_159),
.B1(n_177),
.B2(n_156),
.Y(n_219)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_156),
.B1(n_170),
.B2(n_164),
.Y(n_220)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_227),
.B1(n_229),
.B2(n_233),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_175),
.B1(n_157),
.B2(n_174),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_211),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_189),
.A2(n_178),
.B1(n_30),
.B2(n_19),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

AO21x2_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_17),
.B(n_1),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_235),
.A2(n_238),
.B1(n_239),
.B2(n_192),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_28),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_28),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_210),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_196),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_243),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_199),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_12),
.B(n_11),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_193),
.B1(n_212),
.B2(n_191),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_213),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_249),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_240),
.B1(n_233),
.B2(n_15),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_237),
.B(n_209),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_209),
.C(n_204),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_257),
.C(n_262),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_197),
.C(n_187),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_194),
.B1(n_15),
.B2(n_14),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_260),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_225),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_239),
.C(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_0),
.C(n_2),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_263),
.B(n_278),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_277),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_226),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_269),
.C(n_275),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_2),
.C(n_3),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_276),
.C(n_254),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_14),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_249),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_12),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_3),
.C(n_4),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_259),
.C(n_254),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_292),
.C(n_293),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_252),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_274),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_242),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_280),
.Y(n_297)
);

OAI221xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_242),
.B1(n_250),
.B2(n_248),
.C(n_247),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_289),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_279),
.B1(n_273),
.B2(n_251),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_3),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_257),
.C(n_11),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_11),
.C(n_10),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_269),
.A2(n_10),
.B(n_4),
.Y(n_295)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_5),
.B(n_6),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_296),
.Y(n_311)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_275),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_276),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_304),
.A2(n_307),
.B1(n_283),
.B2(n_6),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_306),
.C(n_281),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_3),
.C(n_4),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_308),
.B(n_285),
.Y(n_309)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_309),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_293),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_315),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_7),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_301),
.A2(n_304),
.B1(n_296),
.B2(n_299),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_308),
.B1(n_7),
.B2(n_8),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_282),
.C(n_288),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_5),
.Y(n_322)
);

XNOR2x1_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_297),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_324),
.B(n_326),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_321),
.A2(n_322),
.B(n_325),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_311),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_7),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_314),
.B(n_317),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_329),
.A2(n_319),
.B(n_9),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_323),
.A2(n_318),
.B(n_315),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_326),
.B(n_312),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_327),
.B(n_332),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_328),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_9),
.Y(n_337)
);


endmodule