module real_jpeg_15950_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_541),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_0),
.B(n_542),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_1),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_1),
.B(n_54),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_1),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_1),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_1),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_1),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_1),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g350 ( 
.A(n_1),
.B(n_351),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_2),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g396 ( 
.A(n_2),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_3),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_3),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_3),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_3),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_3),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_3),
.B(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_3),
.B(n_458),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_3),
.B(n_488),
.Y(n_487)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_4),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_4),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_5),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_5),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_5),
.Y(n_314)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_5),
.Y(n_360)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_6),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_7),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_7),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_7),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_7),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_161),
.Y(n_160)
);

AND2x4_ASAP7_75t_SL g193 ( 
.A(n_7),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_7),
.B(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_8),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g255 ( 
.A(n_8),
.Y(n_255)
);

BUFx4f_ASAP7_75t_L g517 ( 
.A(n_8),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_9),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_9),
.B(n_235),
.Y(n_234)
);

AOI22x1_ASAP7_75t_SL g281 ( 
.A1(n_9),
.A2(n_17),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_9),
.B(n_91),
.Y(n_355)
);

AOI31xp33_ASAP7_75t_L g391 ( 
.A1(n_9),
.A2(n_281),
.A3(n_392),
.B(n_397),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_9),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_9),
.B(n_470),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_9),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_9),
.B(n_100),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_10),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_10),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_10),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_10),
.B(n_54),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_10),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_10),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_10),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_10),
.B(n_395),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_11),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_11),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_11),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_11),
.B(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_12),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_12),
.B(n_79),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_12),
.B(n_242),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_12),
.B(n_262),
.Y(n_261)
);

AND2x4_ASAP7_75t_SL g306 ( 
.A(n_12),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_12),
.B(n_357),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_12),
.B(n_404),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_12),
.B(n_352),
.Y(n_459)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_13),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_14),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_14),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_14),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_14),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_14),
.B(n_506),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_14),
.B(n_510),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_14),
.B(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_15),
.Y(n_118)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_15),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_15),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_15),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_16),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_17),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_17),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_17),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_17),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_17),
.B(n_253),
.Y(n_252)
);

NAND2x1_ASAP7_75t_L g256 ( 
.A(n_17),
.B(n_257),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_17),
.Y(n_393)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_18),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_18),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_171),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_169),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_150),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_R g170 ( 
.A(n_23),
.B(n_150),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_113),
.C(n_127),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_24),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_74),
.C(n_96),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_26),
.B(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.C(n_58),
.Y(n_26)
);

XNOR2x2_ASAP7_75t_SL g226 ( 
.A(n_27),
.B(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_28),
.B(n_35),
.C(n_39),
.Y(n_125)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_31),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_32),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_32),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g429 ( 
.A(n_32),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_34),
.A2(n_35),
.B1(n_116),
.B2(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_35),
.B(n_116),
.C(n_120),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_37),
.Y(n_454)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_38),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_39),
.A2(n_40),
.B1(n_99),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_40),
.B(n_99),
.C(n_102),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_42),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_44),
.B(n_58),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.C(n_53),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_45),
.B(n_53),
.Y(n_187)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_47),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_48),
.Y(n_308)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_49),
.B(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_57),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_64),
.C(n_70),
.Y(n_126)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_62),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_75),
.B(n_96),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_82),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_76),
.B(n_89),
.C(n_95),
.Y(n_149)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_89),
.B1(n_90),
.B2(n_95),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.C(n_109),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_97),
.A2(n_98),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_99),
.B(n_189),
.C(n_193),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_99),
.Y(n_202)
);

AOI22x1_ASAP7_75t_L g231 ( 
.A1(n_99),
.A2(n_193),
.B1(n_202),
.B2(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_102),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_102),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_102),
.A2(n_199),
.B1(n_294),
.B2(n_344),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_105),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_106),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_107),
.B(n_109),
.Y(n_217)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_108),
.B(n_249),
.C(n_252),
.Y(n_248)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_109),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_109),
.A2(n_212),
.B1(n_215),
.B2(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_112),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_113),
.A2(n_127),
.B1(n_128),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_125),
.C(n_126),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_119),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_132),
.C(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_140),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_131),
.C(n_140),
.Y(n_168)
);

XOR2x1_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_137),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_139),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_144),
.C(n_149),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_147),
.Y(n_317)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_147),
.Y(n_400)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_168),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_163),
.B2(n_164),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_219),
.B(n_537),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_173),
.A2(n_539),
.B(n_540),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_174),
.B(n_177),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.C(n_183),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_181),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_183),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_203),
.C(n_216),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_198),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_186),
.B(n_188),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

BUFx2_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_197),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_198),
.B(n_326),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_199),
.B(n_289),
.C(n_294),
.Y(n_288)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_216),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_212),
.C(n_215),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_211),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_211),
.Y(n_246)
);

XOR2x1_ASAP7_75t_SL g245 ( 
.A(n_207),
.B(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_212),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_214),
.Y(n_305)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_217),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_271),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_268),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_222),
.B(n_268),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g371 ( 
.A(n_224),
.B(n_226),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_228),
.B(n_371),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_247),
.C(n_264),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_229),
.B(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.C(n_245),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_230),
.B(n_233),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_240),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_234),
.A2(n_240),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_234),
.Y(n_368)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_237),
.B(n_366),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_240),
.B(n_426),
.C(n_430),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_240),
.A2(n_367),
.B1(n_426),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_241),
.Y(n_367)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_245),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_247),
.B(n_265),
.Y(n_324)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_256),
.C(n_260),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_248),
.B(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_252),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_250),
.Y(n_488)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_255),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_255),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_256),
.A2(n_260),
.B1(n_261),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_260),
.A2(n_261),
.B1(n_407),
.B2(n_408),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_261),
.B(n_402),
.C(n_407),
.Y(n_401)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AO21x2_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_376),
.B(n_534),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_369),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_329),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_274),
.B(n_329),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_322),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_275),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_297),
.C(n_318),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_277),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.C(n_288),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_278),
.B(n_412),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_280),
.A2(n_281),
.B1(n_288),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_288),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_291),
.Y(n_468)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_296),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_298),
.A2(n_318),
.B1(n_319),
.B2(n_334),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_298),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_309),
.C(n_315),
.Y(n_298)
);

XOR2x2_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_364),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_304),
.C(n_306),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_300),
.A2(n_306),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_300),
.Y(n_390)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_L g480 ( 
.A(n_306),
.B(n_481),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_308),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_310),
.B(n_315),
.Y(n_364)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_313),
.Y(n_472)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_325),
.B1(n_327),
.B2(n_328),
.Y(n_322)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.C(n_338),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_331),
.A2(n_332),
.B1(n_336),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_380),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_363),
.C(n_365),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.C(n_354),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_L g435 ( 
.A(n_342),
.B(n_436),
.Y(n_435)
);

XNOR2x1_ASAP7_75t_L g436 ( 
.A(n_345),
.B(n_354),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_350),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_346),
.B(n_350),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.C(n_361),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_355),
.A2(n_356),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_355),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_356),
.A2(n_423),
.B1(n_504),
.B2(n_505),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_356),
.B(n_500),
.C(n_504),
.Y(n_524)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_361),
.B(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_365),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_369),
.A2(n_535),
.B(n_536),
.Y(n_534)
);

AND2x2_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_372),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_370),
.B(n_372),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.C(n_375),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_439),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_382),
.C(n_414),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_379),
.B(n_383),
.Y(n_533)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.C(n_410),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_384),
.B(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_411),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_391),
.C(n_401),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_391),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_389),
.B(n_467),
.C(n_469),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_402),
.B(n_449),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_403),
.B(n_406),
.Y(n_452)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_403),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_403),
.A2(n_497),
.B1(n_498),
.B2(n_512),
.Y(n_511)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_437),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_437),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.C(n_435),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_416),
.B(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_419),
.B(n_435),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_424),
.C(n_433),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_420),
.B(n_462),
.Y(n_461)
);

INVxp33_ASAP7_75t_SL g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_434),
.Y(n_462)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

XOR2x1_ASAP7_75t_L g474 ( 
.A(n_430),
.B(n_475),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.C(n_533),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_442),
.A2(n_528),
.B(n_532),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_477),
.B(n_527),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_463),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_444),
.B(n_463),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_460),
.B2(n_461),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_447),
.B(n_451),
.C(n_460),
.Y(n_529)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

MAJx2_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.C(n_455),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_452),
.B(n_453),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

AO22x1_ASAP7_75t_SL g489 ( 
.A1(n_456),
.A2(n_457),
.B1(n_459),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_459),
.Y(n_490)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_466),
.C(n_473),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_492),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_466),
.B(n_474),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_467),
.B(n_469),
.Y(n_481)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

OAI21x1_ASAP7_75t_SL g477 ( 
.A1(n_478),
.A2(n_493),
.B(n_526),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_491),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_479),
.B(n_491),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_482),
.C(n_489),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_480),
.B(n_522),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_482),
.A2(n_483),
.B1(n_489),
.B2(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_484),
.B(n_487),
.Y(n_501)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_514),
.Y(n_513)
);

AOI21x1_ASAP7_75t_SL g493 ( 
.A1(n_494),
.A2(n_520),
.B(n_525),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_495),
.A2(n_507),
.B(n_519),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_499),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_499),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_498),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_513),
.B(n_518),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_511),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_511),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

NOR2x1_ASAP7_75t_SL g525 ( 
.A(n_521),
.B(n_524),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_SL g528 ( 
.A(n_529),
.B(n_530),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_530),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);


endmodule