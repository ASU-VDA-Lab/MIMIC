module fake_jpeg_10506_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_7),
.B(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_45),
.B1(n_24),
.B2(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_25),
.B(n_8),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_42),
.B(n_17),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_52),
.B(n_68),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_54),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_31),
.B1(n_34),
.B2(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_45),
.B1(n_34),
.B2(n_32),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_18),
.B1(n_20),
.B2(n_31),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_60),
.A2(n_21),
.B1(n_22),
.B2(n_28),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_67),
.Y(n_78)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_17),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_75),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_18),
.C(n_21),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_44),
.Y(n_104)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

OR2x2_ASAP7_75t_SL g84 ( 
.A(n_60),
.B(n_49),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_108),
.B(n_109),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_92),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_97),
.B1(n_101),
.B2(n_113),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_31),
.B1(n_45),
.B2(n_29),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_91),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_96),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_29),
.B1(n_20),
.B2(n_19),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_32),
.Y(n_96)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_44),
.B1(n_38),
.B2(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_70),
.A2(n_19),
.B1(n_32),
.B2(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_114),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_54),
.B(n_38),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_44),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_28),
.B1(n_26),
.B2(n_35),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_28),
.B1(n_26),
.B2(n_35),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_119),
.A2(n_143),
.B1(n_89),
.B2(n_105),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_97),
.B(n_0),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_120),
.A2(n_27),
.B(n_33),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_78),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_132),
.Y(n_150)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_22),
.B1(n_35),
.B2(n_28),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_81),
.B1(n_99),
.B2(n_103),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_140),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_139),
.B(n_142),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_85),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_91),
.A2(n_35),
.B1(n_22),
.B2(n_44),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_33),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_33),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_87),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_151),
.Y(n_185)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_152),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_110),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_147),
.A2(n_97),
.B1(n_108),
.B2(n_84),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_153),
.A2(n_171),
.B1(n_180),
.B2(n_128),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_97),
.B1(n_92),
.B2(n_86),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_158),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_114),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_118),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_160),
.A2(n_162),
.B(n_178),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_88),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_88),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_165),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_81),
.B1(n_99),
.B2(n_98),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_117),
.A2(n_112),
.B1(n_100),
.B2(n_113),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_117),
.A2(n_107),
.B1(n_116),
.B2(n_80),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_173),
.B1(n_137),
.B2(n_128),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_146),
.Y(n_170)
);

AO21x2_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_109),
.B(n_89),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_175),
.B1(n_176),
.B2(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_102),
.B1(n_80),
.B2(n_115),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_110),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_122),
.A2(n_105),
.B1(n_109),
.B2(n_115),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_95),
.B1(n_41),
.B2(n_33),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_0),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_41),
.B1(n_33),
.B2(n_27),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_135),
.B1(n_141),
.B2(n_143),
.Y(n_180)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_187),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_186),
.B(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_134),
.C(n_140),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_190),
.C(n_205),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_138),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_178),
.A3(n_173),
.B1(n_158),
.B2(n_174),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_134),
.B1(n_136),
.B2(n_121),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_152),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_201),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_137),
.B(n_121),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_206),
.B(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_166),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_202),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_144),
.B(n_123),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_210),
.B(n_177),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_168),
.B1(n_169),
.B2(n_154),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_161),
.B1(n_148),
.B2(n_155),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_144),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_123),
.B(n_27),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_123),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_213),
.Y(n_221)
);

OAI21x1_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_8),
.B(n_14),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_1),
.B(n_2),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_8),
.Y(n_212)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_167),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_9),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_211),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_219),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_185),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_231),
.Y(n_259)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_229),
.B1(n_235),
.B2(n_238),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_188),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_195),
.B1(n_189),
.B2(n_171),
.Y(n_248)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

AOI22x1_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_206),
.B1(n_184),
.B2(n_195),
.Y(n_234)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_237),
.B(n_197),
.C(n_204),
.Y(n_246)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_214),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_210),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_184),
.A2(n_175),
.B(n_151),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_179),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_246),
.A2(n_237),
.B(n_224),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_190),
.C(n_205),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_253),
.C(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_252),
.B1(n_260),
.B2(n_235),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_232),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_254),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_182),
.B1(n_189),
.B2(n_194),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_236),
.C(n_223),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_261),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_197),
.B1(n_182),
.B2(n_200),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_256),
.A2(n_217),
.B1(n_215),
.B2(n_218),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_196),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_200),
.B1(n_196),
.B2(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_212),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_224),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_239),
.C(n_217),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_225),
.B(n_227),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_221),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_271),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_275),
.B(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_220),
.C(n_223),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_262),
.C(n_256),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_241),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_278),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_220),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_246),
.B1(n_248),
.B2(n_244),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_228),
.Y(n_280)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_280),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_252),
.B(n_15),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_15),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_286),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_254),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_14),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_282),
.B1(n_276),
.B2(n_271),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_250),
.B1(n_249),
.B2(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_245),
.C(n_266),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_300),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_275),
.A2(n_257),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_300),
.B1(n_290),
.B2(n_301),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_286),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_307),
.B(n_309),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_283),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_294),
.B(n_291),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_312),
.C(n_314),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_269),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_315),
.B(n_296),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_274),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_278),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_289),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_10),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_312),
.C(n_305),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_317),
.A2(n_322),
.B(n_316),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_12),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_304),
.A2(n_301),
.B(n_302),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_302),
.B1(n_10),
.B2(n_11),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_323),
.A2(n_13),
.B1(n_5),
.B2(n_6),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_313),
.A2(n_10),
.B(n_12),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_308),
.B(n_303),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_326),
.B(n_329),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_331),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_330),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_321),
.B(n_13),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_327),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_332),
.A2(n_331),
.B(n_317),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_337),
.Y(n_338)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_333),
.B1(n_334),
.B2(n_325),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_325),
.B(n_318),
.Y(n_340)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_331),
.C2(n_338),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_6),
.B(n_7),
.Y(n_342)
);


endmodule