module fake_jpeg_24970_n_168 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_42),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_41),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_9),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

OR2x2_ASAP7_75t_SL g42 ( 
.A(n_20),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_9),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_21),
.Y(n_52)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_47),
.B(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_54),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_21),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_28),
.B1(n_23),
.B2(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_35),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_14),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_17),
.Y(n_75)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_13),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_75),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_33),
.C(n_22),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_77),
.C(n_29),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_78),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_17),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_34),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_48),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_87),
.B(n_88),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_91),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_13),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_27),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_100),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_104),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_72),
.Y(n_120)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_29),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_64),
.B1(n_61),
.B2(n_51),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_81),
.B1(n_65),
.B2(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_64),
.B1(n_61),
.B2(n_27),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_80),
.B1(n_89),
.B2(n_90),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_119),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_83),
.B1(n_79),
.B2(n_84),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_114),
.B1(n_95),
.B2(n_53),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_106),
.B1(n_101),
.B2(n_107),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_74),
.B(n_73),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_122),
.B(n_108),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_121),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_97),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_70),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_137),
.B(n_132),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_130),
.A2(n_120),
.B(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_133),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_123),
.A2(n_110),
.A3(n_106),
.B1(n_102),
.B2(n_87),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_136),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_1),
.B(n_2),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_114),
.B1(n_112),
.B2(n_116),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_140),
.B1(n_127),
.B2(n_53),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_142),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_1),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_136),
.B(n_53),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_129),
.C(n_137),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_149),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_146),
.C(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_153),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_145),
.B(n_4),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_6),
.Y(n_162)
);

OAI31xp33_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_2),
.A3(n_4),
.B(n_5),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_2),
.B(n_4),
.Y(n_161)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_159),
.A2(n_161),
.B(n_162),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_150),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_147),
.C(n_157),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_155),
.B(n_160),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_166),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_6),
.B1(n_66),
.B2(n_148),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_66),
.Y(n_168)
);


endmodule