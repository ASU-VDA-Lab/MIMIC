module fake_jpeg_10271_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVxp67_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_4),
.A2(n_7),
.B(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_22),
.B1(n_14),
.B2(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_11),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_22)
);

CKINVDCx6p67_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_22),
.B1(n_19),
.B2(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_21),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_32),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_17),
.B1(n_20),
.B2(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_26),
.B1(n_17),
.B2(n_25),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_18),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_36),
.B1(n_38),
.B2(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_28),
.B(n_32),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_42),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_26),
.C(n_24),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_8),
.B1(n_15),
.B2(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_38),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_37),
.C(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_49),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_8),
.C(n_9),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_23),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_34),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_41),
.B1(n_23),
.B2(n_24),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_23),
.B(n_9),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_48),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_51),
.B1(n_9),
.B2(n_6),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_2),
.B(n_6),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_58),
.Y(n_60)
);

AOI221xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_57),
.B1(n_54),
.B2(n_7),
.C(n_6),
.Y(n_61)
);


endmodule