module fake_jpeg_22621_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx24_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_11),
.B(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_16),
.B1(n_10),
.B2(n_12),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_16),
.B1(n_21),
.B2(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_47),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_12),
.B(n_20),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_53),
.B(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_48),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_49),
.B1(n_18),
.B2(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.C(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_13),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_17),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_20),
.B(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_64),
.B(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_60),
.B1(n_52),
.B2(n_48),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_21),
.B1(n_14),
.B2(n_11),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_68),
.Y(n_77)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_74),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_58),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_45),
.B1(n_52),
.B2(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_29),
.C(n_19),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_78),
.C(n_56),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_29),
.C(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_2),
.Y(n_79)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

AOI21x1_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_64),
.B(n_57),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_57),
.B1(n_62),
.B2(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_87),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_69),
.B1(n_77),
.B2(n_76),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_83),
.B1(n_62),
.B2(n_86),
.Y(n_97)
);

AO221x1_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_77),
.B1(n_71),
.B2(n_4),
.C(n_5),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_60),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_82),
.C(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_92),
.B1(n_88),
.B2(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_98),
.B(n_66),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

AOI31xp67_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_67),
.A3(n_89),
.B(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_94),
.C(n_95),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_103),
.A2(n_73),
.B(n_89),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

AOI21x1_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_9),
.B(n_2),
.Y(n_108)
);

OAI321xp33_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_108),
.A3(n_106),
.B1(n_9),
.B2(n_3),
.C(n_104),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_3),
.Y(n_110)
);


endmodule