module fake_jpeg_3081_n_564 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_564);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_564;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_62),
.B(n_115),
.Y(n_124)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_66),
.B(n_68),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_67),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_72),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_80),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_74),
.Y(n_193)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_32),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_15),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_90),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_85),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_87),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_93),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_42),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g94 ( 
.A(n_23),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_95),
.B(n_98),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_21),
.B(n_16),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_104),
.B(n_105),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_49),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_49),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_111),
.Y(n_138)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_26),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_19),
.Y(n_112)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_113),
.Y(n_164)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_57),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_26),
.B(n_0),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_47),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_57),
.Y(n_141)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_23),
.Y(n_118)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_62),
.A2(n_37),
.B1(n_31),
.B2(n_22),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_121),
.B(n_131),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

NAND2x1_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_57),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_57),
.B1(n_46),
.B2(n_39),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_137),
.A2(n_149),
.B1(n_159),
.B2(n_180),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_37),
.B1(n_31),
.B2(n_22),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_139),
.A2(n_158),
.B1(n_138),
.B2(n_174),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_141),
.B(n_46),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_58),
.A2(n_29),
.B1(n_56),
.B2(n_47),
.Y(n_149)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_155),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_77),
.B(n_29),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_158),
.B(n_170),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_87),
.A2(n_21),
.B1(n_52),
.B2(n_51),
.Y(n_159)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_163),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_91),
.B(n_56),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_165),
.B(n_181),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_116),
.B(n_57),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_97),
.A2(n_36),
.B1(n_52),
.B2(n_51),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_171),
.A2(n_75),
.B1(n_107),
.B2(n_84),
.Y(n_204)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_60),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_173),
.Y(n_197)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_114),
.A2(n_35),
.B1(n_45),
.B2(n_36),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_108),
.B(n_45),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_69),
.A2(n_35),
.B1(n_16),
.B2(n_46),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_89),
.B1(n_81),
.B2(n_103),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_94),
.A2(n_46),
.B1(n_54),
.B2(n_28),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_112),
.B1(n_118),
.B2(n_100),
.Y(n_225)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_113),
.B(n_46),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_187),
.B(n_71),
.Y(n_200)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_63),
.Y(n_188)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_64),
.Y(n_189)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_71),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_65),
.Y(n_192)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_198),
.Y(n_323)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_199),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_219),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_201),
.B(n_202),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_122),
.B(n_79),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_204),
.A2(n_215),
.B1(n_227),
.B2(n_262),
.Y(n_267)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_205),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_170),
.A2(n_109),
.B(n_54),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_210),
.A2(n_235),
.B(n_251),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_101),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_211),
.B(n_222),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_132),
.Y(n_214)
);

INVx8_ASAP7_75t_L g270 ( 
.A(n_214),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_139),
.A2(n_67),
.B1(n_61),
.B2(n_110),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_216),
.A2(n_193),
.B1(n_144),
.B2(n_135),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_217),
.Y(n_318)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_125),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_125),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_221),
.B(n_231),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_88),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_225),
.A2(n_194),
.B1(n_145),
.B2(n_151),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_124),
.B(n_99),
.C(n_96),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_226),
.B(n_9),
.C(n_11),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_124),
.A2(n_86),
.B1(n_83),
.B2(n_74),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_228),
.B(n_205),
.Y(n_322)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_230),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_169),
.Y(n_231)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_136),
.Y(n_233)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_147),
.Y(n_234)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_235),
.B(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_127),
.B(n_1),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_169),
.B(n_2),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_243),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_150),
.Y(n_239)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_127),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_156),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_133),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_247),
.Y(n_268)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_153),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_254),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_126),
.A2(n_25),
.B(n_4),
.C(n_6),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_251),
.B(n_9),
.Y(n_299)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_162),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_253),
.Y(n_276)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_164),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_120),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_256),
.Y(n_304)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_258),
.B(n_260),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_156),
.B(n_129),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_261),
.Y(n_312)
);

INVx3_ASAP7_75t_SL g260 ( 
.A(n_119),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_178),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_149),
.A2(n_25),
.B1(n_4),
.B2(n_6),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_123),
.B(n_3),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_263),
.B(n_220),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_264),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_210),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_265),
.B(n_314),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_206),
.A2(n_131),
.B(n_137),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_271),
.B(n_302),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_273),
.A2(n_292),
.B1(n_306),
.B2(n_310),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g367 ( 
.A1(n_274),
.A2(n_297),
.B(n_299),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_209),
.A2(n_144),
.B1(n_140),
.B2(n_134),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_277),
.A2(n_316),
.B1(n_242),
.B2(n_247),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

O2A1O1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_206),
.A2(n_123),
.B(n_166),
.C(n_130),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_286),
.A2(n_213),
.B(n_249),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_248),
.A2(n_152),
.B1(n_146),
.B2(n_143),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_290),
.A2(n_256),
.B1(n_255),
.B2(n_212),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_228),
.A2(n_185),
.B1(n_175),
.B2(n_148),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_291),
.A2(n_268),
.B1(n_280),
.B2(n_286),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_226),
.A2(n_148),
.B1(n_175),
.B2(n_7),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_227),
.B(n_4),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_298),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_196),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_296),
.Y(n_341)
);

OA22x2_ASAP7_75t_L g297 ( 
.A1(n_204),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_244),
.B(n_7),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_299),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_207),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_196),
.B(n_12),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_216),
.A2(n_12),
.B1(n_13),
.B2(n_224),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_223),
.B(n_195),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_307),
.B(n_313),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_233),
.A2(n_240),
.B1(n_252),
.B2(n_234),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_203),
.B(n_207),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_257),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_253),
.A2(n_258),
.B1(n_197),
.B2(n_203),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_249),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_261),
.B1(n_213),
.B2(n_232),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_324),
.B(n_293),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_325),
.B(n_347),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g377 ( 
.A1(n_329),
.A2(n_351),
.B1(n_315),
.B2(n_303),
.Y(n_377)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

INVx13_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_332),
.B(n_339),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_265),
.B(n_197),
.C(n_212),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_356),
.C(n_361),
.Y(n_375)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_275),
.Y(n_334)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_307),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_343),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_269),
.B(n_260),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_342),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_239),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_304),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_284),
.B(n_264),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_355),
.Y(n_390)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_275),
.Y(n_346)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_346),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_305),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_279),
.B(n_208),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_348),
.B(n_350),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_322),
.A2(n_214),
.B1(n_217),
.B2(n_230),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_349),
.A2(n_268),
.B1(n_280),
.B2(n_320),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_276),
.Y(n_350)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_287),
.B(n_323),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_301),
.B(n_300),
.C(n_271),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_322),
.A2(n_267),
.B1(n_277),
.B2(n_274),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_359),
.B1(n_360),
.B2(n_304),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_266),
.B(n_287),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_364),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_292),
.A2(n_273),
.B1(n_288),
.B2(n_294),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_312),
.B(n_283),
.C(n_289),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_362),
.Y(n_403)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_276),
.Y(n_363)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_276),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_288),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_368),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_304),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_366),
.B(n_272),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_367),
.A2(n_296),
.B(n_278),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_289),
.B(n_309),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_369),
.A2(n_383),
.B(n_391),
.Y(n_422)
);

OA22x2_ASAP7_75t_L g370 ( 
.A1(n_357),
.A2(n_297),
.B1(n_316),
.B2(n_306),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_370),
.B(n_401),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_326),
.A2(n_302),
.B1(n_298),
.B2(n_297),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_371),
.A2(n_378),
.B1(n_384),
.B2(n_400),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_356),
.B(n_302),
.Y(n_372)
);

XNOR2x1_ASAP7_75t_L g433 ( 
.A(n_372),
.B(n_405),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_377),
.B1(n_396),
.B2(n_399),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_368),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_381),
.B(n_325),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_328),
.A2(n_336),
.B(n_355),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_326),
.A2(n_297),
.B1(n_317),
.B2(n_309),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_324),
.B(n_317),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_333),
.C(n_338),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_332),
.A2(n_314),
.B(n_285),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_339),
.B(n_352),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_328),
.A2(n_283),
.B(n_308),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_336),
.A2(n_285),
.B(n_308),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_394),
.A2(n_344),
.B(n_362),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_359),
.A2(n_320),
.B1(n_318),
.B2(n_310),
.Y(n_396)
);

AOI22x1_ASAP7_75t_SL g399 ( 
.A1(n_367),
.A2(n_315),
.B1(n_293),
.B2(n_303),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_337),
.A2(n_318),
.B1(n_282),
.B2(n_270),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_330),
.B(n_335),
.Y(n_401)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_393),
.Y(n_408)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_408),
.Y(n_442)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_393),
.Y(n_409)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_410),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_361),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_427),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_430),
.C(n_388),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_383),
.A2(n_366),
.B(n_350),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_414),
.A2(n_425),
.B(n_434),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_401),
.A2(n_335),
.B1(n_327),
.B2(n_365),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_417),
.A2(n_420),
.B1(n_421),
.B2(n_386),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_418),
.A2(n_384),
.B(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_379),
.A2(n_396),
.B1(n_380),
.B2(n_395),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_379),
.A2(n_340),
.B1(n_341),
.B2(n_364),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_373),
.B(n_347),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_424),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_382),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_358),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_432),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_340),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_392),
.Y(n_428)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_395),
.A2(n_374),
.B1(n_399),
.B2(n_397),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_415),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_375),
.B(n_354),
.C(n_363),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_380),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_431),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_394),
.A2(n_369),
.B(n_389),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_435),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_372),
.B(n_375),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_388),
.Y(n_444)
);

FAx1_ASAP7_75t_SL g437 ( 
.A(n_371),
.B(n_391),
.CI(n_376),
.CON(n_437),
.SN(n_437)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_402),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_390),
.B(n_348),
.Y(n_438)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_438),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_431),
.B(n_380),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_444),
.C(n_446),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_438),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_462),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_436),
.B(n_403),
.C(n_402),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_450),
.A2(n_456),
.B1(n_460),
.B2(n_416),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_412),
.B(n_390),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_453),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_403),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_SL g484 ( 
.A(n_455),
.B(n_464),
.C(n_437),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_430),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_345),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_420),
.A2(n_415),
.B1(n_416),
.B2(n_411),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_414),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_413),
.B(n_386),
.C(n_404),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_422),
.C(n_425),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_421),
.Y(n_466)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_466),
.Y(n_472)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_451),
.Y(n_467)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_467),
.Y(n_495)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_468),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_453),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_448),
.B(n_342),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_473),
.B(n_475),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_407),
.Y(n_474)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_474),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_449),
.B(n_417),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_407),
.Y(n_476)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_476),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_441),
.B(n_427),
.C(n_422),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_483),
.C(n_485),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_440),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_478),
.B(n_282),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_404),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_479),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_456),
.Y(n_480)
);

INVx13_ASAP7_75t_L g505 ( 
.A(n_480),
.Y(n_505)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_454),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_481),
.B(n_484),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_460),
.A2(n_418),
.B1(n_437),
.B2(n_434),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_482),
.A2(n_457),
.B1(n_464),
.B2(n_455),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_435),
.C(n_419),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_428),
.C(n_410),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_443),
.B(n_370),
.C(n_353),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_444),
.C(n_463),
.Y(n_504)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_447),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_446),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_491),
.B(n_502),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_492),
.A2(n_370),
.B1(n_334),
.B2(n_346),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_470),
.A2(n_450),
.B1(n_439),
.B2(n_452),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_493),
.A2(n_498),
.B1(n_508),
.B2(n_489),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_482),
.A2(n_457),
.B(n_439),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_494),
.A2(n_331),
.B(n_295),
.Y(n_521)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_496),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_472),
.A2(n_474),
.B1(n_486),
.B2(n_476),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_507),
.C(n_469),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_442),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_489),
.A2(n_400),
.B1(n_349),
.B2(n_351),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_398),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_521),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_512),
.A2(n_501),
.B1(n_498),
.B2(n_497),
.Y(n_534)
);

AOI21xp33_ASAP7_75t_L g513 ( 
.A1(n_493),
.A2(n_484),
.B(n_479),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_517),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_500),
.A2(n_471),
.B1(n_477),
.B2(n_490),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_514),
.B(n_520),
.Y(n_535)
);

OAI221xp5_ASAP7_75t_L g515 ( 
.A1(n_503),
.A2(n_469),
.B1(n_483),
.B2(n_485),
.C(n_488),
.Y(n_515)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_515),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_487),
.Y(n_516)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_516),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_500),
.A2(n_467),
.B1(n_341),
.B2(n_370),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_518),
.B(n_519),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_510),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_311),
.C(n_331),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_522),
.B(n_499),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_311),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_495),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_494),
.A2(n_295),
.B(n_270),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_524),
.A2(n_496),
.B(n_495),
.Y(n_530)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_527),
.Y(n_540)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_530),
.Y(n_546)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_532),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_534),
.B(n_536),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_514),
.A2(n_497),
.B(n_501),
.Y(n_536)
);

XNOR2x1_ASAP7_75t_SL g537 ( 
.A(n_519),
.B(n_491),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_537),
.B(n_507),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_511),
.B(n_504),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_522),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_531),
.B(n_525),
.C(n_502),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_541),
.B(n_543),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_544),
.B(n_537),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_528),
.B(n_526),
.C(n_524),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_545),
.B(n_547),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_520),
.C(n_521),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_533),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_549),
.A2(n_554),
.B(n_517),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_529),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_551),
.B(n_552),
.Y(n_557)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_546),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_555),
.B(n_556),
.C(n_558),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_553),
.B(n_541),
.C(n_542),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_550),
.B(n_534),
.C(n_539),
.Y(n_558)
);

NOR3xp33_ASAP7_75t_L g559 ( 
.A(n_557),
.B(n_549),
.C(n_523),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_559),
.B(n_516),
.Y(n_561)
);

OAI321xp33_ASAP7_75t_L g562 ( 
.A1(n_561),
.A2(n_560),
.A3(n_535),
.B1(n_505),
.B2(n_547),
.C(n_508),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_535),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_563),
.B(n_505),
.Y(n_564)
);


endmodule