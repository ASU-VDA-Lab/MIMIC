module fake_jpeg_1652_n_594 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_594);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_594;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_483;
wire n_236;
wire n_291;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_59),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_60),
.Y(n_127)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_61),
.Y(n_149)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_64),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_24),
.B(n_7),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_65),
.B(n_78),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_68),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_73),
.Y(n_207)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx10_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_77),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_15),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_33),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_82),
.B(n_84),
.Y(n_128)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_29),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_23),
.B(n_15),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_85),
.B(n_87),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_36),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_88),
.B(n_94),
.Y(n_184)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_90),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_92),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_93),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_17),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_39),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_96),
.B(n_100),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_99),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_39),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_101),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_30),
.B(n_10),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_30),
.B(n_10),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_107),
.Y(n_208)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_44),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_116),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_112),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_44),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_41),
.B(n_9),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_122),
.Y(n_214)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_41),
.B(n_8),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_124),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_21),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_27),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

INVx2_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_130),
.B(n_141),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_133),
.B(n_160),
.Y(n_216)
);

INVx2_ASAP7_75t_R g141 ( 
.A(n_71),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_64),
.B(n_31),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_147),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_76),
.B(n_51),
.C(n_49),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_148),
.B(n_55),
.C(n_49),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_80),
.B(n_26),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_165),
.B(n_173),
.Y(n_229)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_79),
.Y(n_169)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_93),
.B(n_48),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_171),
.B(n_200),
.Y(n_231)
);

BUFx16f_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

BUFx24_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_91),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_97),
.Y(n_176)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_176),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_104),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_177),
.B(n_190),
.Y(n_242)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_60),
.Y(n_187)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_187),
.Y(n_288)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_66),
.Y(n_188)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_107),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_68),
.A2(n_21),
.B1(n_26),
.B2(n_52),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_192),
.A2(n_125),
.B1(n_113),
.B2(n_32),
.Y(n_237)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_69),
.Y(n_195)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_198),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g199 ( 
.A(n_112),
.B(n_86),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_199),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_115),
.B(n_51),
.Y(n_200)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_90),
.A2(n_50),
.B1(n_31),
.B2(n_26),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_45),
.B(n_32),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_119),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_124),
.B1(n_114),
.B2(n_55),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_219),
.Y(n_310)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_220),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_175),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_221),
.B(n_241),
.Y(n_301)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_127),
.Y(n_226)
);

INVx3_ASAP7_75t_SL g308 ( 
.A(n_226),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_227),
.A2(n_134),
.B(n_152),
.Y(n_300)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_232),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_233),
.B(n_138),
.Y(n_305)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_234),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_199),
.A2(n_81),
.B1(n_75),
.B2(n_34),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_235),
.A2(n_237),
.B1(n_239),
.B2(n_243),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_238),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_161),
.A2(n_45),
.B1(n_34),
.B2(n_44),
.Y(n_239)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_150),
.Y(n_240)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_240),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_0),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_142),
.A2(n_81),
.B1(n_40),
.B2(n_27),
.Y(n_243)
);

INVx6_ASAP7_75t_SL g245 ( 
.A(n_172),
.Y(n_245)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_247),
.Y(n_293)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_128),
.A2(n_44),
.B1(n_40),
.B2(n_56),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_249),
.A2(n_279),
.B1(n_210),
.B2(n_163),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_128),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_250),
.B(n_258),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_142),
.A2(n_44),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

BUFx8_ASAP7_75t_L g320 ( 
.A(n_251),
.Y(n_320)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_252),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_151),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_253),
.B(n_271),
.Y(n_296)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_137),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_254),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_154),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_255),
.A2(n_265),
.B1(n_278),
.B2(n_289),
.Y(n_322)
);

BUFx16f_ASAP7_75t_L g257 ( 
.A(n_132),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_257),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_178),
.B(n_0),
.Y(n_258)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_137),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_260),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_200),
.B(n_22),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_165),
.C(n_135),
.Y(n_295)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_136),
.Y(n_262)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_262),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_151),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_263),
.B(n_267),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_167),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_265)
);

CKINVDCx12_ASAP7_75t_R g266 ( 
.A(n_132),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_266),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_178),
.B(n_205),
.Y(n_267)
);

INVx11_ASAP7_75t_L g270 ( 
.A(n_170),
.Y(n_270)
);

BUFx4f_ASAP7_75t_L g291 ( 
.A(n_270),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_211),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_4),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_275),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_213),
.B(n_4),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_181),
.Y(n_276)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_276),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_184),
.B(n_5),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_280),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_155),
.A2(n_6),
.B1(n_22),
.B2(n_56),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_206),
.A2(n_6),
.B1(n_56),
.B2(n_184),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_141),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_130),
.B(n_6),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_157),
.B(n_56),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_180),
.Y(n_283)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_171),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_285),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_193),
.B(n_201),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_196),
.B(n_168),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_287),
.B(n_182),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_215),
.A2(n_149),
.B1(n_166),
.B2(n_186),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_134),
.Y(n_290)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_231),
.B(n_131),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_294),
.B(n_223),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_295),
.B(n_255),
.Y(n_372)
);

OAI21xp33_ASAP7_75t_SL g353 ( 
.A1(n_300),
.A2(n_312),
.B(n_243),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_305),
.B(n_316),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_216),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_315),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_261),
.B(n_146),
.C(n_202),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_219),
.C(n_246),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_242),
.Y(n_315)
);

AOI32xp33_ASAP7_75t_L g316 ( 
.A1(n_261),
.A2(n_159),
.A3(n_179),
.B1(n_132),
.B2(n_158),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_222),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_317),
.B(n_326),
.Y(n_358)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_217),
.Y(n_324)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_324),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_222),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

AO21x2_ASAP7_75t_L g332 ( 
.A1(n_237),
.A2(n_163),
.B(n_158),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g377 ( 
.A1(n_332),
.A2(n_289),
.B1(n_251),
.B2(n_283),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_253),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_339),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_233),
.B(n_162),
.CI(n_158),
.CON(n_338),
.SN(n_338)
);

NOR2x1_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_344),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_269),
.A2(n_194),
.B1(n_207),
.B2(n_197),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_340),
.A2(n_341),
.B1(n_342),
.B2(n_228),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_230),
.A2(n_194),
.B1(n_207),
.B2(n_197),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_230),
.A2(n_153),
.B1(n_212),
.B2(n_144),
.Y(n_342)
);

AO22x1_ASAP7_75t_L g344 ( 
.A1(n_229),
.A2(n_246),
.B1(n_235),
.B2(n_220),
.Y(n_344)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_347),
.Y(n_412)
);

CKINVDCx11_ASAP7_75t_R g348 ( 
.A(n_297),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_382),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_296),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_349),
.B(n_355),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_310),
.A2(n_232),
.B1(n_247),
.B2(n_234),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_351),
.A2(n_236),
.B1(n_293),
.B2(n_299),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_367),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_354),
.B(n_322),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_301),
.B(n_274),
.Y(n_355)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_357),
.Y(n_396)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_319),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_359),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_294),
.B(n_314),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_365),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_264),
.C(n_273),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_362),
.B(n_372),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_218),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_364),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_294),
.B(n_288),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_345),
.A2(n_310),
.B1(n_300),
.B2(n_344),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_366),
.A2(n_369),
.B1(n_332),
.B2(n_312),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_224),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_368),
.B(n_383),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_300),
.A2(n_244),
.B1(n_256),
.B2(n_268),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_320),
.A2(n_332),
.B(n_338),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_370),
.A2(n_320),
.B(n_332),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_320),
.A2(n_270),
.B1(n_236),
.B2(n_262),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_371),
.Y(n_414)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_297),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_276),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_375),
.A2(n_342),
.B(n_341),
.Y(n_397)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_336),
.Y(n_376)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_376),
.Y(n_393)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_378),
.Y(n_420)
);

BUFx12f_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

INVx6_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_380),
.A2(n_386),
.B1(n_365),
.B2(n_358),
.Y(n_401)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_295),
.B(n_257),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_292),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_384),
.B(n_385),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_333),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_327),
.B(n_252),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_386),
.B(n_309),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_304),
.B(n_286),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_387),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_303),
.B(n_260),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_388),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_323),
.B(n_254),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_389),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_368),
.B1(n_366),
.B2(n_372),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_390),
.A2(n_377),
.B1(n_352),
.B2(n_308),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_419),
.B1(n_402),
.B2(n_354),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_418),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_398),
.B(n_403),
.Y(n_442)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_363),
.A2(n_298),
.A3(n_293),
.B1(n_322),
.B2(n_302),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_337),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_404),
.B(n_416),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_350),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_406),
.B(n_408),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_374),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_360),
.A2(n_367),
.B1(n_383),
.B2(n_369),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_373),
.Y(n_424)
);

INVx13_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_426),
.A2(n_453),
.B1(n_411),
.B2(n_425),
.Y(n_464)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_410),
.Y(n_427)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_422),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_429),
.B(n_434),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_362),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_430),
.B(n_432),
.Y(n_462)
);

AO22x1_ASAP7_75t_L g431 ( 
.A1(n_402),
.A2(n_375),
.B1(n_360),
.B2(n_367),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_443),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_399),
.B(n_409),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_413),
.Y(n_433)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_433),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_415),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g435 ( 
.A1(n_414),
.A2(n_375),
.B1(n_378),
.B2(n_347),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_423),
.Y(n_439)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_439),
.Y(n_457)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_423),
.Y(n_440)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_440),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_394),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_446),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_407),
.B(n_257),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_420),
.Y(n_444)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_356),
.Y(n_445)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_445),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_396),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_420),
.Y(n_447)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_447),
.Y(n_471)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

OA22x2_ASAP7_75t_L g450 ( 
.A1(n_390),
.A2(n_391),
.B1(n_411),
.B2(n_395),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_451),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_377),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_393),
.Y(n_452)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_452),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_416),
.A2(n_377),
.B1(n_376),
.B2(n_357),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_456),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_455),
.A2(n_411),
.B1(n_397),
.B2(n_392),
.Y(n_463)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_412),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_463),
.A2(n_469),
.B1(n_465),
.B2(n_481),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_464),
.A2(n_455),
.B1(n_431),
.B2(n_425),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_428),
.A2(n_392),
.B(n_403),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_465),
.B(n_480),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_400),
.C(n_404),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_482),
.C(n_485),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_428),
.A2(n_414),
.B(n_424),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_468),
.A2(n_469),
.B(n_481),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_453),
.A2(n_400),
.B(n_421),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_398),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_439),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_410),
.Y(n_479)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_479),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_437),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_431),
.A2(n_382),
.B(n_330),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_426),
.B(n_442),
.C(n_450),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_442),
.A2(n_343),
.B(n_318),
.Y(n_483)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_483),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_321),
.C(n_346),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_436),
.A2(n_421),
.B(n_291),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_456),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_462),
.B(n_427),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_488),
.B(n_458),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_489),
.A2(n_490),
.B1(n_491),
.B2(n_492),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_464),
.A2(n_436),
.B1(n_451),
.B2(n_450),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_470),
.A2(n_436),
.B1(n_443),
.B2(n_440),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_479),
.B(n_447),
.Y(n_493)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_493),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g514 ( 
.A(n_495),
.Y(n_514)
);

INVx3_ASAP7_75t_SL g496 ( 
.A(n_458),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_504),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_506),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_466),
.B(n_325),
.C(n_306),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_500),
.C(n_502),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_473),
.B(n_308),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_478),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_325),
.C(n_292),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_470),
.B(n_438),
.Y(n_501)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_501),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_313),
.C(n_319),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_478),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_463),
.B(n_438),
.Y(n_506)
);

CKINVDCx14_ASAP7_75t_R g507 ( 
.A(n_472),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_507),
.A2(n_476),
.B1(n_477),
.B2(n_484),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_313),
.C(n_212),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_508),
.B(n_486),
.C(n_468),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_460),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_509),
.B(n_510),
.Y(n_525)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_471),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_527),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_511),
.A2(n_459),
.B1(n_475),
.B2(n_474),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_516),
.A2(n_495),
.B1(n_504),
.B2(n_502),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_517),
.B(n_528),
.Y(n_536)
);

AOI21xp33_ASAP7_75t_L g520 ( 
.A1(n_494),
.A2(n_459),
.B(n_475),
.Y(n_520)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_520),
.Y(n_533)
);

FAx1_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_474),
.CI(n_471),
.CON(n_521),
.SN(n_521)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_521),
.A2(n_496),
.B(n_457),
.Y(n_543)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_524),
.Y(n_538)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_526),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_484),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_487),
.B(n_477),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_494),
.A2(n_461),
.B1(n_457),
.B2(n_467),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_529),
.A2(n_495),
.B1(n_493),
.B2(n_501),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_497),
.B(n_467),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_530),
.B(n_500),
.C(n_499),
.Y(n_535)
);

XNOR2x1_ASAP7_75t_L g531 ( 
.A(n_506),
.B(n_461),
.Y(n_531)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_531),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_525),
.B(n_498),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_537),
.Y(n_549)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_534),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_522),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_505),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_516),
.A2(n_503),
.B(n_489),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_539),
.A2(n_515),
.B(n_523),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_542),
.B(n_517),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_543),
.B(n_544),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_528),
.B(n_359),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_519),
.A2(n_508),
.B1(n_334),
.B2(n_291),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_546),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_512),
.B(n_530),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_541),
.B(n_512),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_550),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_536),
.B(n_522),
.C(n_531),
.Y(n_550)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_551),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_533),
.B(n_536),
.C(n_540),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_553),
.B(n_555),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_513),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_556),
.B(n_558),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_557),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_535),
.B(n_514),
.C(n_521),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g560 ( 
.A(n_547),
.B(n_521),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_542),
.Y(n_561)
);

CKINVDCx14_ASAP7_75t_R g573 ( 
.A(n_561),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_554),
.A2(n_538),
.B1(n_518),
.B2(n_529),
.Y(n_562)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_562),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_549),
.B(n_543),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_564),
.B(n_568),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_557),
.B(n_539),
.C(n_547),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_566),
.B(n_569),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_534),
.Y(n_568)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_552),
.Y(n_571)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_571),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_565),
.B(n_558),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_572),
.A2(n_563),
.B(n_566),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_570),
.B(n_550),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_575),
.B(n_576),
.Y(n_582)
);

MAJx2_ASAP7_75t_L g576 ( 
.A(n_567),
.B(n_560),
.C(n_545),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_579),
.B(n_563),
.C(n_562),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_580),
.A2(n_584),
.B(n_572),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_581),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_577),
.A2(n_379),
.B1(n_291),
.B2(n_248),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_583),
.Y(n_586)
);

O2A1O1Ixp33_ASAP7_75t_L g584 ( 
.A1(n_574),
.A2(n_379),
.B(n_225),
.C(n_226),
.Y(n_584)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_587),
.A2(n_225),
.B(n_145),
.C(n_156),
.Y(n_589)
);

AOI322xp5_ASAP7_75t_L g588 ( 
.A1(n_585),
.A2(n_578),
.A3(n_582),
.B1(n_586),
.B2(n_573),
.C1(n_238),
.C2(n_240),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_588),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_590),
.B(n_589),
.C(n_164),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_140),
.C(n_203),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_592),
.B(n_225),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_593),
.B(n_209),
.Y(n_594)
);


endmodule