module fake_jpeg_27880_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_55),
.Y(n_69)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_24),
.C(n_20),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_61),
.C(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_21),
.Y(n_73)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_22),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_73),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_41),
.B1(n_37),
.B2(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_74),
.B1(n_75),
.B2(n_84),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_41),
.B1(n_42),
.B2(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_42),
.B1(n_31),
.B2(n_32),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_76),
.Y(n_92)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_80),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2x1_ASAP7_75t_R g81 ( 
.A(n_56),
.B(n_31),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_86),
.B(n_22),
.C(n_30),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_38),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_35),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_42),
.B1(n_56),
.B2(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_32),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_38),
.B1(n_35),
.B2(n_30),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_54),
.B1(n_44),
.B2(n_64),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_108),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_19),
.B1(n_54),
.B2(n_22),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_95),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_96),
.A2(n_114),
.B(n_16),
.Y(n_137)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_90),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_68),
.A2(n_16),
.B1(n_27),
.B2(n_19),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_102),
.B(n_107),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_110),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_35),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_116),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_35),
.C(n_33),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_75),
.C(n_68),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_30),
.B(n_27),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_69),
.A2(n_44),
.B1(n_53),
.B2(n_48),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_83),
.B1(n_58),
.B2(n_59),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_113),
.C(n_94),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_140),
.B1(n_146),
.B2(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_134),
.B(n_136),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_72),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_96),
.B(n_104),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_141),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_110),
.A2(n_91),
.B1(n_47),
.B2(n_77),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_63),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_118),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_99),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_47),
.B1(n_86),
.B2(n_79),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_148),
.Y(n_151)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_154),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_138),
.C(n_133),
.Y(n_186)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_168),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_124),
.A3(n_145),
.B1(n_120),
.B2(n_128),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_170),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_102),
.B1(n_108),
.B2(n_98),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_164),
.B1(n_79),
.B2(n_33),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_102),
.B1(n_98),
.B2(n_100),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_167),
.B1(n_26),
.B2(n_25),
.Y(n_205)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_169),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_100),
.B1(n_116),
.B2(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_118),
.B(n_105),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_177),
.B(n_26),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_174),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_114),
.B1(n_101),
.B2(n_88),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_123),
.B1(n_137),
.B2(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_179),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_33),
.B(n_29),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_203),
.B1(n_208),
.B2(n_159),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_146),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_183),
.A2(n_189),
.B(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_155),
.C(n_160),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_122),
.B1(n_148),
.B2(n_134),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_177),
.B1(n_24),
.B2(n_23),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_139),
.B1(n_129),
.B2(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_190),
.B(n_192),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_191),
.B(n_29),
.C(n_23),
.Y(n_233)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_193),
.B(n_194),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_151),
.B(n_29),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_88),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_165),
.A2(n_90),
.B1(n_26),
.B2(n_25),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_90),
.B1(n_26),
.B2(n_25),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_152),
.B1(n_150),
.B2(n_153),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_24),
.B1(n_23),
.B2(n_20),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_215),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_187),
.C(n_1),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g212 ( 
.A(n_198),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_214),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_156),
.C(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_216),
.C(n_228),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_156),
.B1(n_180),
.B2(n_152),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_180),
.C(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_218),
.B(n_222),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_220),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_24),
.C(n_23),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_201),
.B1(n_183),
.B2(n_181),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_204),
.C(n_208),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_206),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_239),
.Y(n_262)
);

NAND4xp25_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_188),
.C(n_196),
.D(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_197),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_189),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_249),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_244),
.A2(n_219),
.B(n_226),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_183),
.C(n_203),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_247),
.C(n_250),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_8),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_8),
.C(n_1),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_7),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_220),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_209),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_249),
.C(n_235),
.Y(n_282)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_230),
.Y(n_265)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_248),
.B(n_227),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_214),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_269),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_237),
.A2(n_211),
.B(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_228),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_217),
.B(n_0),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_234),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_281),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_241),
.Y(n_278)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_239),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_260),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_256),
.A2(n_245),
.B1(n_253),
.B2(n_236),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_284),
.B1(n_260),
.B2(n_262),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_238),
.B1(n_2),
.B2(n_3),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_270),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_290),
.Y(n_298)
);

AOI21xp33_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_269),
.B(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_10),
.C(n_11),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_288),
.A2(n_294),
.B(n_278),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_275),
.B1(n_271),
.B2(n_11),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_5),
.B(n_9),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_5),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_274),
.Y(n_300)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_302),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_301),
.B(n_303),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_9),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_10),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_12),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_296),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_287),
.B(n_291),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_306),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_308),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_312),
.C(n_298),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_296),
.B(n_13),
.Y(n_312)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_314),
.A2(n_307),
.B(n_297),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_311),
.B(n_309),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_317),
.C(n_313),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_12),
.B(n_13),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_12),
.B(n_13),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_15),
.Y(n_321)
);


endmodule