module fake_jpeg_3030_n_226 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_54),
.C(n_53),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_90),
.Y(n_92)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_93),
.B1(n_100),
.B2(n_104),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_101),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_70),
.B1(n_56),
.B2(n_55),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_77),
.B1(n_63),
.B2(n_65),
.Y(n_109)
);

OA22x2_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_62),
.B1(n_60),
.B2(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_81),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_55),
.B1(n_56),
.B2(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_101),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_120),
.Y(n_141)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_83),
.B1(n_82),
.B2(n_60),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_110),
.B1(n_95),
.B2(n_99),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_41),
.B1(n_34),
.B2(n_33),
.Y(n_132)
);

OAI22x1_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_82),
.B1(n_75),
.B2(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_115),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_67),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_5),
.Y(n_138)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_63),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_117),
.A2(n_49),
.B(n_42),
.Y(n_131)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_121),
.Y(n_136)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_32),
.Y(n_145)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_79),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_77),
.B1(n_66),
.B2(n_65),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_66),
.B1(n_95),
.B2(n_78),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_126),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_74),
.B(n_62),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_10),
.B(n_12),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_0),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_134),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_133),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_2),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_122),
.B1(n_113),
.B2(n_11),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_26),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_6),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_7),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_113),
.B1(n_121),
.B2(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

AO22x2_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_149),
.B(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_169),
.B1(n_171),
.B2(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_156),
.Y(n_190)
);

AOI31xp33_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_13),
.A3(n_14),
.B(n_15),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_24),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_163),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_16),
.B(n_17),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_172),
.B(n_173),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_17),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_144),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_18),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_170),
.B(n_23),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_25),
.B1(n_20),
.B2(n_21),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_19),
.B(n_22),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_22),
.B(n_23),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_133),
.B1(n_145),
.B2(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_184),
.B1(n_192),
.B2(n_168),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_178),
.B(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

OAI321xp33_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_189),
.A3(n_172),
.B1(n_156),
.B2(n_163),
.C(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_147),
.B1(n_140),
.B2(n_144),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_165),
.C(n_167),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_187),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_150),
.B(n_162),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_167),
.B1(n_168),
.B2(n_151),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_196),
.B1(n_182),
.B2(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_177),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_185),
.Y(n_203)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_207),
.Y(n_213)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_208),
.B1(n_192),
.B2(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_174),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_184),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_196),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_210),
.B(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_210),
.A2(n_202),
.B(n_193),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_215),
.B1(n_204),
.B2(n_188),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_218),
.B1(n_209),
.B2(n_176),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_193),
.B1(n_188),
.B2(n_155),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_214),
.C(n_213),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_203),
.C(n_191),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_186),
.C(n_153),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_180),
.B(n_169),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_180),
.Y(n_226)
);


endmodule