module fake_jpeg_1470_n_611 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_611);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_611;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_26),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_61),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_60),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_26),
.B(n_0),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_96),
.Y(n_137)
);

BUFx12f_ASAP7_75t_SL g75 ( 
.A(n_54),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_57),
.Y(n_136)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_87),
.Y(n_132)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_81),
.Y(n_217)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_82),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_84),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_48),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_92),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_21),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_50),
.B(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_17),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_101),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_17),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_105),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_33),
.B(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_112),
.Y(n_157)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_21),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_110),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_34),
.B(n_3),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_57),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_113),
.B(n_119),
.Y(n_186)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_38),
.B(n_4),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_37),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_41),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_121),
.B(n_126),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

AND2x4_ASAP7_75t_SL g123 ( 
.A(n_41),
.B(n_4),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_123),
.B(n_22),
.Y(n_160)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_125),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_43),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_43),
.Y(n_127)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_22),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_119),
.B(n_56),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_131),
.B(n_140),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_57),
.B1(n_51),
.B2(n_45),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_134),
.A2(n_173),
.B1(n_179),
.B2(n_194),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_136),
.B(n_160),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_63),
.B(n_55),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_43),
.B1(n_45),
.B2(n_51),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_142),
.A2(n_159),
.B1(n_169),
.B2(n_177),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_71),
.A2(n_51),
.B1(n_45),
.B2(n_55),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_154),
.A2(n_198),
.B1(n_221),
.B2(n_118),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_75),
.A2(n_51),
.B1(n_45),
.B2(n_49),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_107),
.A2(n_22),
.B1(n_49),
.B2(n_35),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_123),
.A2(n_24),
.B1(n_46),
.B2(n_44),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_175),
.B(n_193),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_99),
.A2(n_37),
.B1(n_46),
.B2(n_44),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_176),
.A2(n_209),
.B(n_210),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_76),
.A2(n_53),
.B1(n_35),
.B2(n_49),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_73),
.A2(n_42),
.B1(n_25),
.B2(n_24),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_83),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_181),
.B(n_183),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_78),
.B(n_42),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_68),
.B(n_25),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_188),
.B(n_189),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_93),
.B(n_53),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_129),
.B(n_53),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_81),
.A2(n_35),
.B1(n_40),
.B2(n_52),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_84),
.A2(n_40),
.B1(n_52),
.B2(n_7),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_204),
.Y(n_293)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

INVx4_ASAP7_75t_SL g277 ( 
.A(n_208),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_125),
.A2(n_52),
.B1(n_6),
.B2(n_7),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_60),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_85),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_91),
.B(n_5),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_212),
.B(n_216),
.Y(n_296)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_58),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_220),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_95),
.B(n_8),
.Y(n_216)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_69),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_111),
.B(n_17),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_77),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_102),
.Y(n_222)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_224),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_197),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_225),
.B(n_232),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_226),
.A2(n_234),
.B1(n_251),
.B2(n_255),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_142),
.A2(n_100),
.B1(n_105),
.B2(n_62),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_229),
.A2(n_238),
.B1(n_252),
.B2(n_304),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_197),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_160),
.B(n_115),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_233),
.B(n_262),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_134),
.A2(n_82),
.B1(n_111),
.B2(n_104),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_235),
.Y(n_311)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_236),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_136),
.A2(n_70),
.B1(n_103),
.B2(n_98),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_237),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_142),
.A2(n_104),
.B1(n_67),
.B2(n_66),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_239),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_240),
.Y(n_334)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_241),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_165),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_242),
.B(n_266),
.Y(n_313)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_246),
.Y(n_314)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_167),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_248),
.Y(n_357)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_158),
.Y(n_250)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_250),
.Y(n_318)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_205),
.B(n_117),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_252),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_11),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_253),
.B(n_301),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_147),
.A2(n_117),
.B1(n_15),
.B2(n_16),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_159),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_256),
.A2(n_275),
.B1(n_281),
.B2(n_289),
.Y(n_310)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

INVx3_ASAP7_75t_SL g319 ( 
.A(n_257),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_171),
.Y(n_258)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_258),
.Y(n_339)
);

AND2x2_ASAP7_75t_SL g259 ( 
.A(n_188),
.B(n_14),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_280),
.C(n_244),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_261),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_143),
.B(n_14),
.Y(n_262)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_263),
.A2(n_270),
.B1(n_278),
.B2(n_295),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_174),
.Y(n_264)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_264),
.Y(n_360)
);

OR2x4_ASAP7_75t_L g265 ( 
.A(n_186),
.B(n_16),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_265),
.A2(n_253),
.B(n_269),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_157),
.B(n_16),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_272),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_156),
.Y(n_268)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_200),
.Y(n_269)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_149),
.A2(n_162),
.B1(n_182),
.B2(n_187),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_138),
.B(n_168),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_145),
.B(n_164),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_284),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_190),
.B(n_141),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_274),
.B(n_279),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_130),
.A2(n_137),
.B1(n_177),
.B2(n_169),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_215),
.A2(n_132),
.B1(n_150),
.B2(n_192),
.Y(n_276)
);

OA22x2_ASAP7_75t_L g362 ( 
.A1(n_276),
.A2(n_293),
.B1(n_260),
.B2(n_241),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_149),
.A2(n_187),
.B1(n_182),
.B2(n_162),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_153),
.B(n_166),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_180),
.B(n_155),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_196),
.A2(n_215),
.B1(n_135),
.B2(n_151),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_144),
.Y(n_282)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_282),
.Y(n_351)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_174),
.Y(n_283)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_199),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_156),
.Y(n_285)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

NAND2x1p5_ASAP7_75t_L g286 ( 
.A(n_133),
.B(n_184),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_286),
.A2(n_290),
.B(n_300),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_191),
.B(n_202),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_291),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_207),
.A2(n_135),
.B1(n_151),
.B2(n_161),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_202),
.B(n_195),
.Y(n_291)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_294),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_161),
.A2(n_223),
.B1(n_217),
.B2(n_172),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_217),
.B(n_223),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_300),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_172),
.A2(n_152),
.B1(n_218),
.B2(n_139),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_298),
.A2(n_302),
.B1(n_234),
.B2(n_295),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_158),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_148),
.B(n_170),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_170),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_152),
.A2(n_218),
.B1(n_148),
.B2(n_201),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_143),
.B(n_138),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_197),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_286),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_244),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_315),
.B(n_322),
.C(n_328),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_246),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_244),
.B(n_280),
.Y(n_322)
);

A2O1A1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_233),
.A2(n_265),
.B(n_266),
.C(n_245),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_324),
.B(n_340),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_272),
.Y(n_328)
);

OAI22x1_ASAP7_75t_SL g330 ( 
.A1(n_238),
.A2(n_254),
.B1(n_229),
.B2(n_226),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_330),
.A2(n_335),
.B1(n_350),
.B2(n_361),
.Y(n_370)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_331),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_239),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_296),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_344),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_248),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_286),
.A2(n_243),
.B(n_227),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_341),
.A2(n_354),
.B(n_336),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_259),
.B(n_279),
.Y(n_344)
);

NOR3xp33_ASAP7_75t_L g347 ( 
.A(n_287),
.B(n_262),
.C(n_243),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_254),
.Y(n_363)
);

OAI22x1_ASAP7_75t_SL g350 ( 
.A1(n_254),
.A2(n_230),
.B1(n_259),
.B2(n_252),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_253),
.B(n_267),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_293),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_355),
.B(n_277),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_254),
.A2(n_297),
.B1(n_294),
.B2(n_281),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_362),
.Y(n_367)
);

NAND3xp33_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_384),
.C(n_318),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_364),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_365),
.B(n_378),
.C(n_401),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_328),
.B(n_249),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_366),
.B(n_405),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_371),
.A2(n_372),
.B(n_385),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_331),
.A2(n_231),
.B(n_260),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_374),
.B(n_397),
.Y(n_419)
);

INVx6_ASAP7_75t_SL g375 ( 
.A(n_321),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_375),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_316),
.B(n_228),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_377),
.B(n_379),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_322),
.B(n_235),
.C(n_283),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_316),
.B(n_228),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_329),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_383),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_306),
.B(n_344),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_381),
.B(n_382),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_306),
.B(n_236),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_326),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_350),
.A2(n_307),
.B1(n_330),
.B2(n_310),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_386),
.A2(n_393),
.B1(n_400),
.B2(n_335),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_341),
.A2(n_324),
.B(n_354),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_387),
.A2(n_352),
.B(n_357),
.Y(n_425)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_327),
.Y(n_391)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_391),
.Y(n_415)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_309),
.Y(n_392)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_392),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_307),
.A2(n_257),
.B1(n_285),
.B2(n_268),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_357),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_404),
.Y(n_443)
);

INVx4_ASAP7_75t_SL g396 ( 
.A(n_318),
.Y(n_396)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_396),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_337),
.B(n_282),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_398),
.Y(n_426)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_342),
.Y(n_399)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_399),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_310),
.A2(n_289),
.B1(n_298),
.B2(n_301),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_315),
.B(n_299),
.C(n_264),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_402),
.Y(n_433)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_403),
.Y(n_444)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_311),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_349),
.B(n_224),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_313),
.B(n_247),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_406),
.B(n_339),
.Y(n_431)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_311),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_407),
.B(n_348),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_408),
.A2(n_412),
.B1(n_413),
.B2(n_418),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_386),
.A2(n_361),
.B1(n_345),
.B2(n_308),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_410),
.A2(n_414),
.B1(n_416),
.B2(n_441),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_367),
.A2(n_312),
.B1(n_305),
.B2(n_343),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_370),
.A2(n_305),
.B1(n_352),
.B2(n_353),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_370),
.A2(n_352),
.B1(n_343),
.B2(n_320),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_393),
.A2(n_367),
.B1(n_400),
.B2(n_388),
.Y(n_416)
);

OAI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_389),
.A2(n_323),
.B1(n_362),
.B2(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_365),
.B(n_323),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_439),
.C(n_442),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_425),
.A2(n_432),
.B(n_372),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_429),
.B(n_371),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_431),
.B(n_383),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_385),
.A2(n_334),
.B(n_362),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_388),
.A2(n_362),
.B1(n_319),
.B2(n_325),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_435),
.A2(n_380),
.B1(n_395),
.B2(n_398),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_375),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_436),
.B(n_333),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_368),
.B(n_346),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_387),
.A2(n_397),
.B1(n_382),
.B2(n_373),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_369),
.B(n_346),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_408),
.A2(n_389),
.B1(n_385),
.B2(n_377),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_447),
.A2(n_454),
.B1(n_457),
.B2(n_470),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_422),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_468),
.Y(n_482)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_450),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_451),
.A2(n_465),
.B(n_431),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_379),
.Y(n_453)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_453),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_455),
.B(n_475),
.Y(n_495)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_411),
.Y(n_456)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_456),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_416),
.A2(n_389),
.B1(n_368),
.B2(n_381),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_392),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_458),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_378),
.C(n_369),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_463),
.C(n_469),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_460),
.B(n_471),
.Y(n_488)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_415),
.Y(n_461)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_461),
.Y(n_504)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_401),
.C(n_364),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_409),
.B(n_374),
.Y(n_464)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_438),
.A2(n_390),
.B(n_391),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_423),
.B(n_366),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_428),
.Y(n_483)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_420),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_394),
.C(n_402),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_410),
.A2(n_399),
.B1(n_396),
.B2(n_403),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_443),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_441),
.A2(n_396),
.B1(n_325),
.B2(n_319),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_472),
.A2(n_473),
.B1(n_480),
.B2(n_435),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_414),
.A2(n_358),
.B1(n_407),
.B2(n_351),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_351),
.C(n_404),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_444),
.C(n_421),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_428),
.B(n_376),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_477),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_360),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_437),
.A2(n_333),
.B1(n_250),
.B2(n_263),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_427),
.B1(n_436),
.B2(n_421),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_443),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_417),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_437),
.A2(n_360),
.B1(n_334),
.B2(n_247),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_SL g513 ( 
.A1(n_481),
.A2(n_470),
.B1(n_464),
.B2(n_450),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_483),
.B(n_486),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_413),
.B1(n_419),
.B2(n_425),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_484),
.A2(n_487),
.B1(n_489),
.B2(n_507),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_438),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_466),
.A2(n_447),
.B1(n_452),
.B2(n_457),
.Y(n_489)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_492),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_446),
.B(n_440),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_501),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_448),
.B(n_419),
.Y(n_494)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_494),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_449),
.Y(n_496)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_496),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_499),
.B(n_461),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_446),
.B(n_417),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_427),
.Y(n_503)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_503),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_505),
.B(n_506),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_458),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_452),
.A2(n_454),
.B1(n_479),
.B2(n_465),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_453),
.B(n_426),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_473),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_467),
.B(n_424),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_511),
.B(n_430),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_513),
.A2(n_531),
.B1(n_490),
.B2(n_496),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_495),
.B(n_469),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_514),
.B(n_526),
.C(n_527),
.Y(n_542)
);

OAI221xp5_ASAP7_75t_L g515 ( 
.A1(n_494),
.A2(n_458),
.B1(n_451),
.B2(n_463),
.C(n_426),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_520),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_500),
.A2(n_476),
.B(n_472),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_517),
.A2(n_529),
.B(n_535),
.Y(n_540)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_519),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_474),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_480),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_522),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_505),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_523),
.B(n_528),
.Y(n_549)
);

AO22x1_ASAP7_75t_SL g524 ( 
.A1(n_507),
.A2(n_478),
.B1(n_456),
.B2(n_468),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_524),
.B(n_525),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_434),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_484),
.B(n_434),
.Y(n_527)
);

CKINVDCx14_ASAP7_75t_R g528 ( 
.A(n_492),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_493),
.B(n_430),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_503),
.B(n_462),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_490),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_483),
.B(n_420),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g538 ( 
.A(n_516),
.B(n_486),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_538),
.B(n_541),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_501),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_530),
.A2(n_489),
.B1(n_481),
.B2(n_510),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_544),
.Y(n_560)
);

OAI322xp33_ASAP7_75t_L g544 ( 
.A1(n_515),
.A2(n_500),
.A3(n_510),
.B1(n_497),
.B2(n_511),
.C1(n_482),
.C2(n_485),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_485),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_545),
.B(n_548),
.Y(n_567)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_546),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_516),
.B(n_499),
.C(n_482),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_551),
.C(n_556),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_521),
.B(n_502),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_531),
.C(n_512),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_552),
.B(n_517),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_497),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_553),
.B(n_554),
.Y(n_572)
);

AOI322xp5_ASAP7_75t_L g554 ( 
.A1(n_518),
.A2(n_491),
.A3(n_504),
.B1(n_498),
.B2(n_509),
.C1(n_433),
.C2(n_444),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_531),
.B(n_491),
.C(n_498),
.Y(n_556)
);

O2A1O1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_537),
.A2(n_536),
.B(n_530),
.C(n_518),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_557),
.B(n_558),
.Y(n_585)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_549),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_559),
.B(n_562),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_552),
.A2(n_536),
.B1(n_533),
.B2(n_519),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_561),
.A2(n_539),
.B1(n_550),
.B2(n_553),
.Y(n_576)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_546),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_556),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_563),
.B(n_570),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_534),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_539),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_545),
.B(n_522),
.C(n_524),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_568),
.B(n_569),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_522),
.C(n_524),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_542),
.Y(n_570)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_573),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_565),
.B(n_547),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_574),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_565),
.B(n_548),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_581),
.Y(n_586)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_576),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_561),
.A2(n_550),
.B1(n_551),
.B2(n_533),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_580),
.B(n_567),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_560),
.B(n_433),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_572),
.B(n_504),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_583),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_557),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_567),
.B(n_538),
.C(n_540),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_584),
.A2(n_571),
.B(n_509),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g588 ( 
.A1(n_578),
.A2(n_558),
.B(n_564),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_588),
.B(n_590),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_585),
.A2(n_568),
.B(n_569),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_576),
.C(n_573),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_579),
.A2(n_564),
.B(n_566),
.Y(n_590)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_592),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_595),
.B(n_584),
.C(n_574),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_596),
.B(n_597),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_587),
.B(n_577),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_586),
.B(n_580),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_598),
.B(n_599),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_600),
.B(n_593),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_602),
.A2(n_592),
.B(n_591),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_601),
.B(n_587),
.C(n_589),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_604),
.B(n_599),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g608 ( 
.A(n_606),
.B(n_607),
.C(n_603),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_608),
.B(n_605),
.C(n_594),
.Y(n_609)
);

BUFx24_ASAP7_75t_SL g610 ( 
.A(n_609),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_610),
.A2(n_575),
.B(n_571),
.Y(n_611)
);


endmodule