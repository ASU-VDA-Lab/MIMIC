module fake_jpeg_10523_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_49),
.B1(n_37),
.B2(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_57),
.Y(n_78)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_1),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_2),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_3),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_69),
.B1(n_76),
.B2(n_24),
.Y(n_93)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g97 ( 
.A(n_70),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_46),
.B1(n_38),
.B2(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_73),
.B1(n_83),
.B2(n_22),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_79),
.Y(n_87)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_75),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_76)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_23),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_26),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_98),
.Y(n_102)
);

XNOR2x2_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_97),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_103),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_92),
.B1(n_94),
.B2(n_63),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_87),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_64),
.B(n_98),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_84),
.C(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_96),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_72),
.B(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_87),
.Y(n_111)
);

OAI21x1_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_100),
.B(n_89),
.Y(n_112)
);

AOI321xp33_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_95),
.A3(n_86),
.B1(n_93),
.B2(n_67),
.C(n_30),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_95),
.Y(n_114)
);


endmodule