module fake_netlist_5_8_n_1769 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1769);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1769;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_696;
wire n_550;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g163 ( 
.A(n_35),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_63),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_66),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_104),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_58),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_93),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_49),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_85),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_64),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_50),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_7),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_41),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_17),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_111),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_73),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_52),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_37),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_84),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_74),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_18),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_99),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_69),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_105),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_13),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_122),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_109),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_46),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_60),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_62),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_77),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_142),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_108),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_90),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_70),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_13),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_42),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_71),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_88),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_56),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_101),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_161),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_42),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_19),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_94),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_10),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_43),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_151),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_124),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_39),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_144),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_41),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_61),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_98),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_106),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_2),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_32),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_45),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_147),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_53),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_50),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_18),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_10),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_8),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_107),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_33),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_155),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_67),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_33),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_91),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_30),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_0),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_12),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_9),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_112),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_15),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_89),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_126),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_47),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_38),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_20),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_16),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_59),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_128),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_113),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_49),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_40),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_141),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_17),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_15),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_156),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_54),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_114),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_162),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_76),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_36),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_27),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_87),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_131),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_46),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_81),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_51),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_133),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_158),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_118),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_103),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_116),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_75),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_119),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_148),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_135),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_72),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_25),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_95),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_14),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_26),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_14),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_136),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_39),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_127),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_145),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_96),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_8),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_47),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_97),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_43),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_40),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_129),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_32),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_52),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_51),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_80),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_37),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_35),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_79),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_21),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_82),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_57),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_0),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_68),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_6),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_86),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_9),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_160),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_34),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_311),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_182),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_210),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_239),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_210),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_210),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_210),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_210),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_167),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_179),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_187),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_181),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_189),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_196),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_200),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_163),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_168),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_199),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_222),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_163),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_295),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_192),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_218),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_219),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_223),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_174),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_175),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_186),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_228),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_226),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_227),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_230),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_229),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_234),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_243),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_183),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_276),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_269),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_174),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_270),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_299),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_274),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_184),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_197),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_293),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_191),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_301),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_191),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_268),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_235),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_240),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_305),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_231),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_279),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_305),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_323),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_228),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_237),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_237),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_259),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_259),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_320),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_241),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_242),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_312),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_236),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g401 ( 
.A(n_169),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_222),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_320),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_236),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_255),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_255),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_222),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_318),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_326),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_377),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g412 ( 
.A1(n_377),
.A2(n_201),
.B(n_202),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_380),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_326),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_357),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_201),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_341),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_330),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_340),
.A2(n_306),
.B1(n_248),
.B2(n_212),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_371),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_389),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_334),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_401),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_R g429 ( 
.A(n_341),
.B(n_312),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_401),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_344),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_336),
.A2(n_327),
.B1(n_325),
.B2(n_321),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_348),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_342),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_342),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_345),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_394),
.B(n_164),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_201),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_369),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_401),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_396),
.B(n_202),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_403),
.B(n_257),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_357),
.B(n_257),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_401),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_346),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_369),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_400),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_400),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_401),
.B(n_164),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_405),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_405),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_337),
.B(n_165),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_406),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_406),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_355),
.A2(n_388),
.B1(n_364),
.B2(n_373),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_374),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_408),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_339),
.B(n_165),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_328),
.B(n_280),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_408),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_338),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_329),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_361),
.B(n_166),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

OA21x2_ASAP7_75t_L g474 ( 
.A1(n_409),
.A2(n_292),
.B(n_265),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_338),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_362),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_346),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_363),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_367),
.B(n_166),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_368),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_370),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_351),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_372),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_415),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_447),
.B(n_382),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_426),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_447),
.B(n_328),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_415),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_439),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_447),
.B(n_365),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_439),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_417),
.B(n_375),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_447),
.B(n_356),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_419),
.B(n_317),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_351),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_424),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

NAND3xp33_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_353),
.C(n_352),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_413),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_426),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_482),
.B(n_343),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_413),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_470),
.B(n_366),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_426),
.Y(n_507)
);

AND3x2_ASAP7_75t_L g508 ( 
.A(n_471),
.B(n_292),
.C(n_265),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_411),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_417),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_417),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_435),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_435),
.Y(n_516)
);

AND3x2_ASAP7_75t_L g517 ( 
.A(n_471),
.B(n_402),
.C(n_347),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_437),
.B(n_438),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_448),
.B(n_366),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_422),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_422),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_435),
.Y(n_524)
);

AO21x2_ASAP7_75t_L g525 ( 
.A1(n_455),
.A2(n_412),
.B(n_440),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_450),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_435),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_446),
.A2(n_281),
.B1(n_180),
.B2(n_277),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_413),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_425),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_435),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_420),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_452),
.Y(n_539)
);

NOR3xp33_ASAP7_75t_L g540 ( 
.A(n_421),
.B(n_407),
.C(n_331),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_420),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_475),
.A2(n_383),
.B1(n_398),
.B2(n_397),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_482),
.B(n_352),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_465),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_471),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_452),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_425),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_416),
.Y(n_550)
);

BUFx10_ASAP7_75t_L g551 ( 
.A(n_477),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_465),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_448),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_440),
.B(n_399),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_482),
.B(n_353),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_452),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_455),
.B(n_358),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_468),
.B(n_358),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_416),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_416),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_420),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_448),
.Y(n_564)
);

INVxp33_ASAP7_75t_L g565 ( 
.A(n_421),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_468),
.B(n_349),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_461),
.B(n_386),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_441),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_461),
.B(n_359),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_474),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_474),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_453),
.B(n_205),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_452),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_459),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_L g575 ( 
.A(n_467),
.B(n_205),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_441),
.B(n_359),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_416),
.Y(n_577)
);

OA22x2_ASAP7_75t_L g578 ( 
.A1(n_418),
.A2(n_277),
.B1(n_281),
.B2(n_180),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_464),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_474),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_446),
.A2(n_399),
.B1(n_385),
.B2(n_376),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_474),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_459),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_429),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_460),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_460),
.Y(n_587)
);

BUFx6f_ASAP7_75t_SL g588 ( 
.A(n_446),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_460),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_416),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_441),
.B(n_360),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_441),
.B(n_360),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_384),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_453),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_474),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_412),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_423),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_427),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_472),
.B(n_384),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_479),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_479),
.Y(n_601)
);

CKINVDCx6p67_ASAP7_75t_R g602 ( 
.A(n_446),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_423),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_418),
.B(n_378),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_432),
.B(n_397),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_464),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_429),
.Y(n_607)
);

AND3x1_ASAP7_75t_L g608 ( 
.A(n_410),
.B(n_381),
.C(n_379),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_481),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_453),
.B(n_205),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_423),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_418),
.B(n_390),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_412),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_446),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_443),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_445),
.B(n_398),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_423),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_423),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_410),
.B(n_329),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_414),
.B(n_331),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_481),
.Y(n_622)
);

INVx5_ASAP7_75t_L g623 ( 
.A(n_445),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_476),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_445),
.B(n_206),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_R g626 ( 
.A(n_443),
.B(n_170),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_432),
.B(n_280),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_414),
.B(n_350),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_476),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_427),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_478),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_600),
.A2(n_387),
.B1(n_211),
.B2(n_209),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_624),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_628),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_624),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_574),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_566),
.B(n_313),
.C(n_480),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_629),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_600),
.B(n_445),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_601),
.B(n_445),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_520),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_601),
.B(n_205),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_567),
.B(n_480),
.Y(n_644)
);

INVxp33_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_629),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_520),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_564),
.B(n_428),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_559),
.B(n_554),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_505),
.B(n_483),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_578),
.A2(n_205),
.B1(n_221),
.B2(n_273),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_554),
.B(n_428),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_568),
.B(n_428),
.Y(n_653)
);

OAI221xp5_ASAP7_75t_L g654 ( 
.A1(n_529),
.A2(n_490),
.B1(n_493),
.B2(n_582),
.C(n_495),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_585),
.B(n_483),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_578),
.A2(n_307),
.B1(n_221),
.B2(n_273),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_505),
.B(n_315),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_574),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_579),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_576),
.B(n_221),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_591),
.B(n_221),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_569),
.B(n_430),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_630),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_620),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_592),
.B(n_191),
.Y(n_666)
);

NOR2x1_ASAP7_75t_L g667 ( 
.A(n_499),
.B(n_172),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_593),
.B(n_170),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_L g669 ( 
.A(n_617),
.B(n_191),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_596),
.B(n_221),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_584),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_555),
.B(n_171),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_584),
.Y(n_673)
);

OAI221xp5_ASAP7_75t_L g674 ( 
.A1(n_578),
.A2(n_319),
.B1(n_177),
.B2(n_178),
.C(n_185),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_625),
.B(n_430),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_596),
.B(n_273),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_630),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_596),
.B(n_273),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_616),
.B(n_449),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_621),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_632),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_599),
.A2(n_249),
.B1(n_198),
.B2(n_195),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_596),
.B(n_273),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_586),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_492),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_616),
.B(n_449),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_615),
.B(n_449),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_511),
.B(n_473),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_546),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_615),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_515),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_521),
.B(n_261),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_570),
.B(n_456),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_570),
.B(n_456),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_571),
.B(n_581),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_586),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_571),
.B(n_456),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_581),
.B(n_173),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_496),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_583),
.B(n_595),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_583),
.B(n_188),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_596),
.B(n_307),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_595),
.A2(n_307),
.B1(n_191),
.B2(n_244),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_485),
.B(n_171),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_487),
.B(n_176),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_594),
.B(n_213),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_587),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_496),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_522),
.B(n_261),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_587),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_533),
.B(n_261),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_589),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_614),
.B(n_307),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_594),
.B(n_247),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_511),
.B(n_254),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_614),
.B(n_191),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_497),
.Y(n_717)
);

AO22x2_ASAP7_75t_L g718 ( 
.A1(n_627),
.A2(n_256),
.B1(n_285),
.B2(n_286),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_614),
.A2(n_307),
.B1(n_191),
.B2(n_296),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_497),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_484),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_512),
.B(n_288),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_515),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_512),
.B(n_291),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_484),
.B(n_310),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_488),
.B(n_324),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_544),
.B(n_176),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_488),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_492),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_533),
.B(n_431),
.Y(n_730)
);

NAND2x1_ASAP7_75t_L g731 ( 
.A(n_614),
.B(n_427),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_492),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_589),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_607),
.B(n_431),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_604),
.B(n_433),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_557),
.B(n_284),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_604),
.B(n_613),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_613),
.Y(n_738)
);

O2A1O1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_575),
.A2(n_473),
.B(n_469),
.C(n_466),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_609),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_623),
.A2(n_427),
.B(n_466),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_565),
.A2(n_191),
.B1(n_315),
.B2(n_316),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_609),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_612),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_531),
.B(n_427),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_494),
.B(n_433),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_597),
.Y(n_747)
);

O2A1O1Ixp5_ASAP7_75t_L g748 ( 
.A1(n_536),
.A2(n_469),
.B(n_463),
.C(n_462),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_612),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_622),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_536),
.B(n_427),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_538),
.B(n_427),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_597),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_538),
.B(n_434),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_622),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_542),
.B(n_284),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_541),
.B(n_563),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_580),
.A2(n_316),
.B1(n_321),
.B2(n_325),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_541),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_623),
.B(n_190),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_563),
.B(n_434),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_603),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_518),
.B(n_436),
.Y(n_763)
);

BUFx5_ASAP7_75t_L g764 ( 
.A(n_572),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_603),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_513),
.B(n_436),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_560),
.B(n_503),
.Y(n_767)
);

AND2x6_ASAP7_75t_SL g768 ( 
.A(n_489),
.B(n_327),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_606),
.B(n_245),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_626),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_513),
.B(n_442),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_602),
.B(n_287),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_602),
.B(n_605),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_513),
.B(n_519),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_608),
.Y(n_775)
);

INVx3_ASAP7_75t_R g776 ( 
.A(n_489),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_611),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_486),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_611),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_519),
.B(n_442),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_618),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_588),
.A2(n_287),
.B1(n_322),
.B2(n_314),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_486),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_491),
.B(n_250),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_618),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_519),
.B(n_444),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_575),
.A2(n_463),
.B(n_462),
.C(n_458),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_508),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_537),
.B(n_444),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_517),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_537),
.B(n_451),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_588),
.A2(n_540),
.B1(n_525),
.B2(n_504),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_619),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_623),
.B(n_193),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_501),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_623),
.B(n_194),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_537),
.B(n_451),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_759),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_644),
.B(n_525),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_689),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_703),
.A2(n_525),
.B1(n_588),
.B2(n_610),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_644),
.B(n_556),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_740),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_635),
.B(n_526),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_740),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_691),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_649),
.B(n_556),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_668),
.B(n_556),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_703),
.A2(n_610),
.B1(n_572),
.B2(n_507),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_737),
.B(n_526),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_743),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_743),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_690),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_744),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_744),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_750),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_750),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_721),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_728),
.Y(n_819)
);

AND2x2_ASAP7_75t_SL g820 ( 
.A(n_719),
.B(n_514),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_668),
.B(n_561),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_778),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_749),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_692),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_650),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_742),
.A2(n_610),
.B1(n_572),
.B2(n_507),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_665),
.B(n_561),
.Y(n_827)
);

NAND3xp33_ASAP7_75t_SL g828 ( 
.A(n_742),
.B(n_491),
.C(n_545),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_680),
.B(n_561),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_778),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_795),
.Y(n_831)
);

NOR3xp33_ASAP7_75t_SL g832 ( 
.A(n_758),
.B(n_545),
.C(n_553),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_709),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_663),
.B(n_562),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_634),
.B(n_636),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_767),
.A2(n_562),
.B1(n_498),
.B2(n_504),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_690),
.B(n_623),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_685),
.B(n_454),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_690),
.B(n_526),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_755),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_732),
.B(n_454),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_690),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_762),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_765),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_688),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_693),
.A2(n_590),
.B(n_502),
.Y(n_846)
);

AO22x1_ASAP7_75t_L g847 ( 
.A1(n_756),
.A2(n_553),
.B1(n_262),
.B2(n_260),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_792),
.B(n_551),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_777),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_770),
.B(n_551),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_637),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_672),
.B(n_251),
.C(n_258),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_642),
.B(n_551),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_639),
.B(n_498),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_637),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_646),
.B(n_500),
.Y(n_856)
);

NOR2x1p5_ASAP7_75t_L g857 ( 
.A(n_769),
.B(n_252),
.Y(n_857)
);

INVx6_ASAP7_75t_L g858 ( 
.A(n_730),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_723),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_764),
.B(n_502),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_779),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_738),
.B(n_457),
.Y(n_862)
);

BUFx4f_ASAP7_75t_L g863 ( 
.A(n_790),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_781),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_647),
.B(n_500),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_658),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_785),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_764),
.B(n_502),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_793),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_654),
.A2(n_619),
.B1(n_509),
.B2(n_530),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_664),
.B(n_509),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_677),
.B(n_530),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_729),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_735),
.B(n_457),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_681),
.B(n_502),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_688),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_645),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_764),
.B(n_502),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_718),
.A2(n_651),
.B1(n_656),
.B2(n_698),
.Y(n_879)
);

AO22x1_ASAP7_75t_L g880 ( 
.A1(n_756),
.A2(n_283),
.B1(n_253),
.B2(n_266),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_734),
.B(n_590),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_658),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_730),
.Y(n_883)
);

OR2x2_ASAP7_75t_SL g884 ( 
.A(n_784),
.B(n_280),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_699),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_788),
.B(n_458),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_659),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_767),
.A2(n_590),
.B1(n_514),
.B2(n_543),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_708),
.B(n_534),
.Y(n_889)
);

OAI21xp33_ASAP7_75t_L g890 ( 
.A1(n_672),
.A2(n_278),
.B(n_290),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_717),
.B(n_534),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_747),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_720),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_705),
.A2(n_543),
.B1(n_524),
.B2(n_527),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_763),
.B(n_516),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_730),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_764),
.B(n_534),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_659),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_SL g899 ( 
.A(n_758),
.B(n_633),
.C(n_674),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_757),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_705),
.B(n_534),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_711),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_655),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_662),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_662),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_671),
.Y(n_906)
);

BUFx4f_ASAP7_75t_L g907 ( 
.A(n_746),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_753),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_704),
.B(n_534),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_704),
.B(n_577),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_731),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_L g912 ( 
.A(n_764),
.B(n_572),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_640),
.B(n_577),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_764),
.B(n_641),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_695),
.B(n_577),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_727),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_671),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_700),
.B(n_577),
.Y(n_918)
);

O2A1O1Ixp5_ASAP7_75t_L g919 ( 
.A1(n_660),
.A2(n_547),
.B(n_516),
.C(n_524),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_667),
.B(n_527),
.Y(n_920)
);

AOI21x1_ASAP7_75t_L g921 ( 
.A1(n_670),
.A2(n_548),
.B(n_528),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_773),
.B(n_577),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_L g923 ( 
.A(n_772),
.B(n_528),
.Y(n_923)
);

CKINVDCx11_ASAP7_75t_R g924 ( 
.A(n_768),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_753),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_679),
.B(n_631),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_694),
.A2(n_697),
.B(n_652),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_673),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_673),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_684),
.Y(n_930)
);

AND2x4_ASAP7_75t_SL g931 ( 
.A(n_773),
.B(n_532),
.Y(n_931)
);

AO22x1_ASAP7_75t_L g932 ( 
.A1(n_727),
.A2(n_289),
.B1(n_290),
.B2(n_294),
.Y(n_932)
);

BUFx4f_ASAP7_75t_L g933 ( 
.A(n_657),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_696),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_696),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_686),
.B(n_532),
.Y(n_936)
);

NAND2x1_ASAP7_75t_L g937 ( 
.A(n_707),
.B(n_631),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_775),
.B(n_289),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_648),
.B(n_631),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_754),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_718),
.A2(n_610),
.B1(n_572),
.B2(n_501),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_736),
.A2(n_558),
.B1(n_535),
.B2(n_573),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_707),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_736),
.B(n_294),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_653),
.B(n_535),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_772),
.B(n_300),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_718),
.A2(n_610),
.B1(n_572),
.B2(n_573),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_719),
.B(n_539),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_710),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_715),
.B(n_300),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_651),
.A2(n_610),
.B1(n_572),
.B2(n_547),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_675),
.B(n_548),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_687),
.B(n_552),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_656),
.A2(n_552),
.B(n_558),
.C(n_322),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_701),
.A2(n_610),
.B1(n_302),
.B2(n_303),
.Y(n_955)
);

AO22x1_ASAP7_75t_L g956 ( 
.A1(n_638),
.A2(n_314),
.B1(n_304),
.B2(n_303),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_706),
.Y(n_957)
);

AND2x6_ASAP7_75t_SL g958 ( 
.A(n_776),
.B(n_302),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_712),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_722),
.B(n_304),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_643),
.B(n_598),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_783),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_761),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_714),
.B(n_598),
.Y(n_964)
);

INVx2_ASAP7_75t_SL g965 ( 
.A(n_724),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_766),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_733),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_774),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_771),
.B(n_598),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_643),
.B(n_203),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_780),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_748),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_786),
.B(n_506),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_670),
.A2(n_523),
.B(n_510),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_725),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_789),
.Y(n_976)
);

NAND2x1_ASAP7_75t_L g977 ( 
.A(n_745),
.B(n_506),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_782),
.B(n_204),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_791),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_944),
.A2(n_666),
.B(n_669),
.C(n_660),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_900),
.B(n_726),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_927),
.A2(n_678),
.B(n_676),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_944),
.A2(n_796),
.B1(n_794),
.B2(n_760),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_963),
.B(n_682),
.Y(n_984)
);

OAI21xp33_ASAP7_75t_SL g985 ( 
.A1(n_801),
.A2(n_713),
.B(n_702),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_916),
.A2(n_683),
.B(n_676),
.C(n_678),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_SL g987 ( 
.A1(n_946),
.A2(n_881),
.B(n_804),
.C(n_950),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_946),
.A2(n_713),
.B(n_787),
.C(n_661),
.Y(n_988)
);

OAI22xp33_ASAP7_75t_L g989 ( 
.A1(n_907),
.A2(n_797),
.B1(n_796),
.B2(n_794),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_810),
.B(n_760),
.Y(n_990)
);

INVx6_ASAP7_75t_L g991 ( 
.A(n_958),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_803),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_814),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_804),
.B(n_661),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_800),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_848),
.A2(n_899),
.B(n_902),
.C(n_824),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_848),
.A2(n_716),
.B1(n_207),
.B2(n_263),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_978),
.A2(n_739),
.B(n_787),
.C(n_751),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_806),
.B(n_752),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_828),
.B(n_208),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_877),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_881),
.B(n_741),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_890),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_L g1004 ( 
.A(n_978),
.B(n_238),
.C(n_215),
.Y(n_1004)
);

BUFx4f_ASAP7_75t_SL g1005 ( 
.A(n_859),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_825),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_SL g1007 ( 
.A(n_853),
.B(n_214),
.C(n_216),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_850),
.A2(n_1),
.B(n_3),
.C(n_5),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_950),
.A2(n_264),
.B(n_220),
.C(n_224),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_901),
.A2(n_523),
.B(n_510),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_883),
.B(n_100),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_975),
.B(n_940),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_858),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_911),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_960),
.A2(n_272),
.B(n_225),
.C(n_232),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_896),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_903),
.B(n_217),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_940),
.B(n_282),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_832),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_957),
.B(n_233),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_845),
.B(n_275),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_SL g1022 ( 
.A(n_850),
.B(n_246),
.C(n_271),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_858),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_845),
.B(n_523),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_922),
.A2(n_523),
.B(n_510),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_909),
.A2(n_523),
.B(n_510),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_816),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_799),
.B(n_550),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_817),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_883),
.B(n_550),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_805),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_813),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_960),
.A2(n_510),
.B(n_550),
.C(n_506),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_852),
.A2(n_550),
.B(n_506),
.C(n_11),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_910),
.A2(n_550),
.B(n_506),
.Y(n_1035)
);

OAI21xp33_ASAP7_75t_SL g1036 ( 
.A1(n_801),
.A2(n_6),
.B(n_7),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_858),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_876),
.A2(n_506),
.B(n_12),
.C(n_19),
.Y(n_1038)
);

AND2x6_ASAP7_75t_L g1039 ( 
.A(n_966),
.B(n_159),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_873),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_938),
.A2(n_11),
.B(n_20),
.C(n_21),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_811),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_915),
.A2(n_55),
.B(n_152),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_863),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_933),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_815),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_918),
.A2(n_154),
.B(n_143),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_933),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_833),
.B(n_22),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_965),
.B(n_874),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_813),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_863),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_834),
.A2(n_134),
.B(n_121),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_815),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_913),
.A2(n_117),
.B(n_110),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_938),
.B(n_847),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_822),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_818),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_819),
.B(n_22),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_921),
.A2(n_846),
.B(n_919),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_830),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_842),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_842),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_SL g1064 ( 
.A(n_886),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_827),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_839),
.B(n_23),
.C(n_24),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_879),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_971),
.B(n_979),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_874),
.A2(n_102),
.B1(n_83),
.B2(n_78),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_862),
.B(n_65),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_979),
.B(n_28),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_895),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_802),
.B(n_29),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_862),
.A2(n_31),
.B(n_34),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_886),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_873),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_835),
.B(n_36),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_892),
.B(n_44),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_838),
.B(n_44),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_895),
.B(n_45),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_885),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_838),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_879),
.A2(n_48),
.B1(n_951),
.B2(n_809),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_924),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_857),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_841),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_829),
.A2(n_48),
.B(n_839),
.C(n_893),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_841),
.B(n_920),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_970),
.B(n_823),
.Y(n_1089)
);

AO32x1_ASAP7_75t_L g1090 ( 
.A1(n_870),
.A2(n_972),
.A3(n_931),
.B1(n_959),
.B2(n_849),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_SL g1091 ( 
.A(n_954),
.B(n_820),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_798),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_840),
.B(n_923),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_830),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_865),
.B(n_976),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_831),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_865),
.B(n_920),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_976),
.B(n_807),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_964),
.A2(n_808),
.B(n_821),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_968),
.A2(n_869),
.B(n_867),
.C(n_864),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_931),
.A2(n_844),
.B1(n_843),
.B2(n_861),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_951),
.A2(n_809),
.B1(n_954),
.B2(n_820),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_964),
.A2(n_952),
.B(n_945),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_892),
.B(n_908),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_956),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_880),
.B(n_932),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_812),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_962),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_831),
.Y(n_1109)
);

NOR2x1p5_ASAP7_75t_L g1110 ( 
.A(n_884),
.B(n_854),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_836),
.A2(n_856),
.B(n_872),
.C(n_871),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_926),
.A2(n_969),
.B(n_948),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_955),
.A2(n_889),
.B(n_891),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_908),
.Y(n_1114)
);

BUFx12f_ASAP7_75t_L g1115 ( 
.A(n_911),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_875),
.A2(n_953),
.B(n_936),
.C(n_925),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_826),
.A2(n_947),
.B1(n_941),
.B2(n_955),
.Y(n_1117)
);

OAI21xp33_ASAP7_75t_SL g1118 ( 
.A1(n_826),
.A2(n_897),
.B(n_878),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_935),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_967),
.B(n_943),
.Y(n_1120)
);

INVx5_ASAP7_75t_L g1121 ( 
.A(n_1115),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_981),
.B(n_917),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_1005),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_981),
.B(n_917),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1056),
.B(n_888),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1083),
.A2(n_947),
.B1(n_941),
.B2(n_972),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1060),
.A2(n_936),
.B(n_977),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1025),
.A2(n_973),
.B(n_974),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_982),
.A2(n_912),
.B(n_969),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1058),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1082),
.B(n_905),
.Y(n_1131)
);

NAND3x1_ASAP7_75t_L g1132 ( 
.A(n_1106),
.B(n_942),
.C(n_894),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1112),
.A2(n_973),
.B(n_939),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_985),
.A2(n_914),
.B(n_961),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1031),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1014),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1103),
.A2(n_937),
.B(n_851),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1002),
.A2(n_878),
.B(n_860),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1068),
.B(n_904),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1035),
.A2(n_904),
.B(n_855),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1010),
.A2(n_905),
.B(n_866),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1068),
.B(n_906),
.Y(n_1142)
);

BUFx8_ASAP7_75t_L g1143 ( 
.A(n_995),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1026),
.A2(n_906),
.B(n_934),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1088),
.B(n_837),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1044),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1050),
.B(n_928),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_988),
.A2(n_868),
.B(n_949),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_999),
.B(n_928),
.Y(n_1149)
);

AO21x1_ASAP7_75t_L g1150 ( 
.A1(n_994),
.A2(n_868),
.B(n_882),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1116),
.A2(n_882),
.B(n_887),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1028),
.A2(n_887),
.B(n_898),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1028),
.A2(n_929),
.B(n_930),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1108),
.B(n_934),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1048),
.B(n_1040),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1081),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_1001),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_996),
.A2(n_983),
.B(n_1000),
.C(n_987),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1012),
.B(n_1095),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_1033),
.A2(n_1102),
.A3(n_998),
.B(n_980),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1098),
.B(n_984),
.Y(n_1161)
);

NOR4xp25_ASAP7_75t_L g1162 ( 
.A(n_1041),
.B(n_1003),
.C(n_1065),
.D(n_1067),
.Y(n_1162)
);

OAI22x1_ASAP7_75t_L g1163 ( 
.A1(n_1110),
.A2(n_1101),
.B1(n_1105),
.B2(n_1019),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1111),
.A2(n_1014),
.B(n_986),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1118),
.A2(n_1102),
.B(n_1091),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1075),
.B(n_1086),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1087),
.A2(n_1089),
.B(n_1083),
.C(n_1091),
.Y(n_1167)
);

AO31x2_ASAP7_75t_L g1168 ( 
.A1(n_1100),
.A2(n_1117),
.A3(n_1034),
.B(n_1073),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1006),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1088),
.B(n_1076),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1036),
.A2(n_1004),
.B(n_1077),
.C(n_990),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1117),
.A2(n_1073),
.A3(n_1038),
.B(n_1071),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1008),
.A2(n_1074),
.B(n_1113),
.C(n_1059),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1071),
.A2(n_1090),
.A3(n_1043),
.B(n_1047),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_1113),
.A2(n_989),
.B(n_1093),
.C(n_1015),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1088),
.B(n_1076),
.Y(n_1176)
);

O2A1O1Ixp5_ASAP7_75t_L g1177 ( 
.A1(n_1009),
.A2(n_1097),
.B(n_1024),
.C(n_1053),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1119),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1064),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1090),
.A2(n_1054),
.A3(n_1042),
.B(n_1046),
.Y(n_1180)
);

AOI221xp5_ASAP7_75t_SL g1181 ( 
.A1(n_1072),
.A2(n_1080),
.B1(n_992),
.B2(n_993),
.C(n_1027),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1057),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1090),
.A2(n_1055),
.A3(n_1029),
.B(n_1061),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1014),
.Y(n_1184)
);

BUFx10_ASAP7_75t_L g1185 ( 
.A(n_1020),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1092),
.B(n_1018),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1030),
.A2(n_1021),
.B(n_1120),
.Y(n_1187)
);

BUFx2_ASAP7_75t_R g1188 ( 
.A(n_1084),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_SL g1189 ( 
.A(n_1052),
.B(n_1045),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1070),
.A2(n_1079),
.B1(n_1066),
.B2(n_1069),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_1007),
.A2(n_997),
.B(n_1022),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1094),
.A2(n_1096),
.A3(n_1109),
.B(n_1107),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1023),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1040),
.B(n_1070),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1079),
.A2(n_1040),
.B1(n_1011),
.B2(n_1013),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1016),
.B(n_1017),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1049),
.A2(n_1085),
.B(n_1114),
.C(n_1051),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1030),
.A2(n_1104),
.B(n_1051),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1032),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1013),
.B(n_1037),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1062),
.A2(n_1063),
.B(n_1037),
.Y(n_1201)
);

NAND2x1p5_ASAP7_75t_L g1202 ( 
.A(n_1037),
.B(n_1039),
.Y(n_1202)
);

NOR4xp25_ASAP7_75t_L g1203 ( 
.A(n_1078),
.B(n_1041),
.C(n_1003),
.D(n_1065),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_991),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1039),
.A2(n_1060),
.B(n_921),
.Y(n_1205)
);

CKINVDCx11_ASAP7_75t_R g1206 ( 
.A(n_991),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1039),
.A2(n_1060),
.B(n_921),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1039),
.B(n_1068),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1060),
.A2(n_921),
.B(n_1025),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1068),
.B(n_900),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_982),
.A2(n_1103),
.B(n_1099),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_982),
.A2(n_1103),
.B(n_1099),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1060),
.A2(n_921),
.B(n_1025),
.Y(n_1213)
);

AO32x2_ASAP7_75t_L g1214 ( 
.A1(n_1102),
.A2(n_1117),
.A3(n_1083),
.B1(n_870),
.B2(n_633),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1060),
.A2(n_921),
.B(n_1025),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1068),
.B(n_900),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1068),
.B(n_900),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1056),
.A2(n_668),
.B(n_944),
.C(n_566),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1068),
.B(n_900),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1014),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1037),
.Y(n_1221)
);

NAND3xp33_ASAP7_75t_L g1222 ( 
.A(n_1056),
.B(n_944),
.C(n_668),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1056),
.A2(n_565),
.B(n_566),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1001),
.B(n_642),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_995),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1068),
.B(n_900),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1060),
.A2(n_921),
.B(n_1025),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1083),
.A2(n_879),
.B1(n_801),
.B2(n_1117),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1082),
.B(n_635),
.Y(n_1229)
);

OR2x6_ASAP7_75t_L g1230 ( 
.A(n_1088),
.B(n_1115),
.Y(n_1230)
);

AO21x1_ASAP7_75t_L g1231 ( 
.A1(n_994),
.A2(n_1091),
.B(n_944),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_982),
.A2(n_1025),
.B(n_1028),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1060),
.A2(n_921),
.B(n_1025),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_981),
.B(n_635),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1058),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1014),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_SL g1237 ( 
.A1(n_996),
.A2(n_1068),
.B(n_1071),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_982),
.A2(n_1103),
.B(n_1099),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1005),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_985),
.A2(n_1112),
.B(n_988),
.Y(n_1240)
);

AOI221x1_ASAP7_75t_L g1241 ( 
.A1(n_1067),
.A2(n_944),
.B1(n_1056),
.B2(n_668),
.C(n_982),
.Y(n_1241)
);

AOI21x1_ASAP7_75t_L g1242 ( 
.A1(n_982),
.A2(n_1025),
.B(n_1028),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_982),
.A2(n_1103),
.B(n_1099),
.Y(n_1243)
);

AO21x1_ASAP7_75t_L g1244 ( 
.A1(n_994),
.A2(n_1091),
.B(n_944),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1058),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1056),
.A2(n_668),
.B(n_944),
.C(n_566),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_981),
.B(n_635),
.Y(n_1247)
);

OA22x2_ASAP7_75t_L g1248 ( 
.A1(n_1074),
.A2(n_627),
.B1(n_432),
.B2(n_605),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_982),
.A2(n_1103),
.B(n_1099),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_981),
.B(n_635),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1082),
.B(n_635),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_995),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_981),
.B(n_635),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1058),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_985),
.A2(n_1112),
.B(n_988),
.Y(n_1255)
);

O2A1O1Ixp5_ASAP7_75t_L g1256 ( 
.A1(n_1056),
.A2(n_944),
.B(n_668),
.C(n_946),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1001),
.B(n_642),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_981),
.B(n_635),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1083),
.A2(n_1111),
.B(n_1117),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_985),
.A2(n_1112),
.B(n_988),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1001),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1083),
.A2(n_879),
.B1(n_801),
.B2(n_1117),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_982),
.A2(n_1103),
.B(n_1099),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1005),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_982),
.A2(n_1103),
.B(n_1099),
.Y(n_1265)
);

INVx6_ASAP7_75t_L g1266 ( 
.A(n_1121),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1206),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1130),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1145),
.B(n_1170),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1127),
.A2(n_1153),
.B(n_1152),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1256),
.A2(n_1246),
.B(n_1218),
.Y(n_1271)
);

AOI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1164),
.A2(n_1125),
.B(n_1232),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1223),
.A2(n_1222),
.B1(n_1190),
.B2(n_1163),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1123),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_SL g1275 ( 
.A1(n_1173),
.A2(n_1158),
.B(n_1167),
.C(n_1262),
.Y(n_1275)
);

AOI222xp33_ASAP7_75t_L g1276 ( 
.A1(n_1223),
.A2(n_1262),
.B1(n_1228),
.B2(n_1222),
.C1(n_1165),
.C2(n_1190),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_SL g1277 ( 
.A(n_1188),
.B(n_1239),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1156),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1264),
.Y(n_1279)
);

NOR2xp67_ASAP7_75t_L g1280 ( 
.A(n_1157),
.B(n_1261),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1211),
.A2(n_1238),
.B(n_1212),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1192),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1213),
.A2(n_1227),
.B(n_1215),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1234),
.B(n_1247),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_1143),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1231),
.A2(n_1244),
.A3(n_1150),
.B(n_1241),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1175),
.A2(n_1171),
.B(n_1177),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1131),
.B(n_1229),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1240),
.A2(n_1255),
.B(n_1260),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1151),
.Y(n_1290)
);

CKINVDCx16_ASAP7_75t_R g1291 ( 
.A(n_1204),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1240),
.A2(n_1255),
.B(n_1260),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1235),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1145),
.B(n_1170),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1243),
.A2(n_1265),
.A3(n_1249),
.B(n_1263),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1245),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1259),
.A2(n_1129),
.B(n_1228),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1165),
.A2(n_1233),
.B(n_1133),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1121),
.B(n_1136),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1141),
.A2(n_1144),
.B(n_1140),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1176),
.B(n_1230),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1254),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1242),
.A2(n_1128),
.B(n_1137),
.Y(n_1303)
);

NOR3xp33_ASAP7_75t_L g1304 ( 
.A(n_1186),
.B(n_1197),
.C(n_1258),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1138),
.A2(n_1219),
.B(n_1226),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1185),
.Y(n_1306)
);

BUFx12f_ASAP7_75t_L g1307 ( 
.A(n_1143),
.Y(n_1307)
);

AOI22x1_ASAP7_75t_L g1308 ( 
.A1(n_1237),
.A2(n_1187),
.B1(n_1202),
.B2(n_1198),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1178),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1210),
.A2(n_1226),
.B(n_1219),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1250),
.B(n_1253),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1210),
.A2(n_1216),
.B(n_1217),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1251),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1203),
.A2(n_1132),
.B(n_1161),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1172),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1134),
.A2(n_1148),
.B(n_1181),
.Y(n_1316)
);

OR2x6_ASAP7_75t_L g1317 ( 
.A(n_1202),
.B(n_1230),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1225),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1126),
.A2(n_1208),
.B(n_1122),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1159),
.B(n_1166),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1135),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1195),
.A2(n_1248),
.B1(n_1194),
.B2(n_1196),
.Y(n_1323)
);

BUFx2_ASAP7_75t_R g1324 ( 
.A(n_1252),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1191),
.A2(n_1126),
.B1(n_1149),
.B2(n_1195),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_L g1326 ( 
.A(n_1203),
.B(n_1162),
.C(n_1181),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1139),
.A2(n_1142),
.B(n_1124),
.Y(n_1327)
);

AO31x2_ASAP7_75t_L g1328 ( 
.A1(n_1139),
.A2(n_1174),
.A3(n_1160),
.B(n_1214),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1169),
.B(n_1154),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1182),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1200),
.Y(n_1331)
);

NOR2xp67_ASAP7_75t_L g1332 ( 
.A(n_1224),
.B(n_1257),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1179),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1147),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1162),
.A2(n_1191),
.B(n_1201),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1221),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1230),
.B(n_1155),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1199),
.A2(n_1236),
.B(n_1220),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_1221),
.Y(n_1339)
);

BUFx12f_ASAP7_75t_L g1340 ( 
.A(n_1121),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1174),
.A2(n_1160),
.A3(n_1214),
.B(n_1183),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1189),
.B(n_1146),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1184),
.B(n_1214),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1168),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1183),
.A2(n_1174),
.B(n_1180),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1168),
.A2(n_1255),
.B(n_1240),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1168),
.A2(n_1256),
.B(n_1246),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1180),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1180),
.A2(n_1207),
.B(n_1205),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1222),
.A2(n_944),
.B1(n_1248),
.B2(n_1056),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1222),
.A2(n_944),
.B1(n_1248),
.B2(n_1056),
.Y(n_1351)
);

OR2x6_ASAP7_75t_L g1352 ( 
.A(n_1259),
.B(n_1202),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1259),
.B(n_1202),
.Y(n_1353)
);

AOI22x1_ASAP7_75t_L g1354 ( 
.A1(n_1237),
.A2(n_665),
.B1(n_680),
.B2(n_1110),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1228),
.A2(n_1262),
.B1(n_1248),
.B2(n_1223),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1211),
.A2(n_1238),
.B(n_1212),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1192),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1256),
.A2(n_1246),
.B(n_1218),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1209),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1123),
.Y(n_1360)
);

OAI211xp5_ASAP7_75t_L g1361 ( 
.A1(n_1218),
.A2(n_1246),
.B(n_1223),
.C(n_566),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1209),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1192),
.Y(n_1363)
);

CKINVDCx16_ASAP7_75t_R g1364 ( 
.A(n_1239),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_1206),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1209),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1256),
.A2(n_1246),
.B(n_1218),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1193),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1209),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1172),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1218),
.B(n_1246),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1123),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1130),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1130),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1121),
.B(n_1014),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1130),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1240),
.A2(n_1255),
.B(n_1260),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1234),
.B(n_1247),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1130),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1211),
.A2(n_1238),
.B(n_1212),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1172),
.Y(n_1381)
);

CKINVDCx9p33_ASAP7_75t_R g1382 ( 
.A(n_1234),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1193),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1193),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1209),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1205),
.A2(n_1207),
.B(n_1209),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1131),
.B(n_1229),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1240),
.A2(n_1255),
.B(n_1260),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1297),
.A2(n_1356),
.B(n_1281),
.Y(n_1389)
);

O2A1O1Ixp5_ASAP7_75t_L g1390 ( 
.A1(n_1361),
.A2(n_1371),
.B(n_1367),
.C(n_1358),
.Y(n_1390)
);

INVxp67_ASAP7_75t_L g1391 ( 
.A(n_1313),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1365),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1329),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1371),
.A2(n_1273),
.B(n_1350),
.C(n_1351),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1284),
.B(n_1311),
.Y(n_1395)
);

AOI211xp5_ASAP7_75t_L g1396 ( 
.A1(n_1271),
.A2(n_1355),
.B(n_1275),
.C(n_1314),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1310),
.A2(n_1312),
.B(n_1352),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1350),
.A2(n_1351),
.B(n_1287),
.C(n_1326),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1355),
.A2(n_1319),
.B1(n_1378),
.B2(n_1292),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1268),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1332),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1289),
.A2(n_1388),
.B1(n_1292),
.B2(n_1377),
.Y(n_1402)
);

CKINVDCx6p67_ASAP7_75t_R g1403 ( 
.A(n_1365),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1275),
.A2(n_1304),
.B(n_1347),
.C(n_1276),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1320),
.B(n_1305),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1323),
.B(n_1278),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1342),
.A2(n_1325),
.B(n_1301),
.C(n_1334),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1339),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1293),
.B(n_1296),
.Y(n_1409)
);

AOI211xp5_ASAP7_75t_L g1410 ( 
.A1(n_1342),
.A2(n_1280),
.B(n_1333),
.C(n_1382),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1302),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1269),
.B(n_1294),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1289),
.A2(n_1388),
.B1(n_1292),
.B2(n_1377),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1352),
.A2(n_1353),
.B(n_1377),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1337),
.A2(n_1317),
.B(n_1309),
.C(n_1379),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1317),
.B(n_1337),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1289),
.A2(n_1388),
.B1(n_1325),
.B2(n_1346),
.Y(n_1418)
);

AOI221x1_ASAP7_75t_SL g1419 ( 
.A1(n_1376),
.A2(n_1382),
.B1(n_1343),
.B2(n_1322),
.C(n_1330),
.Y(n_1419)
);

O2A1O1Ixp5_ASAP7_75t_L g1420 ( 
.A1(n_1272),
.A2(n_1344),
.B(n_1343),
.C(n_1380),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1346),
.A2(n_1352),
.B1(n_1353),
.B2(n_1337),
.Y(n_1421)
);

NOR2xp67_ASAP7_75t_L g1422 ( 
.A(n_1274),
.B(n_1360),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1353),
.A2(n_1375),
.B(n_1317),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1346),
.A2(n_1308),
.B(n_1316),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1291),
.Y(n_1425)
);

BUFx12f_ASAP7_75t_L g1426 ( 
.A(n_1267),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1267),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1335),
.A2(n_1315),
.B(n_1370),
.C(n_1381),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1354),
.A2(n_1316),
.B1(n_1327),
.B2(n_1266),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1349),
.A2(n_1303),
.B(n_1270),
.Y(n_1430)
);

AOI21x1_ASAP7_75t_SL g1431 ( 
.A1(n_1306),
.A2(n_1340),
.B(n_1324),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1336),
.B(n_1338),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1433)
);

OA22x2_ASAP7_75t_L g1434 ( 
.A1(n_1368),
.A2(n_1384),
.B1(n_1372),
.B2(n_1344),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1383),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1383),
.B(n_1286),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1336),
.B(n_1299),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1279),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1364),
.B(n_1266),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1339),
.B(n_1277),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1298),
.A2(n_1363),
.B(n_1282),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1375),
.A2(n_1298),
.B(n_1363),
.Y(n_1443)
);

O2A1O1Ixp5_ASAP7_75t_L g1444 ( 
.A1(n_1290),
.A2(n_1357),
.B(n_1348),
.C(n_1295),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1285),
.A2(n_1357),
.B1(n_1348),
.B2(n_1318),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1341),
.B(n_1295),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1341),
.B(n_1345),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1290),
.A2(n_1318),
.B(n_1307),
.C(n_1295),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1359),
.A2(n_1362),
.B(n_1366),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1366),
.A2(n_1369),
.B1(n_1385),
.B2(n_1386),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1369),
.A2(n_1287),
.B(n_1300),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1283),
.B(n_1310),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1283),
.B(n_1321),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1310),
.B(n_1312),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1361),
.A2(n_1246),
.B(n_1218),
.C(n_1256),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1297),
.A2(n_1246),
.B(n_1218),
.Y(n_1456)
);

OAI211xp5_ASAP7_75t_L g1457 ( 
.A1(n_1350),
.A2(n_1246),
.B(n_1218),
.C(n_1223),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1297),
.A2(n_1246),
.B(n_1218),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1291),
.Y(n_1459)
);

O2A1O1Ixp5_ASAP7_75t_L g1460 ( 
.A1(n_1361),
.A2(n_1256),
.B(n_1371),
.C(n_1358),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1310),
.B(n_1312),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1288),
.B(n_1387),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1321),
.B(n_1331),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1371),
.A2(n_1218),
.B(n_1246),
.C(n_1056),
.Y(n_1464)
);

AOI221xp5_ASAP7_75t_L g1465 ( 
.A1(n_1355),
.A2(n_1246),
.B1(n_1218),
.B2(n_1275),
.C(n_1223),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1268),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1350),
.A2(n_1262),
.B1(n_1228),
.B2(n_1351),
.Y(n_1467)
);

INVx5_ASAP7_75t_L g1468 ( 
.A(n_1447),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1399),
.B(n_1454),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1418),
.B(n_1402),
.Y(n_1470)
);

AO21x1_ASAP7_75t_SL g1471 ( 
.A1(n_1454),
.A2(n_1461),
.B(n_1405),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1461),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1397),
.B(n_1414),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1453),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1413),
.B(n_1446),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1400),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1416),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1433),
.B(n_1438),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1449),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1465),
.A2(n_1467),
.B1(n_1458),
.B2(n_1456),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1424),
.A2(n_1389),
.B(n_1442),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1436),
.B(n_1444),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1443),
.B(n_1423),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1430),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1432),
.B(n_1405),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1420),
.A2(n_1452),
.B(n_1460),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1429),
.A2(n_1464),
.B(n_1450),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1451),
.B(n_1466),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1428),
.A2(n_1398),
.B(n_1394),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1411),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1399),
.B(n_1395),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1409),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1451),
.B(n_1406),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1421),
.B(n_1404),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1417),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1393),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1455),
.A2(n_1465),
.B(n_1448),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1415),
.B(n_1467),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1434),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1434),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1419),
.Y(n_1501)
);

NOR2x1_ASAP7_75t_L g1502 ( 
.A(n_1457),
.B(n_1407),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1396),
.B(n_1390),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1419),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1401),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1471),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1476),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1472),
.B(n_1463),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1472),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1470),
.B(n_1445),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1470),
.B(n_1445),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1488),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1485),
.B(n_1412),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1478),
.B(n_1391),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1478),
.B(n_1435),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1473),
.A2(n_1480),
.B(n_1497),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1493),
.B(n_1462),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1485),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1485),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1491),
.B(n_1410),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1474),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1493),
.B(n_1439),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1491),
.B(n_1440),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1469),
.B(n_1437),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1479),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1493),
.B(n_1459),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1474),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1522),
.Y(n_1528)
);

AOI211xp5_ASAP7_75t_L g1529 ( 
.A1(n_1516),
.A2(n_1503),
.B(n_1501),
.C(n_1504),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1516),
.A2(n_1502),
.B1(n_1503),
.B2(n_1480),
.Y(n_1530)
);

OAI222xp33_ASAP7_75t_L g1531 ( 
.A1(n_1520),
.A2(n_1502),
.B1(n_1503),
.B2(n_1498),
.C1(n_1494),
.C2(n_1501),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1520),
.A2(n_1489),
.B1(n_1498),
.B2(n_1494),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1518),
.B(n_1485),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1526),
.Y(n_1534)
);

AOI322xp5_ASAP7_75t_L g1535 ( 
.A1(n_1510),
.A2(n_1504),
.A3(n_1469),
.B1(n_1499),
.B2(n_1500),
.C1(n_1482),
.C2(n_1475),
.Y(n_1535)
);

AOI221xp5_ASAP7_75t_L g1536 ( 
.A1(n_1523),
.A2(n_1489),
.B1(n_1496),
.B2(n_1490),
.C(n_1482),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1518),
.B(n_1485),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1521),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_SL g1539 ( 
.A(n_1506),
.B(n_1473),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1525),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1523),
.A2(n_1498),
.B1(n_1494),
.B2(n_1500),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1518),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1519),
.B(n_1468),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1526),
.B(n_1498),
.C(n_1494),
.Y(n_1544)
);

AND2x4_ASAP7_75t_SL g1545 ( 
.A(n_1513),
.B(n_1483),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1524),
.A2(n_1489),
.B1(n_1498),
.B2(n_1494),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1519),
.B(n_1468),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_R g1548 ( 
.A(n_1526),
.B(n_1392),
.Y(n_1548)
);

OAI211xp5_ASAP7_75t_L g1549 ( 
.A1(n_1510),
.A2(n_1482),
.B(n_1496),
.C(n_1500),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1522),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1524),
.A2(n_1498),
.B1(n_1494),
.B2(n_1500),
.Y(n_1551)
);

AO22x1_ASAP7_75t_L g1552 ( 
.A1(n_1509),
.A2(n_1505),
.B1(n_1499),
.B2(n_1511),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1519),
.B(n_1468),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1510),
.A2(n_1489),
.B1(n_1498),
.B2(n_1494),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1511),
.A2(n_1473),
.B1(n_1477),
.B2(n_1499),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1521),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1517),
.B(n_1515),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1512),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1517),
.A2(n_1473),
.B1(n_1483),
.B2(n_1477),
.Y(n_1559)
);

AOI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1511),
.A2(n_1490),
.B1(n_1505),
.B2(n_1495),
.C(n_1492),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1507),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1514),
.A2(n_1473),
.B1(n_1483),
.B2(n_1477),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1508),
.A2(n_1505),
.B1(n_1492),
.B2(n_1495),
.C(n_1527),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1561),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1534),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1540),
.Y(n_1566)
);

INVx4_ASAP7_75t_L g1567 ( 
.A(n_1545),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1534),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1561),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1538),
.Y(n_1570)
);

BUFx8_ASAP7_75t_L g1571 ( 
.A(n_1549),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1532),
.B(n_1506),
.Y(n_1572)
);

NAND3xp33_ASAP7_75t_L g1573 ( 
.A(n_1530),
.B(n_1486),
.C(n_1473),
.Y(n_1573)
);

BUFx8_ASAP7_75t_L g1574 ( 
.A(n_1542),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1540),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1556),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1556),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1558),
.Y(n_1578)
);

INVx2_ASAP7_75t_SL g1579 ( 
.A(n_1543),
.Y(n_1579)
);

NOR2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1544),
.B(n_1403),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1534),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1557),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1547),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1528),
.Y(n_1584)
);

NAND2xp33_ASAP7_75t_R g1585 ( 
.A(n_1531),
.B(n_1483),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1550),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1530),
.B(n_1486),
.C(n_1514),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1483),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1552),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1536),
.A2(n_1481),
.B(n_1484),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1564),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1581),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1584),
.B(n_1563),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1584),
.B(n_1560),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1586),
.B(n_1529),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1565),
.Y(n_1596)
);

AND2x2_ASAP7_75t_SL g1597 ( 
.A(n_1565),
.B(n_1554),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1564),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1569),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1569),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1570),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1566),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1571),
.B(n_1529),
.Y(n_1603)
);

OAI211xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1572),
.A2(n_1535),
.B(n_1546),
.C(n_1514),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1579),
.B(n_1539),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1587),
.A2(n_1544),
.B(n_1535),
.Y(n_1606)
);

NAND2x1_ASAP7_75t_L g1607 ( 
.A(n_1588),
.B(n_1553),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1581),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1579),
.B(n_1539),
.Y(n_1609)
);

INVx3_ASAP7_75t_SL g1610 ( 
.A(n_1572),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1566),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1566),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1579),
.B(n_1553),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1571),
.B(n_1506),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1570),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1583),
.B(n_1533),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1583),
.B(n_1533),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1567),
.B(n_1426),
.Y(n_1618)
);

NAND4xp25_ASAP7_75t_L g1619 ( 
.A(n_1587),
.B(n_1548),
.C(n_1551),
.D(n_1541),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1573),
.A2(n_1562),
.B(n_1559),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1577),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1575),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1589),
.B(n_1537),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1586),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1577),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1574),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1578),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1575),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1618),
.B(n_1427),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1626),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1624),
.B(n_1589),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1591),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1626),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1610),
.B(n_1626),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1591),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1592),
.B(n_1568),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1628),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1610),
.B(n_1623),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1598),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1608),
.B(n_1568),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1598),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1603),
.B(n_1580),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1599),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1610),
.A2(n_1573),
.B1(n_1580),
.B2(n_1555),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1596),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1627),
.B(n_1567),
.Y(n_1646)
);

OAI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1606),
.A2(n_1588),
.B(n_1576),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1623),
.B(n_1567),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1597),
.A2(n_1619),
.B(n_1604),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1595),
.B(n_1576),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1614),
.B(n_1567),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1605),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1599),
.Y(n_1653)
);

AOI21xp33_ASAP7_75t_L g1654 ( 
.A1(n_1597),
.A2(n_1585),
.B(n_1571),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1600),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1600),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1605),
.B(n_1567),
.Y(n_1657)
);

OAI21xp33_ASAP7_75t_L g1658 ( 
.A1(n_1597),
.A2(n_1588),
.B(n_1576),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1602),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1601),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1602),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1593),
.A2(n_1585),
.B1(n_1571),
.B2(n_1487),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1627),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1594),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1663),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1633),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1638),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1638),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1631),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1635),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1633),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1634),
.B(n_1609),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1664),
.B(n_1624),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1648),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1634),
.Y(n_1675)
);

NAND2x1_ASAP7_75t_L g1676 ( 
.A(n_1651),
.B(n_1609),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1635),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1639),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1631),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1639),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1645),
.B(n_1601),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1636),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1630),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1640),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1652),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1641),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1652),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1648),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1649),
.B(n_1616),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1641),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1669),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1668),
.B(n_1650),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1669),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1672),
.B(n_1642),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1683),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1675),
.B(n_1630),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1689),
.A2(n_1647),
.B1(n_1658),
.B2(n_1662),
.C(n_1632),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1675),
.B(n_1646),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1676),
.A2(n_1642),
.B1(n_1644),
.B2(n_1654),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1668),
.B(n_1667),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1683),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1679),
.B(n_1684),
.Y(n_1703)
);

AOI32xp33_ASAP7_75t_L g1704 ( 
.A1(n_1679),
.A2(n_1657),
.A3(n_1646),
.B1(n_1613),
.B2(n_1617),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1672),
.B(n_1642),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1682),
.A2(n_1620),
.B1(n_1571),
.B2(n_1646),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1690),
.Y(n_1707)
);

OAI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1684),
.A2(n_1588),
.B1(n_1607),
.B2(n_1590),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1670),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1666),
.B(n_1657),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1696),
.B(n_1666),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1701),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1702),
.B(n_1666),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1694),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1699),
.B(n_1671),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1691),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1697),
.B(n_1671),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1693),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_R g1719 ( 
.A(n_1705),
.B(n_1674),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1703),
.B(n_1671),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1710),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1692),
.B(n_1685),
.Y(n_1722)
);

NOR2x1_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1665),
.Y(n_1723)
);

AOI222xp33_ASAP7_75t_L g1724 ( 
.A1(n_1721),
.A2(n_1700),
.B1(n_1706),
.B2(n_1673),
.C1(n_1665),
.C2(n_1681),
.Y(n_1724)
);

OAI211xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1720),
.A2(n_1704),
.B(n_1706),
.C(n_1698),
.Y(n_1725)
);

OAI211xp5_ASAP7_75t_L g1726 ( 
.A1(n_1723),
.A2(n_1698),
.B(n_1676),
.C(n_1681),
.Y(n_1726)
);

NOR4xp25_ASAP7_75t_L g1727 ( 
.A(n_1721),
.B(n_1709),
.C(n_1707),
.D(n_1687),
.Y(n_1727)
);

AOI211xp5_ASAP7_75t_SL g1728 ( 
.A1(n_1711),
.A2(n_1708),
.B(n_1687),
.C(n_1688),
.Y(n_1728)
);

NOR3xp33_ASAP7_75t_L g1729 ( 
.A(n_1717),
.B(n_1687),
.C(n_1674),
.Y(n_1729)
);

NAND4xp25_ASAP7_75t_SL g1730 ( 
.A(n_1715),
.B(n_1688),
.C(n_1690),
.D(n_1670),
.Y(n_1730)
);

NOR3xp33_ASAP7_75t_L g1731 ( 
.A(n_1713),
.B(n_1688),
.C(n_1629),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1714),
.A2(n_1708),
.B1(n_1655),
.B2(n_1607),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1722),
.A2(n_1678),
.B(n_1677),
.Y(n_1733)
);

NOR3xp33_ASAP7_75t_L g1734 ( 
.A(n_1712),
.B(n_1686),
.C(n_1678),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1732),
.Y(n_1735)
);

AOI21xp33_ASAP7_75t_SL g1736 ( 
.A1(n_1726),
.A2(n_1718),
.B(n_1716),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1734),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1733),
.B(n_1677),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1730),
.Y(n_1739)
);

AOI32xp33_ASAP7_75t_L g1740 ( 
.A1(n_1725),
.A2(n_1719),
.A3(n_1686),
.B1(n_1680),
.B2(n_1656),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1724),
.B1(n_1728),
.B2(n_1727),
.C(n_1729),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1737),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1739),
.Y(n_1743)
);

NOR2x1_ASAP7_75t_L g1744 ( 
.A(n_1735),
.B(n_1680),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1736),
.B(n_1731),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1738),
.B(n_1637),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1739),
.Y(n_1747)
);

XNOR2xp5_ASAP7_75t_L g1748 ( 
.A(n_1741),
.B(n_1425),
.Y(n_1748)
);

NOR3xp33_ASAP7_75t_L g1749 ( 
.A(n_1745),
.B(n_1653),
.C(n_1643),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1747),
.A2(n_1660),
.B1(n_1643),
.B2(n_1656),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1744),
.B(n_1653),
.Y(n_1751)
);

NAND2x1_ASAP7_75t_SL g1752 ( 
.A(n_1742),
.B(n_1660),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1752),
.Y(n_1753)
);

NOR3xp33_ASAP7_75t_L g1754 ( 
.A(n_1749),
.B(n_1743),
.C(n_1746),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1748),
.Y(n_1755)
);

NOR3x2_ASAP7_75t_L g1756 ( 
.A(n_1754),
.B(n_1751),
.C(n_1750),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1756),
.A2(n_1755),
.B1(n_1753),
.B2(n_1637),
.C(n_1661),
.Y(n_1757)
);

OR3x1_ASAP7_75t_L g1758 ( 
.A(n_1757),
.B(n_1621),
.C(n_1615),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1757),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1759),
.B(n_1661),
.Y(n_1760)
);

INVxp67_ASAP7_75t_L g1761 ( 
.A(n_1758),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1659),
.B1(n_1611),
.B2(n_1628),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1760),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1659),
.B1(n_1622),
.B2(n_1612),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1762),
.B1(n_1612),
.B2(n_1611),
.Y(n_1765)
);

OR2x6_ASAP7_75t_L g1766 ( 
.A(n_1765),
.B(n_1422),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1625),
.B1(n_1615),
.B2(n_1621),
.Y(n_1767)
);

AOI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1625),
.B1(n_1622),
.B2(n_1408),
.C(n_1613),
.Y(n_1768)
);

AOI211xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1408),
.B(n_1441),
.C(n_1431),
.Y(n_1769)
);


endmodule