module fake_jpeg_3547_n_686 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_686);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_686;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_461;
wire n_214;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx8_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_40),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_63),
.A2(n_65),
.B(n_80),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_1),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_66),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_67),
.Y(n_160)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g224 ( 
.A(n_68),
.Y(n_224)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_69),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_86),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_19),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_74),
.B(n_106),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx5_ASAP7_75t_SL g76 ( 
.A(n_50),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_76),
.B(n_59),
.Y(n_153)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_79),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_33),
.B(n_1),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_84),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_32),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_89),
.Y(n_189)
);

BUFx16f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_90),
.Y(n_227)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_91),
.Y(n_197)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_93),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_95),
.Y(n_207)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_56),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_100),
.B(n_104),
.Y(n_174)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_56),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_19),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_111),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_47),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_121),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_24),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_21),
.Y(n_122)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_21),
.Y(n_124)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_23),
.Y(n_126)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_126),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

CKINVDCx12_ASAP7_75t_R g186 ( 
.A(n_127),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_23),
.Y(n_128)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_29),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_29),
.Y(n_130)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_29),
.Y(n_131)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_131),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_39),
.Y(n_132)
);

BUFx4f_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_65),
.B(n_80),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_140),
.B(n_151),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_147),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_119),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_153),
.Y(n_264)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_99),
.A2(n_26),
.B1(n_58),
.B2(n_30),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_165),
.A2(n_180),
.B1(n_35),
.B2(n_53),
.Y(n_249)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_167),
.Y(n_247)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_63),
.B(n_46),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_176),
.B(n_179),
.Y(n_232)
);

INVx2_ASAP7_75t_R g178 ( 
.A(n_76),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_178),
.A2(n_185),
.B(n_205),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_112),
.B(n_59),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_60),
.A2(n_26),
.B1(n_58),
.B2(n_30),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_130),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_212),
.Y(n_242)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_182),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_102),
.B(n_46),
.Y(n_185)
);

BUFx4f_ASAP7_75t_L g188 ( 
.A(n_79),
.Y(n_188)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_191),
.Y(n_279)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_192),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_51),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_208),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_103),
.B(n_105),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_81),
.B(n_59),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_206),
.B(n_228),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_111),
.B(n_41),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_115),
.B(n_41),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_209),
.B(n_215),
.Y(n_288)
);

OA22x2_ASAP7_75t_SL g210 ( 
.A1(n_91),
.A2(n_45),
.B1(n_54),
.B2(n_51),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_210),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_277)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_127),
.Y(n_211)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_211),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_116),
.B(n_34),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_64),
.B(n_34),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_67),
.B(n_55),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_219),
.B(n_222),
.Y(n_289)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_96),
.Y(n_220)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_220),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_78),
.B(n_55),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_82),
.B(n_54),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_38),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_85),
.B(n_38),
.Y(n_228)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_233),
.Y(n_355)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_234),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_134),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_235),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_236),
.B(n_270),
.Y(n_332)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_239),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_134),
.Y(n_240)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_240),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_139),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_241),
.Y(n_364)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_162),
.Y(n_243)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_243),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_35),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_244),
.B(n_260),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_245),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_143),
.B(n_93),
.C(n_89),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_248),
.B(n_292),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_249),
.A2(n_255),
.B1(n_273),
.B2(n_275),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_137),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_250),
.B(n_280),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_212),
.A2(n_57),
.B1(n_53),
.B2(n_39),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_252),
.A2(n_272),
.B1(n_293),
.B2(n_298),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_148),
.Y(n_253)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_253),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_180),
.A2(n_210),
.B1(n_193),
.B2(n_206),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_258),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_178),
.B(n_57),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_259),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_187),
.B(n_57),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_153),
.A2(n_53),
.B(n_39),
.C(n_45),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_261),
.A2(n_303),
.B(n_216),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_262),
.Y(n_342)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_160),
.Y(n_263)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_263),
.Y(n_357)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_171),
.Y(n_265)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_265),
.Y(n_328)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_163),
.Y(n_267)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_141),
.B(n_1),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_268),
.B(n_271),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_179),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_291),
.B1(n_224),
.B2(n_223),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_174),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_174),
.B(n_1),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_184),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_193),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_169),
.Y(n_274)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_222),
.A2(n_226),
.B1(n_199),
.B2(n_229),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_161),
.Y(n_276)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_277),
.B(n_296),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_190),
.Y(n_278)
);

CKINVDCx6p67_ASAP7_75t_R g344 ( 
.A(n_278),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_185),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_190),
.Y(n_282)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_194),
.B(n_6),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_283),
.B(n_295),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_217),
.B(n_6),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_284),
.B(n_307),
.Y(n_371)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_162),
.Y(n_285)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_145),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_286),
.Y(n_373)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_138),
.Y(n_287)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_287),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_177),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_290),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_209),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_136),
.B(n_7),
.C(n_10),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_184),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_200),
.B(n_11),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_225),
.B(n_19),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_137),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_297),
.B(n_299),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_230),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_208),
.B(n_12),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_195),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_300),
.Y(n_323)
);

INVx11_ASAP7_75t_L g301 ( 
.A(n_203),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_301),
.A2(n_312),
.B1(n_313),
.B2(n_186),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_213),
.A2(n_12),
.B(n_16),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_177),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_304),
.Y(n_327)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_146),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_305),
.B(n_311),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_133),
.B(n_16),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_172),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_308),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_166),
.A2(n_17),
.B1(n_18),
.B2(n_157),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_205),
.Y(n_335)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_149),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_223),
.A2(n_18),
.B1(n_224),
.B2(n_188),
.Y(n_312)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_204),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_L g402 ( 
.A1(n_316),
.A2(n_317),
.B(n_335),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_288),
.B(n_150),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_322),
.B(n_354),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_237),
.B(n_152),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_334),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_154),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_231),
.B(n_218),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_336),
.B(n_337),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_236),
.B(n_218),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_306),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_347),
.B(n_349),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_250),
.B(n_242),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_259),
.A2(n_203),
.B1(n_142),
.B2(n_155),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_275),
.A2(n_277),
.B1(n_249),
.B2(n_264),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_353),
.A2(n_274),
.B1(n_238),
.B2(n_266),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_296),
.B(n_173),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_296),
.B(n_173),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_367),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_232),
.A2(n_196),
.B1(n_197),
.B2(n_189),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_359),
.A2(n_363),
.B1(n_372),
.B2(n_245),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_259),
.A2(n_221),
.B1(n_207),
.B2(n_175),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_362),
.A2(n_301),
.B1(n_309),
.B2(n_241),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_256),
.A2(n_189),
.B1(n_202),
.B2(n_183),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_306),
.B(n_197),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_303),
.A2(n_202),
.B1(n_183),
.B2(n_201),
.Y(n_372)
);

FAx1_ASAP7_75t_SL g374 ( 
.A(n_302),
.B(n_186),
.CI(n_227),
.CON(n_374),
.SN(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g393 ( 
.A1(n_374),
.A2(n_284),
.B(n_291),
.C(n_292),
.Y(n_393)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_377),
.Y(n_434)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_375),
.Y(n_379)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_379),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_318),
.Y(n_380)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_375),
.Y(n_383)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_261),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_384),
.B(n_405),
.Y(n_465)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_330),
.Y(n_385)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_385),
.Y(n_450)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g451 ( 
.A1(n_386),
.A2(n_387),
.B1(n_400),
.B2(n_404),
.Y(n_451)
);

INVx13_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_340),
.Y(n_390)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_390),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_391),
.A2(n_365),
.B1(n_373),
.B2(n_344),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_392),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_393),
.A2(n_365),
.B(n_371),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_257),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_394),
.B(n_399),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_336),
.B(n_267),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_396),
.A2(n_412),
.B(n_368),
.Y(n_445)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_397),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_322),
.B(n_248),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_407),
.C(n_408),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_324),
.B(n_314),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_317),
.A2(n_246),
.B1(n_254),
.B2(n_279),
.Y(n_400)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_333),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_355),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_339),
.B(n_305),
.C(n_287),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_339),
.B(n_281),
.C(n_311),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_331),
.B(n_310),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_368),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_233),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_410),
.B(n_414),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_411),
.A2(n_417),
.B1(n_419),
.B2(n_372),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_265),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_355),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_420),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g414 ( 
.A(n_341),
.B(n_227),
.Y(n_414)
);

OR2x4_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_278),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_415),
.A2(n_424),
.B(n_367),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_282),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_416),
.B(n_418),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_337),
.A2(n_263),
.B1(n_235),
.B2(n_251),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_343),
.B(n_253),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_347),
.B(n_247),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_334),
.B(n_247),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_422),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_371),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_356),
.B(n_313),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_425),
.Y(n_441)
);

NOR2x1p5_ASAP7_75t_L g424 ( 
.A(n_316),
.B(n_286),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_340),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_427),
.B(n_448),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_428),
.A2(n_432),
.B1(n_435),
.B2(n_458),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_431),
.B(n_456),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_402),
.A2(n_315),
.B1(n_365),
.B2(n_359),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_412),
.A2(n_320),
.B1(n_335),
.B2(n_332),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_436),
.A2(n_395),
.B1(n_417),
.B2(n_383),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_415),
.A2(n_325),
.B(n_346),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_439),
.A2(n_440),
.B(n_452),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_422),
.A2(n_323),
.B(n_346),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_382),
.B(n_354),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_444),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_382),
.B(n_358),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_445),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_381),
.B(n_398),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_448),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_394),
.A2(n_323),
.B(n_366),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_406),
.A2(n_366),
.B(n_325),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_453),
.Y(n_503)
);

FAx1_ASAP7_75t_SL g455 ( 
.A(n_407),
.B(n_351),
.CI(n_361),
.CON(n_455),
.SN(n_455)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_455),
.B(n_408),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_412),
.A2(n_338),
.B(n_294),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_384),
.B(n_328),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_460),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_389),
.A2(n_321),
.B1(n_327),
.B2(n_370),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_401),
.B(n_321),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_389),
.A2(n_327),
.B1(n_370),
.B2(n_326),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_462),
.A2(n_389),
.B1(n_395),
.B2(n_405),
.Y(n_481)
);

AO22x1_ASAP7_75t_SL g466 ( 
.A1(n_411),
.A2(n_361),
.B1(n_345),
.B2(n_333),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_466),
.B(n_445),
.Y(n_492)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_467),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_430),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_468),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_414),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_469),
.B(n_472),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_430),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_470),
.B(n_477),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_433),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_471),
.B(n_490),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_393),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_446),
.Y(n_473)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_473),
.Y(n_518)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_460),
.Y(n_476)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_476),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_478),
.B(n_429),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_441),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_479),
.B(n_461),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_432),
.A2(n_419),
.B1(n_396),
.B2(n_424),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_480),
.A2(n_500),
.B1(n_434),
.B2(n_438),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_481),
.A2(n_447),
.B(n_459),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_452),
.A2(n_395),
.B1(n_424),
.B2(n_377),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_482),
.A2(n_489),
.B1(n_491),
.B2(n_495),
.Y(n_542)
);

INVx13_ASAP7_75t_L g484 ( 
.A(n_447),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_484),
.Y(n_513)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_486),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_429),
.B(n_381),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_455),
.C(n_456),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_428),
.A2(n_388),
.B1(n_396),
.B2(n_409),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_433),
.B(n_388),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_SL g517 ( 
.A1(n_492),
.A2(n_496),
.B(n_466),
.C(n_455),
.Y(n_517)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_463),
.Y(n_493)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_493),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_441),
.B(n_425),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g536 ( 
.A(n_494),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_436),
.A2(n_379),
.B1(n_413),
.B2(n_404),
.Y(n_495)
);

AO22x1_ASAP7_75t_L g496 ( 
.A1(n_465),
.A2(n_390),
.B1(n_397),
.B2(n_403),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_437),
.B(n_328),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_498),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_338),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_442),
.B(n_385),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_450),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_426),
.A2(n_360),
.B1(n_348),
.B2(n_342),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_426),
.A2(n_427),
.B1(n_440),
.B2(n_434),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_501),
.A2(n_462),
.B1(n_451),
.B2(n_466),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_444),
.B(n_360),
.Y(n_504)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_504),
.Y(n_540)
);

NOR4xp25_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_453),
.C(n_443),
.D(n_438),
.Y(n_506)
);

AOI21xp33_ASAP7_75t_L g556 ( 
.A1(n_506),
.A2(n_475),
.B(n_495),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_507),
.B(n_509),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_474),
.A2(n_439),
.B(n_431),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_508),
.A2(n_514),
.B(n_520),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_449),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_486),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_510),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_511),
.A2(n_531),
.B1(n_518),
.B2(n_515),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_499),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_512),
.B(n_539),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_474),
.A2(n_435),
.B(n_443),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_516),
.B(n_522),
.C(n_524),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_517),
.B(n_492),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_519),
.A2(n_503),
.B1(n_480),
.B2(n_502),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_464),
.C(n_459),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_505),
.B(n_464),
.C(n_450),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_489),
.Y(n_527)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_527),
.Y(n_554)
);

CKINVDCx14_ASAP7_75t_R g558 ( 
.A(n_528),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_483),
.A2(n_466),
.B1(n_461),
.B2(n_380),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_505),
.B(n_345),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_SL g569 ( 
.A(n_532),
.B(n_500),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_501),
.A2(n_326),
.B(n_378),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_533),
.A2(n_502),
.B(n_503),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_477),
.B(n_238),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_537),
.B(n_342),
.Y(n_576)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_538),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_490),
.B(n_392),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_488),
.B(n_243),
.C(n_285),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_541),
.B(n_543),
.C(n_493),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_488),
.B(n_364),
.C(n_170),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_544),
.A2(n_546),
.B1(n_547),
.B2(n_549),
.Y(n_579)
);

A2O1A1Ixp33_ASAP7_75t_SL g586 ( 
.A1(n_545),
.A2(n_517),
.B(n_508),
.C(n_526),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_542),
.A2(n_496),
.B1(n_502),
.B2(n_468),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_523),
.B(n_479),
.Y(n_548)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_548),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_519),
.A2(n_485),
.B1(n_476),
.B2(n_496),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_538),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_551),
.B(n_553),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_475),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g582 ( 
.A(n_552),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_536),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_504),
.Y(n_555)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_555),
.Y(n_587)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_556),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_561),
.B(n_565),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_511),
.A2(n_491),
.B1(n_472),
.B2(n_481),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_562),
.Y(n_591)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_510),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_563),
.B(n_566),
.Y(n_590)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_525),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_567),
.B(n_570),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_507),
.B(n_467),
.C(n_473),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_568),
.B(n_522),
.C(n_509),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_SL g597 ( 
.A(n_569),
.B(n_532),
.Y(n_597)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_534),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_513),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_571),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_513),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_572),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_540),
.B(n_469),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_573),
.Y(n_583)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_529),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_574),
.B(n_576),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_580),
.B(n_581),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_564),
.B(n_568),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_586),
.B(n_588),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_524),
.C(n_516),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_559),
.B(n_537),
.C(n_535),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_589),
.B(n_595),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_559),
.B(n_533),
.C(n_514),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_575),
.B(n_561),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_596),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_598),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_SL g598 ( 
.A(n_569),
.B(n_526),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_554),
.B(n_541),
.C(n_543),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_599),
.B(n_600),
.C(n_601),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_554),
.B(n_520),
.C(n_531),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_576),
.B(n_521),
.C(n_513),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_589),
.B(n_573),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_605),
.B(n_611),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_582),
.B(n_558),
.Y(n_606)
);

CKINVDCx14_ASAP7_75t_R g633 ( 
.A(n_606),
.Y(n_633)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_584),
.Y(n_608)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_608),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_580),
.B(n_547),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_609),
.B(n_614),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_583),
.A2(n_562),
.B1(n_560),
.B2(n_549),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_610),
.A2(n_517),
.B1(n_586),
.B2(n_570),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_593),
.Y(n_611)
);

NOR3xp33_ASAP7_75t_SL g612 ( 
.A(n_592),
.B(n_548),
.C(n_545),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_612),
.B(n_613),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_594),
.B(n_546),
.C(n_550),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_594),
.B(n_550),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_595),
.B(n_544),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_615),
.B(n_620),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_579),
.A2(n_572),
.B(n_571),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_616),
.A2(n_618),
.B1(n_619),
.B2(n_590),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_601),
.B(n_574),
.Y(n_617)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_617),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_599),
.A2(n_555),
.B(n_560),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_SL g619 ( 
.A1(n_585),
.A2(n_517),
.B(n_567),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_598),
.B(n_563),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_588),
.B(n_557),
.C(n_566),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_623),
.B(n_577),
.C(n_578),
.Y(n_629)
);

BUFx24_ASAP7_75t_SL g625 ( 
.A(n_622),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_625),
.B(n_629),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_623),
.Y(n_626)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_626),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_610),
.A2(n_591),
.B1(n_587),
.B2(n_602),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_632),
.A2(n_612),
.B1(n_607),
.B2(n_620),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_603),
.B(n_600),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_635),
.B(n_640),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_603),
.B(n_591),
.C(n_597),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_637),
.B(n_319),
.C(n_318),
.Y(n_652)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_638),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_639),
.A2(n_319),
.B1(n_330),
.B2(n_386),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_613),
.A2(n_586),
.B1(n_484),
.B2(n_348),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_621),
.A2(n_586),
.B(n_387),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_641),
.A2(n_614),
.B(n_609),
.Y(n_646)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_619),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_642),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_645),
.A2(n_651),
.B1(n_656),
.B2(n_648),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_646),
.B(n_648),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_636),
.A2(n_615),
.B(n_604),
.Y(n_648)
);

AOI21x1_ASAP7_75t_L g650 ( 
.A1(n_629),
.A2(n_624),
.B(n_604),
.Y(n_650)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_650),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_635),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_652),
.B(n_654),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_626),
.B(n_634),
.C(n_630),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g666 ( 
.A(n_655),
.B(n_329),
.Y(n_666)
);

CKINVDCx16_ASAP7_75t_R g656 ( 
.A(n_628),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_634),
.B(n_262),
.C(n_304),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_657),
.B(n_631),
.C(n_630),
.Y(n_659)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_658),
.Y(n_669)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_659),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_647),
.A2(n_627),
.B1(n_633),
.B2(n_644),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_660),
.A2(n_662),
.B1(n_655),
.B2(n_657),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_651),
.B(n_632),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_661),
.A2(n_663),
.B(n_646),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_643),
.A2(n_637),
.B1(n_639),
.B2(n_276),
.Y(n_662)
);

AOI321xp33_ASAP7_75t_L g663 ( 
.A1(n_650),
.A2(n_286),
.A3(n_329),
.B1(n_239),
.B2(n_294),
.C(n_234),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_666),
.B(n_649),
.C(n_654),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_645),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_667),
.Y(n_671)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_670),
.Y(n_678)
);

AOI31xp33_ASAP7_75t_L g677 ( 
.A1(n_672),
.A2(n_674),
.A3(n_659),
.B(n_667),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_664),
.B(n_653),
.C(n_652),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_675),
.A2(n_668),
.B(n_649),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_676),
.A2(n_677),
.B(n_679),
.Y(n_681)
);

A2O1A1O1Ixp25_ASAP7_75t_L g679 ( 
.A1(n_669),
.A2(n_668),
.B(n_665),
.C(n_666),
.D(n_286),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_678),
.B(n_673),
.C(n_672),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_SL g682 ( 
.A1(n_680),
.A2(n_681),
.B(n_671),
.Y(n_682)
);

AOI222xp33_ASAP7_75t_SL g683 ( 
.A1(n_682),
.A2(n_671),
.B1(n_239),
.B2(n_313),
.C1(n_240),
.C2(n_290),
.Y(n_683)
);

MAJx2_ASAP7_75t_L g684 ( 
.A(n_683),
.B(n_214),
.C(n_144),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_144),
.C(n_198),
.Y(n_685)
);

AO21x1_ASAP7_75t_L g686 ( 
.A1(n_685),
.A2(n_198),
.B(n_18),
.Y(n_686)
);


endmodule