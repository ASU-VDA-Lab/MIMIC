module real_jpeg_4981_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_286;
wire n_176;
wire n_166;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_1),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_1),
.B(n_160),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_2),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_2),
.Y(n_143)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_2),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_3),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_3),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_3),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_3),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_3),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_3),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_4),
.B(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_4),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_4),
.B(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_4),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_5),
.B(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_5),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_5),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_5),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_5),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_5),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_5),
.B(n_396),
.Y(n_395)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_7),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_7),
.Y(n_246)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_7),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_7),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_7),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_8),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_8),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_8),
.B(n_36),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_8),
.B(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_8),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_8),
.B(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_8),
.B(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_11),
.B(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_11),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_11),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_11),
.B(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_12),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_12),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_13),
.B(n_40),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_13),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_13),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_13),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_13),
.B(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_14),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_14),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_14),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_14),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_14),
.B(n_219),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_14),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_14),
.B(n_36),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_14),
.B(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_15),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_15),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_15),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g430 ( 
.A(n_15),
.Y(n_430)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

A2O1A1O1Ixp25_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_113),
.B(n_355),
.C(n_512),
.D(n_514),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_20),
.B(n_72),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_57),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_48),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_22),
.A2(n_23),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_42),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_26),
.A2(n_27),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_26),
.A2(n_27),
.B1(n_232),
.B2(n_239),
.Y(n_231)
);

NOR3xp33_ASAP7_75t_L g514 ( 
.A(n_26),
.B(n_61),
.C(n_66),
.Y(n_514)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_33),
.C(n_39),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_27),
.B(n_320),
.C(n_321),
.Y(n_319)
);

OR2x2_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_30),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_30),
.Y(n_223)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_31),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_31),
.Y(n_334)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_32),
.B(n_108),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_32),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_49),
.C(n_53),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_33),
.A2(n_34),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_34),
.B(n_154),
.C(n_159),
.Y(n_254)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_37),
.Y(n_185)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_38),
.Y(n_385)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_39),
.A2(n_42),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_39),
.B(n_341),
.C(n_344),
.Y(n_487)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_47),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_49),
.B(n_101),
.C(n_106),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_49),
.A2(n_112),
.B1(n_180),
.B2(n_191),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_49),
.B(n_181),
.C(n_187),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_49),
.A2(n_106),
.B1(n_107),
.B2(n_112),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_50),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_51),
.Y(n_372)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_52),
.Y(n_217)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_52),
.Y(n_236)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_52),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_70),
.B2(n_71),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_65),
.B2(n_69),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_60),
.A2(n_61),
.B1(n_479),
.B2(n_480),
.Y(n_478)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_86),
.C(n_90),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_66),
.A2(n_68),
.B1(n_305),
.B2(n_307),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_66),
.B(n_244),
.C(n_278),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_70),
.B(n_513),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.C(n_95),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_78),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.C(n_94),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_80),
.B1(n_94),
.B2(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_82),
.B(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_86),
.A2(n_90),
.B1(n_248),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_86),
.Y(n_481)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_90),
.A2(n_241),
.B1(n_242),
.B2(n_248),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_90),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_90),
.B(n_141),
.C(n_244),
.Y(n_294)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_92),
.Y(n_342)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_94),
.A2(n_99),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_94),
.B(n_318),
.C(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_94),
.A2(n_99),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_95),
.B(n_508),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_110),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_96),
.A2(n_97),
.B1(n_490),
.B2(n_491),
.Y(n_489)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_99),
.B(n_352),
.C(n_355),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_100),
.B(n_110),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_101),
.B(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_105),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_106),
.A2(n_107),
.B1(n_141),
.B2(n_243),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_106),
.A2(n_107),
.B1(n_278),
.B2(n_306),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_136),
.C(n_141),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_107),
.B(n_278),
.C(n_330),
.Y(n_488)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_108),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_109),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_506),
.B(n_511),
.Y(n_113)
);

AOI21x1_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_472),
.B(n_503),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_324),
.B(n_357),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_288),
.B(n_323),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_262),
.B(n_287),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_118),
.B(n_470),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_225),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_119),
.B(n_225),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_178),
.C(n_209),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_120),
.B(n_286),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_120),
.Y(n_515)
);

FAx1_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_151),
.CI(n_162),
.CON(n_120),
.SN(n_120)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_121),
.B(n_151),
.C(n_162),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_135),
.C(n_144),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_122),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_132),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_124),
.B(n_128),
.C(n_132),
.Y(n_224)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_127),
.Y(n_280)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_135),
.A2(n_144),
.B1(n_145),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_135),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_136),
.B(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_141),
.A2(n_243),
.B1(n_244),
.B2(n_247),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_141),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx8_ASAP7_75t_L g367 ( 
.A(n_143),
.Y(n_367)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_281)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_154),
.A2(n_161),
.B1(n_197),
.B2(n_198),
.Y(n_390)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_164),
.B(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_163),
.B(n_169),
.C(n_176),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_167),
.B(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_173),
.Y(n_406)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_174),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_177),
.B(n_374),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_177),
.B(n_388),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_177),
.B(n_423),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_178),
.B(n_209),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_192),
.C(n_194),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_179),
.A2(n_192),
.B1(n_193),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_179),
.Y(n_267)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B1(n_187),
.B2(n_190),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_186),
.A2(n_187),
.B1(n_296),
.B2(n_301),
.Y(n_295)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_187),
.B(n_297),
.C(n_298),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_189),
.Y(n_275)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_194),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.C(n_205),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_195),
.A2(n_196),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_200),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_460)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_224),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_212),
.C(n_224),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_220),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_218),
.C(n_220),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_214),
.A2(n_341),
.B1(n_343),
.B2(n_344),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_214),
.Y(n_344)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_217),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_226),
.B(n_228),
.C(n_261),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_249),
.B1(n_260),
.B2(n_261),
.Y(n_227)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_240),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_230),
.B(n_231),
.C(n_240),
.Y(n_309)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_233),
.Y(n_320)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_237),
.Y(n_321)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_244),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_244),
.A2(n_247),
.B1(n_278),
.B2(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_244),
.A2(n_247),
.B1(n_382),
.B2(n_383),
.Y(n_400)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_247),
.B(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_250),
.B(n_252),
.C(n_253),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_256),
.B(n_258),
.C(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_285),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_263),
.B(n_285),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.C(n_282),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_264),
.A2(n_265),
.B1(n_465),
.B2(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_268),
.B(n_282),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.C(n_281),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_269),
.B(n_452),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_271),
.B(n_281),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_276),
.C(n_278),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_272),
.A2(n_273),
.B1(n_276),
.B2(n_277),
.Y(n_379)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_278),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_278),
.A2(n_306),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_289),
.B(n_324),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_291),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_325),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_291),
.B(n_325),
.Y(n_471)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_308),
.CI(n_322),
.CON(n_291),
.SN(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_304),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_302),
.B2(n_303),
.Y(n_293)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_303),
.C(n_304),
.Y(n_347)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

INVx4_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_311),
.C(n_313),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.Y(n_313)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_319),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_326),
.B(n_328),
.C(n_345),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_345),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_336),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_329),
.B(n_337),
.C(n_338),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_341),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_348),
.B2(n_356),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_346),
.B(n_349),
.C(n_351),
.Y(n_499)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_348),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_355),
.Y(n_354)
);

OAI31xp33_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_468),
.A3(n_469),
.B(n_471),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_462),
.B(n_467),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_447),
.B(n_461),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_401),
.B(n_446),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_391),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_362),
.B(n_391),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_380),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_377),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_364),
.B(n_377),
.C(n_380),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.C(n_373),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_365),
.A2(n_366),
.B1(n_368),
.B2(n_369),
.Y(n_393)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_367),
.Y(n_432)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_373),
.B(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_381),
.B(n_456),
.C(n_457),
.Y(n_455)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_387),
.Y(n_456)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.C(n_400),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_392),
.B(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_394),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_394),
.A2(n_400),
.B1(n_438),
.B2(n_444),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_395),
.Y(n_436)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_398),
.Y(n_437)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_400),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_440),
.B(n_445),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_403),
.A2(n_426),
.B(n_439),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_411),
.B(n_425),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_407),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_422),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_422),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_417),
.B(n_421),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_417),
.Y(n_421)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_421),
.A2(n_428),
.B1(n_433),
.B2(n_434),
.Y(n_427)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_435),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_435),
.Y(n_439)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_428),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_431),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_429),
.A2(n_431),
.B(n_433),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_436),
.A2(n_437),
.B(n_438),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_441),
.B(n_442),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_449),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_451),
.B1(n_453),
.B2(n_454),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_455),
.C(n_458),
.Y(n_463)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.Y(n_454)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_463),
.B(n_464),
.Y(n_467)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_465),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_500),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_473),
.A2(n_504),
.B(n_505),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_492),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_474),
.B(n_492),
.Y(n_505)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_474),
.Y(n_518)
);

FAx1_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_483),
.CI(n_489),
.CON(n_474),
.SN(n_474)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_483),
.C(n_489),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.C(n_482),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_476),
.A2(n_477),
.B1(n_494),
.B2(n_495),
.Y(n_493)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_482),
.Y(n_494)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.C(n_488),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_484),
.A2(n_485),
.B1(n_497),
.B2(n_498),
.Y(n_496)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_488),
.Y(n_498)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_490),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_496),
.C(n_499),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_493),
.B(n_496),
.CI(n_499),
.CON(n_502),
.SN(n_502)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_494),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_501),
.B(n_502),
.Y(n_504)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_502),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_510),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_510),
.Y(n_511)
);


endmodule