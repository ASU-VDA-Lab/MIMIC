module fake_jpeg_1688_n_462 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_462);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_462;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_24),
.B1(n_33),
.B2(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_56),
.A2(n_104),
.B1(n_29),
.B2(n_52),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_60),
.B(n_61),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_16),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_62),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_67),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_15),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_82),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_72),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_35),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_22),
.B(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_78),
.B(n_90),
.Y(n_182)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_15),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_84),
.Y(n_190)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_27),
.B(n_14),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_94),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_88),
.Y(n_186)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_89),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_13),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_25),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_41),
.B(n_0),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_110),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_19),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_106),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_28),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_48),
.B(n_29),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_30),
.B(n_1),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_48),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_32),
.B(n_2),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_113),
.B(n_81),
.Y(n_188)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_28),
.B(n_53),
.Y(n_164)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_21),
.B(n_3),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_54),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_117),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_118),
.A2(n_157),
.B1(n_191),
.B2(n_186),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_119),
.A2(n_120),
.B1(n_128),
.B2(n_130),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_88),
.A2(n_43),
.B1(n_45),
.B2(n_51),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_43),
.B1(n_45),
.B2(n_51),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_21),
.B1(n_52),
.B2(n_42),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_133),
.A2(n_141),
.B1(n_166),
.B2(n_180),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_83),
.A2(n_54),
.B1(n_42),
.B2(n_37),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_143),
.B(n_155),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_56),
.A2(n_37),
.B1(n_53),
.B2(n_20),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_152),
.A2(n_167),
.B1(n_170),
.B2(n_174),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_75),
.B(n_3),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_89),
.A2(n_28),
.B1(n_26),
.B2(n_20),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_74),
.B(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_163),
.B(n_168),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_95),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_57),
.A2(n_53),
.B1(n_20),
.B2(n_26),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_91),
.A2(n_53),
.B1(n_26),
.B2(n_9),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_74),
.B(n_6),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g170 ( 
.A1(n_84),
.A2(n_53),
.B1(n_9),
.B2(n_10),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_92),
.A2(n_53),
.B1(n_9),
.B2(n_10),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_63),
.B(n_7),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_189),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_93),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_179),
.A2(n_187),
.B1(n_181),
.B2(n_165),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_58),
.A2(n_11),
.B1(n_67),
.B2(n_71),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_62),
.A2(n_11),
.B1(n_64),
.B2(n_76),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_99),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_68),
.B(n_111),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_98),
.A2(n_65),
.B1(n_108),
.B2(n_79),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_192),
.A2(n_198),
.B(n_196),
.Y(n_265)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_117),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_196),
.B(n_198),
.Y(n_268)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_197),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_110),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_199),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_201),
.B(n_202),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_140),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_129),
.B(n_97),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_203),
.B(n_205),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_80),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_204),
.B(n_208),
.Y(n_277)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_127),
.A2(n_59),
.B(n_72),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_206),
.A2(n_253),
.B(n_254),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_140),
.B(n_133),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_207),
.B(n_215),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_138),
.B(n_73),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_149),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_209),
.B(n_226),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_122),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_210),
.B(n_211),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_176),
.Y(n_211)
);

INVx4_ASAP7_75t_SL g212 ( 
.A(n_149),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_212),
.B(n_219),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_213),
.Y(n_302)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_85),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_217),
.A2(n_240),
.B1(n_241),
.B2(n_247),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_132),
.B(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_222),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_122),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_223),
.B(n_224),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_159),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_146),
.B(n_131),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_225),
.B(n_233),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_131),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_126),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_227),
.B(n_232),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_126),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_228),
.Y(n_272)
);

INVx4_ASAP7_75t_SL g229 ( 
.A(n_162),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_229),
.B(n_235),
.Y(n_297)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_230),
.Y(n_288)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_160),
.B(n_170),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_147),
.B(n_158),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_158),
.B(n_190),
.Y(n_235)
);

BUFx16f_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_244),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_160),
.B(n_161),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_243),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_171),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_246),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_159),
.A2(n_157),
.B1(n_185),
.B2(n_136),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_161),
.B(n_156),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_173),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_166),
.A2(n_134),
.B1(n_181),
.B2(n_124),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_151),
.B(n_180),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_248),
.B(n_251),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_128),
.A2(n_130),
.B1(n_119),
.B2(n_120),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_165),
.B1(n_148),
.B2(n_153),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_191),
.B(n_124),
.C(n_134),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_254),
.C(n_253),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g251 ( 
.A(n_151),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_156),
.B(n_135),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_226),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_171),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_169),
.A2(n_171),
.B(n_148),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_255),
.A2(n_257),
.B1(n_259),
.B2(n_267),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_221),
.A2(n_135),
.B1(n_153),
.B2(n_242),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_221),
.A2(n_242),
.B1(n_232),
.B2(n_192),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_265),
.A2(n_266),
.B(n_287),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_207),
.A2(n_203),
.B(n_200),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_249),
.B1(n_215),
.B2(n_238),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_252),
.B1(n_227),
.B2(n_218),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_269),
.A2(n_270),
.B1(n_276),
.B2(n_283),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_245),
.B1(n_218),
.B2(n_194),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_281),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_218),
.A2(n_206),
.B1(n_219),
.B2(n_216),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_218),
.A2(n_220),
.B1(n_193),
.B2(n_195),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_230),
.B(n_226),
.C(n_197),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_251),
.C(n_262),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_199),
.A2(n_231),
.B1(n_222),
.B2(n_234),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_296),
.B1(n_300),
.B2(n_280),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_237),
.A2(n_246),
.B1(n_244),
.B2(n_229),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_214),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_275),
.B(n_236),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_303),
.B(n_308),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_236),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_251),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_309),
.Y(n_366)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_284),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_311),
.Y(n_342)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_313),
.C(n_320),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_265),
.B(n_281),
.C(n_275),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_261),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_317),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_268),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_282),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_319),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_271),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_266),
.B(n_270),
.C(n_268),
.Y(n_320)
);

XNOR2x2_ASAP7_75t_L g321 ( 
.A(n_259),
.B(n_286),
.Y(n_321)
);

XNOR2x2_ASAP7_75t_SL g346 ( 
.A(n_321),
.B(n_258),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_315),
.Y(n_367)
);

INVx8_ASAP7_75t_L g323 ( 
.A(n_302),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_326),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_261),
.B(n_269),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_327),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_264),
.A2(n_267),
.B(n_278),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_325),
.A2(n_279),
.B(n_300),
.Y(n_357)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_286),
.B(n_301),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_262),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_329),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_272),
.B(n_295),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_333),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_297),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_331),
.B(n_337),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_289),
.Y(n_333)
);

NOR2x1_ASAP7_75t_L g334 ( 
.A(n_264),
.B(n_274),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_334),
.A2(n_313),
.B(n_320),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_336),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_285),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_272),
.B(n_295),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_278),
.B(n_279),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_338),
.B(n_292),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_316),
.A2(n_257),
.B1(n_255),
.B2(n_283),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_339),
.A2(n_310),
.B1(n_305),
.B2(n_306),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_332),
.A2(n_263),
.B1(n_258),
.B2(n_279),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_345),
.A2(n_361),
.B1(n_303),
.B2(n_337),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_321),
.Y(n_380)
);

AOI22x1_ASAP7_75t_L g350 ( 
.A1(n_332),
.A2(n_290),
.B1(n_298),
.B2(n_291),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_350),
.A2(n_359),
.B1(n_330),
.B2(n_336),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_288),
.C(n_299),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_328),
.C(n_312),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_358),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_316),
.A2(n_296),
.B1(n_293),
.B2(n_298),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_338),
.A2(n_291),
.B1(n_293),
.B2(n_299),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_360),
.B(n_304),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_333),
.A2(n_292),
.B1(n_273),
.B2(n_280),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_314),
.B(n_273),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_327),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_367),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_342),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_371),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_318),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_369),
.B(n_373),
.Y(n_393)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_342),
.Y(n_370)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_362),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_380),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_322),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_351),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_351),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_383),
.Y(n_396)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_365),
.Y(n_376)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_377),
.A2(n_385),
.B1(n_339),
.B2(n_386),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_381),
.Y(n_397)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_345),
.A2(n_317),
.B1(n_324),
.B2(n_321),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_386),
.B1(n_387),
.B2(n_349),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_356),
.A2(n_329),
.B1(n_338),
.B2(n_325),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_SL g388 ( 
.A(n_349),
.B(n_334),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_388),
.B(n_367),
.Y(n_405)
);

OAI32xp33_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_334),
.A3(n_307),
.B1(n_311),
.B2(n_326),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_358),
.Y(n_407)
);

XOR2x2_ASAP7_75t_SL g414 ( 
.A(n_391),
.B(n_378),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_370),
.B(n_353),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_395),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_353),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_402),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_399),
.A2(n_409),
.B1(n_379),
.B2(n_377),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_385),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_401),
.B(n_371),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_343),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_406),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_384),
.B(n_341),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_407),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_376),
.A2(n_341),
.B1(n_350),
.B2(n_357),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_SL g410 ( 
.A(n_403),
.B(n_372),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_410),
.A2(n_417),
.B(n_421),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_354),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_414),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_415),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_407),
.A2(n_389),
.B(n_381),
.Y(n_415)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_382),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_400),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_418),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_354),
.C(n_364),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_355),
.C(n_408),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_378),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_422),
.B(n_411),
.Y(n_432)
);

AOI322xp5_ASAP7_75t_L g424 ( 
.A1(n_392),
.A2(n_343),
.A3(n_363),
.B1(n_390),
.B2(n_364),
.C1(n_346),
.C2(n_388),
.Y(n_424)
);

BUFx24_ASAP7_75t_SL g428 ( 
.A(n_424),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_432),
.Y(n_442)
);

O2A1O1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_423),
.A2(n_409),
.B(n_392),
.C(n_408),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_SL g439 ( 
.A1(n_430),
.A2(n_396),
.B(n_404),
.C(n_417),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_397),
.C(n_361),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_434),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_397),
.C(n_352),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_422),
.B(n_380),
.Y(n_435)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_435),
.B(n_399),
.Y(n_438)
);

BUFx24_ASAP7_75t_SL g436 ( 
.A(n_428),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_438),
.Y(n_450)
);

OAI221xp5_ASAP7_75t_L g437 ( 
.A1(n_426),
.A2(n_419),
.B1(n_415),
.B2(n_413),
.C(n_396),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_437),
.A2(n_383),
.B1(n_359),
.B2(n_340),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_439),
.B(n_347),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_430),
.A2(n_416),
.B1(n_421),
.B2(n_412),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_443),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_429),
.A2(n_393),
.B(n_404),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_441),
.A2(n_360),
.B1(n_362),
.B2(n_348),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_431),
.A2(n_387),
.B1(n_393),
.B2(n_418),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_439),
.A2(n_437),
.B(n_425),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_444),
.A2(n_425),
.B1(n_346),
.B2(n_435),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_446),
.B(n_449),
.Y(n_455)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_447),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_448),
.A2(n_452),
.B(n_366),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_442),
.A2(n_350),
.B1(n_348),
.B2(n_347),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_454),
.B(n_456),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_451),
.C(n_445),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_455),
.A2(n_446),
.B(n_304),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_457),
.A2(n_459),
.B(n_323),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_323),
.C(n_456),
.Y(n_459)
);

BUFx24_ASAP7_75t_SL g461 ( 
.A(n_460),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_458),
.Y(n_462)
);


endmodule