module fake_jpeg_12730_n_601 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_601);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_601;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_5),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_84),
.Y(n_124)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_8),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_69),
.B(n_81),
.Y(n_130)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_78),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_19),
.B(n_8),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_82),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_36),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_89),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_90),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_92),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_36),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_94),
.B(n_97),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_17),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_98),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_99),
.B(n_101),
.Y(n_176)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_36),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx5_ASAP7_75t_SL g180 ( 
.A(n_105),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_41),
.B(n_8),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_12),
.Y(n_182)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx5_ASAP7_75t_SL g193 ( 
.A(n_109),
.Y(n_193)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_110),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_24),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_113),
.Y(n_187)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_114),
.Y(n_171)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_115),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_49),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_116),
.B(n_47),
.Y(n_169)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_42),
.Y(n_119)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_47),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_125),
.B(n_0),
.Y(n_254)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_60),
.B(n_45),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_136),
.B(n_166),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_85),
.A2(n_43),
.B1(n_41),
.B2(n_54),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_137),
.A2(n_145),
.B1(n_33),
.B2(n_31),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_44),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_138),
.B(n_168),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_78),
.A2(n_43),
.B1(n_111),
.B2(n_95),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_60),
.A2(n_47),
.B1(n_55),
.B2(n_43),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_149),
.A2(n_113),
.B1(n_33),
.B2(n_31),
.Y(n_203)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_150),
.Y(n_209)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_161),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_100),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_109),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_191),
.Y(n_201)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_77),
.B(n_54),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_182),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_66),
.Y(n_189)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_114),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_102),
.B(n_48),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_51),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_74),
.B(n_48),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_91),
.Y(n_206)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_198),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_199),
.A2(n_215),
.B1(n_226),
.B2(n_23),
.Y(n_320)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_200),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_203),
.A2(n_217),
.B1(n_221),
.B2(n_236),
.Y(n_308)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_204),
.Y(n_305)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

BUFx2_ASAP7_75t_SL g313 ( 
.A(n_205),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_206),
.B(n_212),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_73),
.C(n_75),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_207),
.B(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_208),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_125),
.A2(n_104),
.B1(n_79),
.B2(n_93),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_210),
.A2(n_229),
.B(n_189),
.Y(n_300)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_211),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_46),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_92),
.B1(n_90),
.B2(n_45),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_138),
.A2(n_108),
.B1(n_29),
.B2(n_34),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_171),
.A2(n_91),
.B1(n_74),
.B2(n_46),
.Y(n_218)
);

OAI22x1_ASAP7_75t_L g288 ( 
.A1(n_218),
.A2(n_230),
.B1(n_235),
.B2(n_189),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_130),
.B(n_51),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_124),
.B(n_164),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_220),
.B(n_223),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_149),
.A2(n_39),
.B1(n_29),
.B2(n_34),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_225),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_52),
.B1(n_35),
.B2(n_56),
.Y(n_226)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g270 ( 
.A(n_227),
.Y(n_270)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_123),
.Y(n_228)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_228),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_196),
.A2(n_83),
.B1(n_58),
.B2(n_52),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_171),
.A2(n_35),
.B1(n_56),
.B2(n_39),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_133),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_231),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_148),
.B(n_105),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_251),
.Y(n_268)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_184),
.A2(n_56),
.B1(n_39),
.B2(n_37),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_173),
.A2(n_56),
.B1(n_39),
.B2(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_131),
.Y(n_237)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_237),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_131),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_238),
.Y(n_275)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_141),
.Y(n_239)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_126),
.B(n_11),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_240),
.B(n_250),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_127),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_242),
.A2(n_195),
.B1(n_174),
.B2(n_186),
.Y(n_280)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_173),
.A2(n_37),
.B1(n_35),
.B2(n_34),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_244),
.A2(n_258),
.B1(n_23),
.B2(n_165),
.Y(n_306)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_162),
.Y(n_245)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

BUFx4f_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_249),
.B(n_252),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_29),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_140),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_254),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_167),
.B(n_9),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_255),
.B(n_264),
.Y(n_317)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

INVx4_ASAP7_75t_SL g299 ( 
.A(n_256),
.Y(n_299)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_178),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_257),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_122),
.A2(n_29),
.B1(n_23),
.B2(n_2),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_129),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_259),
.B(n_195),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_128),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_260),
.Y(n_273)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_135),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_156),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_187),
.B(n_23),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_187),
.B(n_7),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_132),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_207),
.B(n_150),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_266),
.B(n_269),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_151),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_219),
.B(n_201),
.C(n_197),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_278),
.B(n_304),
.C(n_239),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_280),
.A2(n_295),
.B1(n_306),
.B2(n_320),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_288),
.A2(n_152),
.B1(n_263),
.B2(n_213),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_289),
.B(n_292),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_199),
.A2(n_157),
.B1(n_151),
.B2(n_170),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_241),
.B(n_135),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_297),
.B(n_315),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_300),
.A2(n_209),
.B(n_213),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_232),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_312),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_160),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_157),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_311),
.Y(n_338)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_225),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_309),
.Y(n_324)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_216),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_243),
.B(n_245),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_232),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_205),
.B(n_214),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_247),
.B(n_165),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_183),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_319),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_242),
.A2(n_147),
.B1(n_122),
.B2(n_159),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_322),
.A2(n_224),
.B1(n_227),
.B2(n_202),
.Y(n_333)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_285),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_328),
.B(n_345),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_308),
.A2(n_210),
.B1(n_229),
.B2(n_159),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_329),
.A2(n_346),
.B1(n_351),
.B2(n_358),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_279),
.B(n_211),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_330),
.B(n_361),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_333),
.A2(n_348),
.B1(n_362),
.B2(n_272),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g402 ( 
.A1(n_334),
.A2(n_271),
.B1(n_274),
.B2(n_287),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_335),
.A2(n_268),
.B(n_319),
.Y(n_369)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

INVx13_ASAP7_75t_L g339 ( 
.A(n_299),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_339),
.Y(n_400)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_270),
.Y(n_340)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_340),
.Y(n_389)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

BUFx12_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_342),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_344),
.B(n_301),
.Y(n_384)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_308),
.A2(n_251),
.B1(n_233),
.B2(n_253),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_360),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_295),
.A2(n_202),
.B1(n_216),
.B2(n_147),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_349),
.A2(n_352),
.B1(n_281),
.B2(n_267),
.Y(n_385)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_354),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_266),
.A2(n_183),
.B1(n_186),
.B2(n_209),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_293),
.B(n_0),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_356),
.Y(n_377)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_300),
.A2(n_263),
.B(n_148),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_357),
.A2(n_268),
.B(n_319),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_269),
.A2(n_248),
.B1(n_256),
.B2(n_257),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_293),
.B(n_121),
.C(n_261),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_304),
.Y(n_374)
);

BUFx12f_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_291),
.B(n_262),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_280),
.A2(n_262),
.B1(n_246),
.B2(n_146),
.Y(n_362)
);

NAND3xp33_ASAP7_75t_SL g363 ( 
.A(n_289),
.B(n_121),
.C(n_246),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_363),
.B(n_367),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_317),
.A2(n_146),
.B1(n_144),
.B2(n_143),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_364),
.A2(n_294),
.B1(n_283),
.B2(n_275),
.Y(n_395)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_365),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_277),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_284),
.Y(n_381)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_342),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_368),
.B(n_360),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_369),
.A2(n_394),
.B(n_324),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_323),
.A2(n_282),
.B1(n_288),
.B2(n_316),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_370),
.A2(n_382),
.B1(n_397),
.B2(n_404),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_372),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_384),
.C(n_387),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_380),
.A2(n_395),
.B(n_335),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_323),
.A2(n_322),
.B1(n_276),
.B2(n_314),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_385),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_278),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_301),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_390),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_337),
.B(n_301),
.Y(n_390)
);

NOR2x1_ASAP7_75t_L g391 ( 
.A(n_332),
.B(n_268),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_391),
.B(n_358),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_329),
.A2(n_267),
.B1(n_314),
.B2(n_281),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_344),
.B(n_305),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_398),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_367),
.A2(n_291),
.B1(n_283),
.B2(n_296),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_286),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_325),
.B(n_271),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_403),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_340),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_345),
.B(n_274),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_338),
.A2(n_287),
.B1(n_298),
.B2(n_290),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_326),
.B(n_298),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_406),
.B(n_378),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_370),
.A2(n_351),
.B1(n_338),
.B2(n_357),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_408),
.A2(n_427),
.B1(n_376),
.B2(n_377),
.Y(n_446)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_371),
.Y(n_409)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_409),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_410),
.A2(n_440),
.B(n_435),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_379),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_415),
.Y(n_445)
);

OA22x2_ASAP7_75t_L g412 ( 
.A1(n_376),
.A2(n_333),
.B1(n_362),
.B2(n_348),
.Y(n_412)
);

OA22x2_ASAP7_75t_L g449 ( 
.A1(n_412),
.A2(n_405),
.B1(n_393),
.B2(n_389),
.Y(n_449)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_413),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_417),
.Y(n_444)
);

NOR3xp33_ASAP7_75t_SL g467 ( 
.A(n_419),
.B(n_387),
.C(n_365),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_420),
.A2(n_392),
.B1(n_349),
.B2(n_339),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_403),
.B(n_354),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_421),
.B(n_426),
.Y(n_452)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_375),
.Y(n_422)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_422),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_401),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_429),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_383),
.B(n_360),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_350),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_382),
.A2(n_353),
.B1(n_352),
.B2(n_327),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_378),
.B(n_343),
.Y(n_428)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_428),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_388),
.B(n_343),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_404),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_438),
.Y(n_471)
);

INVx13_ASAP7_75t_L g431 ( 
.A(n_400),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_431),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_375),
.B(n_356),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_432),
.B(n_442),
.Y(n_456)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_373),
.Y(n_434)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_435),
.A2(n_436),
.B(n_440),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_369),
.B(n_341),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_368),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_402),
.A2(n_324),
.B1(n_331),
.B2(n_366),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_386),
.B1(n_342),
.B2(n_321),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_380),
.A2(n_395),
.B(n_391),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_399),
.B(n_321),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_384),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_414),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_446),
.A2(n_466),
.B1(n_423),
.B2(n_430),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_416),
.B(n_396),
.C(n_374),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_448),
.B(n_455),
.C(n_414),
.Y(n_492)
);

A2O1A1Ixp33_ASAP7_75t_SL g494 ( 
.A1(n_449),
.A2(n_412),
.B(n_420),
.C(n_434),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_450),
.A2(n_462),
.B(n_472),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_398),
.C(n_390),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_417),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_465),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_377),
.Y(n_459)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_459),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_413),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_460),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_424),
.B(n_389),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_461),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_410),
.A2(n_373),
.B(n_405),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_463),
.A2(n_469),
.B1(n_439),
.B2(n_441),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_386),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_464),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_432),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_467),
.A2(n_415),
.B1(n_419),
.B2(n_408),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_423),
.A2(n_290),
.B1(n_146),
.B2(n_144),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_436),
.A2(n_144),
.B(n_143),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_436),
.A2(n_143),
.B(n_135),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_473),
.B(n_411),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_476),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_493),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_458),
.Y(n_479)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_479),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_448),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_492),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_459),
.Y(n_482)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_482),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_483),
.A2(n_487),
.B1(n_495),
.B2(n_501),
.Y(n_523)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_460),
.B(n_407),
.CI(n_418),
.CON(n_484),
.SN(n_484)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_484),
.B(n_467),
.CI(n_437),
.CON(n_514),
.SN(n_514)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_461),
.Y(n_486)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_486),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_446),
.A2(n_436),
.B1(n_420),
.B2(n_429),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_488),
.A2(n_496),
.B1(n_451),
.B2(n_465),
.Y(n_508)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_449),
.Y(n_489)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_489),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_443),
.B(n_418),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_494),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_444),
.A2(n_433),
.B1(n_422),
.B2(n_412),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_447),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_474),
.A2(n_437),
.B1(n_427),
.B2(n_439),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_497),
.A2(n_503),
.B1(n_502),
.B2(n_462),
.Y(n_507)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_498),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_458),
.B(n_407),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_500),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_442),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_452),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_445),
.B(n_425),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_474),
.A2(n_437),
.B1(n_426),
.B2(n_421),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_457),
.C(n_444),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_506),
.B(n_513),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_507),
.A2(n_508),
.B1(n_515),
.B2(n_521),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_510),
.B(n_484),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_492),
.B(n_450),
.C(n_456),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_514),
.B(n_527),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_497),
.A2(n_503),
.B1(n_477),
.B2(n_489),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_478),
.B(n_456),
.C(n_468),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_519),
.B(n_526),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_491),
.A2(n_453),
.B1(n_454),
.B2(n_466),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_481),
.A2(n_454),
.B1(n_453),
.B2(n_449),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_522),
.A2(n_464),
.B1(n_494),
.B2(n_451),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_490),
.A2(n_468),
.B(n_471),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_524),
.A2(n_470),
.B(n_431),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_525),
.B(n_475),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_493),
.B(n_490),
.C(n_499),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_483),
.A2(n_445),
.B1(n_471),
.B2(n_463),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_512),
.A2(n_485),
.B1(n_496),
.B2(n_488),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_529),
.B(n_537),
.Y(n_561)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_531),
.Y(n_555)
);

AND3x1_ASAP7_75t_L g532 ( 
.A(n_511),
.B(n_494),
.C(n_487),
.Y(n_532)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_532),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_522),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_533),
.B(n_507),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_472),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_534),
.B(n_538),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_536),
.A2(n_524),
.B1(n_516),
.B2(n_517),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_523),
.A2(n_494),
.B1(n_467),
.B2(n_449),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_449),
.C(n_473),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_543),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_513),
.B(n_484),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_540),
.B(n_510),
.Y(n_553)
);

INVx13_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_541),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_518),
.A2(n_420),
.B(n_469),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_514),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_509),
.B(n_475),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_526),
.C(n_525),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_546),
.A2(n_537),
.B(n_521),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_547),
.B(n_548),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_SL g548 ( 
.A(n_530),
.B(n_519),
.C(n_514),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_504),
.C(n_509),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_551),
.B(n_556),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_552),
.A2(n_562),
.B1(n_529),
.B2(n_532),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_553),
.A2(n_557),
.B(n_535),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_554),
.A2(n_535),
.B1(n_536),
.B2(n_546),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_528),
.B(n_520),
.Y(n_556)
);

AND2x2_ASAP7_75t_SL g558 ( 
.A(n_538),
.B(n_515),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_558),
.Y(n_575)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_563),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_564),
.B(n_566),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_565),
.B(n_557),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_561),
.A2(n_540),
.B1(n_539),
.B2(n_470),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_543),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_568),
.B(n_570),
.Y(n_581)
);

A2O1A1Ixp33_ASAP7_75t_SL g569 ( 
.A1(n_559),
.A2(n_541),
.B(n_542),
.C(n_412),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_569),
.A2(n_562),
.B(n_555),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_558),
.A2(n_561),
.B1(n_547),
.B2(n_560),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_551),
.B(n_544),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_573),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_550),
.B(n_534),
.C(n_412),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_552),
.B(n_431),
.C(n_1),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_574),
.B(n_0),
.C(n_1),
.Y(n_582)
);

AOI21xp33_ASAP7_75t_L g578 ( 
.A1(n_575),
.A2(n_548),
.B(n_549),
.Y(n_578)
);

AO21x1_ASAP7_75t_L g590 ( 
.A1(n_578),
.A2(n_579),
.B(n_569),
.Y(n_590)
);

AOI21x1_ASAP7_75t_SL g589 ( 
.A1(n_580),
.A2(n_583),
.B(n_569),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_582),
.B(n_574),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_567),
.A2(n_16),
.B(n_2),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_584),
.B(n_571),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_585),
.B(n_586),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_573),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_SL g591 ( 
.A(n_587),
.B(n_579),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_564),
.C(n_569),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_588),
.B(n_590),
.C(n_10),
.Y(n_594)
);

OAI321xp33_ASAP7_75t_L g593 ( 
.A1(n_589),
.A2(n_580),
.A3(n_590),
.B1(n_581),
.B2(n_5),
.C(n_7),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_591),
.B(n_594),
.C(n_589),
.Y(n_595)
);

AOI322xp5_ASAP7_75t_L g596 ( 
.A1(n_593),
.A2(n_7),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_16),
.C2(n_11),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_595),
.B(n_596),
.C(n_592),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_597),
.A2(n_3),
.B1(n_4),
.B2(n_12),
.Y(n_598)
);

AO21x1_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_3),
.B(n_4),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_599),
.B(n_13),
.C(n_1),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_600),
.A2(n_13),
.B(n_224),
.Y(n_601)
);


endmodule