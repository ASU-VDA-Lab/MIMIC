module fake_jpeg_27929_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_6),
.B(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_7),
.A2(n_10),
.B1(n_14),
.B2(n_11),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_15),
.A2(n_23),
.B1(n_14),
.B2(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_23),
.Y(n_32)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_8),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_21),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_6),
.B1(n_17),
.B2(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_28),
.B1(n_18),
.B2(n_19),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_16),
.A2(n_6),
.B1(n_18),
.B2(n_20),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_31),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_39),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_21),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_22),
.C(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

XNOR2x1_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_25),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_45),
.C(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.C(n_48),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_37),
.C(n_41),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_44),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_44),
.B(n_42),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_49),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_50),
.Y(n_53)
);


endmodule