module fake_ariane_1652_n_1118 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1118);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1118;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_1016;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_958;
wire n_945;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_754;
wire n_336;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_1099;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_458;
wire n_361;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_658;
wire n_617;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_847;
wire n_772;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_1026;
wire n_951;
wire n_213;
wire n_938;
wire n_895;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

BUFx10_ASAP7_75t_L g206 ( 
.A(n_36),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_6),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_15),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_92),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_94),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_35),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_54),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_43),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_107),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_48),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_95),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_154),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_72),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_41),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_139),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_176),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_10),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_108),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_183),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_205),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_113),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_85),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_195),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_142),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_138),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_70),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_96),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_105),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_181),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_141),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_134),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_14),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_76),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_199),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_103),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_186),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_67),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_48),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_39),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_39),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_41),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_140),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_50),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_11),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_152),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_13),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_184),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_124),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_148),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_51),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_131),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_243),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_221),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_233),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_221),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_256),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_271),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_211),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_211),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_206),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_206),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_206),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_230),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_209),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_208),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_222),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_239),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_208),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_223),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_213),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_235),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_213),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_217),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_236),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_217),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_267),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_212),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_267),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_265),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_240),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_212),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_268),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_241),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_244),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_268),
.Y(n_326)
);

OAI22x1_ASAP7_75t_L g327 ( 
.A1(n_287),
.A2(n_259),
.B1(n_227),
.B2(n_219),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_307),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_247),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_323),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_302),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_260),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_289),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_326),
.A2(n_270),
.B1(n_262),
.B2(n_214),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_237),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_300),
.B(n_249),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_286),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_290),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_290),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_277),
.A2(n_288),
.B1(n_291),
.B2(n_294),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_295),
.B(n_237),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

AND2x6_ASAP7_75t_L g361 ( 
.A(n_298),
.B(n_252),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_279),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_280),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_281),
.B(n_269),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_282),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_283),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_284),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_299),
.Y(n_368)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_295),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_288),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_277),
.A2(n_234),
.B1(n_269),
.B2(n_261),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_291),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_306),
.A2(n_252),
.B1(n_253),
.B2(n_273),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_296),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_297),
.A2(n_263),
.B1(n_274),
.B2(n_266),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_312),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_278),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_312),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_210),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_382),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_349),
.B(n_313),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_349),
.B(n_315),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_334),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_329),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_328),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_350),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_349),
.B(n_315),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_350),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_317),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_350),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_351),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_354),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

BUFx8_ASAP7_75t_L g416 ( 
.A(n_333),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_357),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_349),
.B(n_317),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_372),
.A2(n_373),
.B1(n_381),
.B2(n_374),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_372),
.A2(n_319),
.B1(n_248),
.B2(n_246),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_337),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_373),
.A2(n_319),
.B1(n_250),
.B2(n_242),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_335),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_345),
.B(n_218),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_357),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_336),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_SL g437 ( 
.A(n_380),
.B(n_377),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_376),
.A2(n_310),
.B1(n_320),
.B2(n_303),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_376),
.A2(n_275),
.B1(n_264),
.B2(n_257),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_347),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_345),
.B(n_1),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_343),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_340),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_367),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_347),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_347),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_332),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_374),
.A2(n_228),
.B1(n_254),
.B2(n_232),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_367),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_352),
.B(n_1),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_332),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_364),
.B(n_220),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_342),
.A2(n_225),
.B1(n_226),
.B2(n_231),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_332),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_407),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_419),
.B(n_377),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_407),
.Y(n_463)
);

BUFx6f_ASAP7_75t_SL g464 ( 
.A(n_443),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_377),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

NOR3xp33_ASAP7_75t_L g469 ( 
.A(n_459),
.B(n_377),
.C(n_381),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_403),
.B(n_378),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_L g471 ( 
.A(n_437),
.B(n_380),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_403),
.B(n_378),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_380),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_380),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_414),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_402),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_380),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

BUFx6f_ASAP7_75t_SL g479 ( 
.A(n_416),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_420),
.B(n_369),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_387),
.B(n_383),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_394),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_415),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_369),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_L g485 ( 
.A(n_424),
.B(n_352),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_423),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_426),
.B(n_369),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_388),
.B(n_383),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_422),
.B(n_369),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_423),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

BUFx5_ASAP7_75t_L g494 ( 
.A(n_397),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_430),
.B(n_369),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_400),
.B(n_369),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_454),
.B(n_384),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_431),
.B(n_339),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_446),
.B(n_339),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_428),
.B(n_368),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_L g504 ( 
.A(n_418),
.B(n_368),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_439),
.B(n_375),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_396),
.B(n_355),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_342),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_396),
.B(n_356),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_402),
.B(n_379),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_385),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_414),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_385),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_440),
.B(n_379),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_444),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_389),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_L g516 ( 
.A(n_453),
.B(n_370),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_389),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_391),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_386),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_398),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_391),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_416),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_370),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_416),
.B(n_327),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_456),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_392),
.B(n_355),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_457),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_457),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_392),
.B(n_359),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_L g531 ( 
.A(n_417),
.B(n_346),
.C(n_365),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_417),
.B(n_359),
.Y(n_532)
);

BUFx6f_ASAP7_75t_SL g533 ( 
.A(n_456),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_417),
.B(n_341),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_414),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_413),
.B(n_331),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_413),
.B(n_367),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_427),
.B(n_365),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_406),
.B(n_365),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_406),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_408),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_397),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_408),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_470),
.B(n_472),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_513),
.A2(n_429),
.B1(n_434),
.B2(n_427),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_485),
.A2(n_434),
.B1(n_435),
.B2(n_429),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_360),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_507),
.A2(n_327),
.B1(n_353),
.B2(n_348),
.Y(n_550)
);

NAND2x1p5_ASAP7_75t_L g551 ( 
.A(n_532),
.B(n_509),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_472),
.A2(n_469),
.B1(n_464),
.B2(n_481),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_469),
.A2(n_464),
.B1(n_490),
.B2(n_481),
.Y(n_553)
);

NAND2x1p5_ASAP7_75t_L g554 ( 
.A(n_467),
.B(n_360),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_479),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_468),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_478),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_482),
.Y(n_558)
);

CKINVDCx16_ASAP7_75t_R g559 ( 
.A(n_476),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_486),
.B(n_493),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_540),
.Y(n_562)
);

AO22x2_ASAP7_75t_L g563 ( 
.A1(n_462),
.A2(n_348),
.B1(n_358),
.B2(n_353),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_526),
.A2(n_358),
.B1(n_366),
.B2(n_363),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_533),
.A2(n_363),
.B1(n_366),
.B2(n_435),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_512),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_520),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

NAND2x1p5_ASAP7_75t_L g569 ( 
.A(n_475),
.B(n_441),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_475),
.B(n_441),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_520),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_473),
.A2(n_399),
.B1(n_404),
.B2(n_401),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_518),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_521),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_490),
.B(n_367),
.Y(n_575)
);

NAND2x1p5_ASAP7_75t_L g576 ( 
.A(n_475),
.B(n_447),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_541),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_533),
.A2(n_448),
.B1(n_449),
.B2(n_447),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_522),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_519),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_519),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_515),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_475),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_527),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_529),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_474),
.A2(n_449),
.B1(n_450),
.B2(n_448),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_522),
.B(n_450),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_506),
.Y(n_591)
);

AO22x2_ASAP7_75t_L g592 ( 
.A1(n_477),
.A2(n_498),
.B1(n_524),
.B2(n_465),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_499),
.B(n_367),
.Y(n_593)
);

NAND2x1p5_ASAP7_75t_L g594 ( 
.A(n_488),
.B(n_455),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_461),
.Y(n_595)
);

AO22x2_ASAP7_75t_L g596 ( 
.A1(n_524),
.A2(n_455),
.B1(n_411),
.B2(n_412),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_463),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_508),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_501),
.A2(n_508),
.B1(n_505),
.B2(n_466),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_534),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_543),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_543),
.A2(n_399),
.B1(n_401),
.B2(n_404),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_483),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_531),
.A2(n_405),
.B1(n_411),
.B2(n_409),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_505),
.B(n_405),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_487),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_505),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_524),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_492),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_545),
.B(n_503),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g611 ( 
.A1(n_572),
.A2(n_570),
.B(n_569),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_548),
.B(n_537),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_598),
.B(n_537),
.Y(n_613)
);

O2A1O1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_593),
.A2(n_504),
.B(n_531),
.C(n_523),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_601),
.A2(n_471),
.B(n_480),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_553),
.A2(n_491),
.B1(n_535),
.B2(n_484),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_583),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_562),
.A2(n_516),
.B(n_539),
.C(n_535),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_567),
.B(n_494),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_579),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_606),
.Y(n_622)
);

O2A1O1Ixp33_ASAP7_75t_L g623 ( 
.A1(n_561),
.A2(n_495),
.B(n_489),
.C(n_496),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_571),
.B(n_564),
.Y(n_624)
);

NAND2x1p5_ASAP7_75t_L g625 ( 
.A(n_584),
.B(n_488),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_575),
.A2(n_538),
.B(n_511),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_581),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_599),
.B(n_494),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_552),
.B(n_494),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_602),
.A2(n_511),
.B(n_488),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_591),
.B(n_494),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_582),
.B(n_460),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_584),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_560),
.A2(n_511),
.B1(n_525),
.B2(n_488),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_557),
.B(n_558),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_586),
.B(n_494),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_590),
.B(n_511),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_585),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_559),
.B(n_497),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_579),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_564),
.A2(n_550),
.B1(n_565),
.B2(n_578),
.Y(n_641)
);

BUFx4f_ASAP7_75t_L g642 ( 
.A(n_551),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_604),
.A2(n_410),
.B(n_409),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_589),
.A2(n_412),
.B(n_410),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_561),
.A2(n_536),
.B(n_525),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_566),
.B(n_332),
.C(n_390),
.Y(n_646)
);

CKINVDCx11_ASAP7_75t_R g647 ( 
.A(n_580),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_568),
.B(n_494),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_590),
.B(n_525),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_573),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_565),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_605),
.B(n_525),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_574),
.A2(n_502),
.B(n_500),
.Y(n_653)
);

O2A1O1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_577),
.A2(n_514),
.B(n_421),
.C(n_433),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_549),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_588),
.A2(n_536),
.B(n_542),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g657 ( 
.A1(n_546),
.A2(n_421),
.B(n_390),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_550),
.B(n_542),
.Y(n_658)
);

AOI21x1_ASAP7_75t_L g659 ( 
.A1(n_563),
.A2(n_536),
.B(n_542),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_554),
.B(n_605),
.Y(n_660)
);

OAI21xp33_ASAP7_75t_L g661 ( 
.A1(n_563),
.A2(n_421),
.B(n_390),
.Y(n_661)
);

OAI21xp33_ASAP7_75t_L g662 ( 
.A1(n_547),
.A2(n_436),
.B(n_433),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_607),
.A2(n_361),
.B1(n_542),
.B2(n_544),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_600),
.A2(n_433),
.B(n_436),
.C(n_438),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_576),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_609),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_592),
.B(n_544),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_594),
.A2(n_438),
.B(n_436),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_637),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_616),
.Y(n_670)
);

CKINVDCx8_ASAP7_75t_R g671 ( 
.A(n_655),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_610),
.A2(n_592),
.B1(n_588),
.B2(n_596),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_624),
.B(n_627),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_666),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_613),
.B(n_555),
.Y(n_675)
);

BUFx4f_ASAP7_75t_SL g676 ( 
.A(n_621),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_639),
.B(n_595),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_650),
.B(n_612),
.Y(n_678)
);

BUFx8_ASAP7_75t_L g679 ( 
.A(n_640),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_635),
.B(n_596),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_629),
.A2(n_578),
.B1(n_608),
.B2(n_536),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_618),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_647),
.B(n_361),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_622),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_660),
.B(n_597),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_637),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_638),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_SL g688 ( 
.A(n_619),
.B(n_641),
.C(n_614),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_642),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_655),
.B(n_642),
.Y(n_690)
);

AND3x1_ASAP7_75t_SL g691 ( 
.A(n_620),
.B(n_2),
.C(n_3),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_655),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_651),
.B(n_652),
.Y(n_693)
);

AND2x2_ASAP7_75t_SL g694 ( 
.A(n_667),
.B(n_544),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_633),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_649),
.B(n_603),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_648),
.A2(n_609),
.B1(n_587),
.B2(n_544),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_659),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_632),
.B(n_658),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_628),
.B(n_438),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_633),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_SL g702 ( 
.A1(n_663),
.A2(n_625),
.B1(n_633),
.B2(n_631),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_653),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_665),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_665),
.B(n_361),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_636),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_656),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_625),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_644),
.B(n_361),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_668),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_611),
.B(n_442),
.Y(n_711)
);

INVx8_ASAP7_75t_L g712 ( 
.A(n_661),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_619),
.B(n_361),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_617),
.A2(n_361),
.B1(n_451),
.B2(n_442),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_654),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_654),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_634),
.Y(n_717)
);

NAND2x1p5_ASAP7_75t_L g718 ( 
.A(n_656),
.B(n_442),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_645),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_643),
.B(n_451),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_646),
.A2(n_361),
.B1(n_347),
.B2(n_255),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_662),
.A2(n_452),
.B1(n_451),
.B2(n_255),
.Y(n_722)
);

AND3x1_ASAP7_75t_SL g723 ( 
.A(n_614),
.B(n_3),
.C(n_4),
.Y(n_723)
);

CKINVDCx8_ASAP7_75t_R g724 ( 
.A(n_664),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_657),
.B(n_4),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_630),
.A2(n_452),
.B1(n_255),
.B2(n_7),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_645),
.B(n_452),
.Y(n_727)
);

INVx3_ASAP7_75t_SL g728 ( 
.A(n_701),
.Y(n_728)
);

INVx6_ASAP7_75t_SL g729 ( 
.A(n_711),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_674),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_686),
.B(n_630),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_670),
.Y(n_732)
);

NAND2x1p5_ASAP7_75t_L g733 ( 
.A(n_686),
.B(n_626),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_682),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_674),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_706),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_717),
.A2(n_623),
.B(n_615),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_706),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_684),
.Y(n_739)
);

NAND2x1_ASAP7_75t_L g740 ( 
.A(n_711),
.B(n_626),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_689),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_SL g742 ( 
.A1(n_688),
.A2(n_664),
.B(n_623),
.C(n_615),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_675),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_699),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_673),
.B(n_5),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_687),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_679),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_678),
.B(n_8),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_689),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_687),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_698),
.Y(n_751)
);

INVx4_ASAP7_75t_L g752 ( 
.A(n_676),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_685),
.Y(n_753)
);

O2A1O1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_688),
.A2(n_675),
.B(n_725),
.C(n_716),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_717),
.A2(n_8),
.B(n_9),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_698),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_689),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_703),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_727),
.A2(n_9),
.B(n_10),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_704),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_677),
.B(n_11),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_683),
.B(n_12),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_696),
.Y(n_763)
);

AO21x2_ASAP7_75t_L g764 ( 
.A1(n_672),
.A2(n_255),
.B(n_53),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_693),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_704),
.B(n_12),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_669),
.B(n_13),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_689),
.Y(n_768)
);

INVx8_ASAP7_75t_L g769 ( 
.A(n_692),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_669),
.B(n_14),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_719),
.Y(n_771)
);

NAND2x1_ASAP7_75t_L g772 ( 
.A(n_715),
.B(n_255),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_676),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_669),
.B(n_15),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_726),
.A2(n_712),
.B(n_714),
.C(n_700),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_679),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_724),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_702),
.B(n_255),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_692),
.B(n_16),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_719),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_680),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_694),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_669),
.B(n_17),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_690),
.B(n_18),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_694),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_695),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_712),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_695),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_713),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_719),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_720),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_712),
.A2(n_22),
.B(n_23),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_719),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_671),
.B(n_24),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_710),
.A2(n_25),
.B(n_26),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_745),
.B(n_708),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_744),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_753),
.B(n_700),
.Y(n_798)
);

O2A1O1Ixp5_ASAP7_75t_L g799 ( 
.A1(n_737),
.A2(n_710),
.B(n_697),
.C(n_709),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_758),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_728),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_782),
.B(n_785),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_730),
.B(n_707),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_748),
.B(n_681),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_744),
.B(n_707),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_730),
.B(n_735),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_752),
.B(n_722),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_769),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_767),
.B(n_718),
.Y(n_809)
);

CKINVDCx14_ASAP7_75t_R g810 ( 
.A(n_747),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_774),
.B(n_718),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_SL g812 ( 
.A1(n_787),
.A2(n_705),
.B(n_723),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_SL g813 ( 
.A1(n_747),
.A2(n_723),
.B1(n_691),
.B2(n_721),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_732),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_728),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_734),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_787),
.A2(n_691),
.B(n_721),
.C(n_28),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_754),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_752),
.B(n_27),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_763),
.B(n_781),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_755),
.B(n_255),
.C(n_29),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_760),
.B(n_29),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_758),
.Y(n_823)
);

CKINVDCx12_ASAP7_75t_R g824 ( 
.A(n_794),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_792),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_739),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_736),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_765),
.B(n_30),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_788),
.B(n_31),
.Y(n_829)
);

BUFx12f_ASAP7_75t_L g830 ( 
.A(n_776),
.Y(n_830)
);

AOI21x1_ASAP7_75t_SL g831 ( 
.A1(n_766),
.A2(n_32),
.B(n_33),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_771),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_761),
.B(n_33),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_784),
.B(n_34),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_762),
.B(n_34),
.Y(n_835)
);

INVx5_ASAP7_75t_L g836 ( 
.A(n_731),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_771),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_736),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_769),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_SL g840 ( 
.A1(n_775),
.A2(n_35),
.B(n_36),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_746),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_775),
.A2(n_743),
.B1(n_777),
.B2(n_791),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_731),
.B(n_52),
.Y(n_843)
);

OR2x6_ASAP7_75t_SL g844 ( 
.A(n_776),
.B(n_37),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_769),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_733),
.Y(n_846)
);

OAI21x1_ASAP7_75t_SL g847 ( 
.A1(n_789),
.A2(n_37),
.B(n_38),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_770),
.B(n_38),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_779),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_SL g850 ( 
.A1(n_759),
.A2(n_40),
.B(n_42),
.C(n_44),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_784),
.B(n_44),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_742),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_795),
.A2(n_778),
.B(n_770),
.C(n_783),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_742),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_786),
.B(n_49),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_738),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_738),
.B(n_49),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_778),
.A2(n_55),
.B(n_56),
.C(n_57),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_842),
.A2(n_786),
.B1(n_733),
.B2(n_729),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_805),
.B(n_780),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_808),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_804),
.A2(n_764),
.B1(n_750),
.B2(n_746),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_814),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_813),
.A2(n_764),
.B1(n_729),
.B2(n_756),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_802),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_SL g866 ( 
.A1(n_834),
.A2(n_773),
.B1(n_741),
.B2(n_757),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_830),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_L g868 ( 
.A1(n_817),
.A2(n_729),
.B1(n_741),
.B2(n_768),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_821),
.A2(n_751),
.B1(n_756),
.B2(n_780),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_816),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_817),
.A2(n_851),
.B1(n_818),
.B2(n_854),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_847),
.A2(n_757),
.B1(n_741),
.B2(n_749),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_806),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_826),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_797),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_848),
.A2(n_757),
.B1(n_741),
.B2(n_749),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_849),
.A2(n_757),
.B1(n_749),
.B2(n_768),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_818),
.A2(n_768),
.B1(n_749),
.B2(n_740),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_796),
.B(n_790),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_798),
.B(n_790),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_802),
.A2(n_751),
.B1(n_793),
.B2(n_768),
.Y(n_881)
);

OAI22x1_ASAP7_75t_L g882 ( 
.A1(n_822),
.A2(n_793),
.B1(n_772),
.B2(n_60),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_806),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_820),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_836),
.Y(n_885)
);

OAI22xp33_ASAP7_75t_L g886 ( 
.A1(n_833),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_852),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_800),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_809),
.B(n_204),
.Y(n_889)
);

INVx5_ASAP7_75t_SL g890 ( 
.A(n_808),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_808),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_800),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_801),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_843),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_825),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_841),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_839),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_835),
.A2(n_201),
.B1(n_73),
.B2(n_74),
.Y(n_898)
);

OAI21xp33_ASAP7_75t_L g899 ( 
.A1(n_840),
.A2(n_71),
.B(n_75),
.Y(n_899)
);

BUFx4f_ASAP7_75t_SL g900 ( 
.A(n_815),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_823),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_827),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_902)
);

OAI21xp33_ASAP7_75t_L g903 ( 
.A1(n_852),
.A2(n_80),
.B(n_81),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_810),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_836),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_854),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_SL g907 ( 
.A1(n_836),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_907)
);

BUFx8_ASAP7_75t_L g908 ( 
.A(n_855),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_823),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_871),
.A2(n_853),
.B(n_819),
.C(n_850),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_863),
.Y(n_911)
);

NOR2x1_ASAP7_75t_SL g912 ( 
.A(n_894),
.B(n_836),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_875),
.B(n_832),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_860),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_865),
.B(n_885),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_880),
.B(n_832),
.Y(n_916)
);

OA21x2_ASAP7_75t_L g917 ( 
.A1(n_901),
.A2(n_799),
.B(n_856),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_865),
.B(n_845),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_880),
.B(n_846),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_885),
.B(n_803),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_860),
.B(n_888),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_871),
.A2(n_858),
.B(n_843),
.C(n_807),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_896),
.Y(n_923)
);

NAND4xp25_ASAP7_75t_SL g924 ( 
.A(n_864),
.B(n_844),
.C(n_812),
.D(n_829),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_892),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_899),
.A2(n_868),
.B1(n_903),
.B2(n_906),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_887),
.A2(n_799),
.B(n_803),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_887),
.A2(n_828),
.B(n_857),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_879),
.B(n_837),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_893),
.B(n_837),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_861),
.B(n_811),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_894),
.B(n_838),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_868),
.A2(n_906),
.B1(n_878),
.B2(n_895),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_870),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_884),
.B(n_831),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_874),
.B(n_824),
.Y(n_936)
);

AOI221xp5_ASAP7_75t_L g937 ( 
.A1(n_878),
.A2(n_831),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_859),
.A2(n_89),
.B(n_97),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_866),
.B(n_98),
.Y(n_939)
);

AOI221xp5_ASAP7_75t_L g940 ( 
.A1(n_886),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.C(n_102),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_862),
.A2(n_859),
.B(n_877),
.C(n_898),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_905),
.B(n_104),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_909),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_873),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_914),
.B(n_905),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_930),
.B(n_883),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_918),
.B(n_897),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_929),
.B(n_897),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_915),
.B(n_897),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_915),
.B(n_891),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_914),
.B(n_869),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_925),
.B(n_891),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_932),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_925),
.B(n_891),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_924),
.A2(n_882),
.B1(n_908),
.B2(n_907),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_932),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_943),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_917),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_931),
.B(n_904),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_943),
.B(n_876),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_921),
.B(n_881),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_911),
.B(n_908),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_917),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_935),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_934),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_916),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_927),
.B(n_889),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_932),
.B(n_890),
.Y(n_968)
);

AOI211xp5_ASAP7_75t_L g969 ( 
.A1(n_960),
.A2(n_910),
.B(n_922),
.C(n_926),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_958),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_958),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_964),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_965),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_967),
.A2(n_910),
.B(n_922),
.Y(n_974)
);

AOI31xp33_ASAP7_75t_L g975 ( 
.A1(n_955),
.A2(n_933),
.A3(n_938),
.B(n_867),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_967),
.A2(n_941),
.B(n_927),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_965),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_967),
.A2(n_941),
.B(n_939),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_957),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_964),
.B(n_919),
.Y(n_980)
);

BUFx8_ASAP7_75t_L g981 ( 
.A(n_959),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_967),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_958),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_967),
.A2(n_939),
.B(n_928),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_957),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_982),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_969),
.B(n_966),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_974),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_982),
.B(n_953),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_982),
.B(n_953),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_976),
.B(n_956),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_970),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_970),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_972),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_979),
.B(n_956),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_977),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_977),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_979),
.B(n_949),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_988),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_988),
.Y(n_1000)
);

NAND4xp25_ASAP7_75t_L g1001 ( 
.A(n_989),
.B(n_978),
.C(n_984),
.D(n_955),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_992),
.Y(n_1002)
);

OA21x2_ASAP7_75t_L g1003 ( 
.A1(n_987),
.A2(n_971),
.B(n_983),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_998),
.B(n_949),
.Y(n_1004)
);

AO21x2_ASAP7_75t_L g1005 ( 
.A1(n_991),
.A2(n_983),
.B(n_971),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_986),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_989),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_1007),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_1004),
.B(n_990),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_999),
.Y(n_1010)
);

O2A1O1Ixp5_ASAP7_75t_SL g1011 ( 
.A1(n_1006),
.A2(n_986),
.B(n_994),
.C(n_997),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_999),
.B(n_980),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1000),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1000),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_1010),
.B(n_981),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_1012),
.B(n_1007),
.Y(n_1016)
);

AND3x1_ASAP7_75t_L g1017 ( 
.A(n_1008),
.B(n_991),
.C(n_986),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1008),
.B(n_1005),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_1009),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_1009),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_1013),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_1014),
.B(n_981),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1011),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_1010),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_1024),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1021),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_1017),
.A2(n_1003),
.B1(n_1001),
.B2(n_1005),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_1019),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1020),
.A2(n_990),
.B(n_975),
.Y(n_1029)
);

OAI322xp33_ASAP7_75t_L g1030 ( 
.A1(n_1023),
.A2(n_1006),
.A3(n_1002),
.B1(n_963),
.B2(n_997),
.C1(n_996),
.C2(n_1003),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_1018),
.A2(n_1021),
.B(n_1015),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1016),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1028),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1025),
.B(n_1022),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1026),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_1032),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_L g1037 ( 
.A(n_1029),
.B(n_1027),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1031),
.B(n_998),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1030),
.B(n_995),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_SL g1040 ( 
.A(n_1034),
.B(n_1036),
.C(n_1033),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1037),
.A2(n_1003),
.B(n_996),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1035),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_1038),
.B(n_1002),
.C(n_940),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_SL g1044 ( 
.A(n_1039),
.B(n_981),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1041),
.B(n_995),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1042),
.B(n_963),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_1040),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1043),
.Y(n_1048)
);

OAI221xp5_ASAP7_75t_L g1049 ( 
.A1(n_1044),
.A2(n_993),
.B1(n_992),
.B2(n_937),
.C(n_962),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1042),
.B(n_959),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_1050),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1048),
.B(n_985),
.Y(n_1052)
);

OAI21xp33_ASAP7_75t_SL g1053 ( 
.A1(n_1047),
.A2(n_962),
.B(n_985),
.Y(n_1053)
);

AOI211xp5_ASAP7_75t_L g1054 ( 
.A1(n_1045),
.A2(n_1046),
.B(n_1049),
.C(n_993),
.Y(n_1054)
);

AOI322xp5_ASAP7_75t_L g1055 ( 
.A1(n_1048),
.A2(n_951),
.A3(n_960),
.B1(n_961),
.B2(n_872),
.C1(n_945),
.C2(n_973),
.Y(n_1055)
);

OAI221xp5_ASAP7_75t_L g1056 ( 
.A1(n_1045),
.A2(n_951),
.B1(n_936),
.B2(n_945),
.C(n_961),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1051),
.B(n_966),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1053),
.B(n_900),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1052),
.Y(n_1059)
);

NOR2x1_ASAP7_75t_L g1060 ( 
.A(n_1056),
.B(n_968),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1057),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_1059),
.B(n_1054),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1058),
.B(n_1055),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1060),
.B(n_947),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_1058),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1057),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1057),
.B(n_952),
.Y(n_1067)
);

NOR2x1_ASAP7_75t_L g1068 ( 
.A(n_1059),
.B(n_968),
.Y(n_1068)
);

OAI322xp33_ASAP7_75t_L g1069 ( 
.A1(n_1063),
.A2(n_913),
.A3(n_952),
.B1(n_954),
.B2(n_942),
.C1(n_947),
.C2(n_948),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1061),
.Y(n_1070)
);

NAND4xp75_ASAP7_75t_L g1071 ( 
.A(n_1066),
.B(n_954),
.C(n_950),
.D(n_948),
.Y(n_1071)
);

OAI211xp5_ASAP7_75t_SL g1072 ( 
.A1(n_1062),
.A2(n_902),
.B(n_890),
.C(n_912),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1068),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1064),
.B(n_950),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1067),
.A2(n_890),
.B1(n_946),
.B2(n_944),
.Y(n_1075)
);

OAI211xp5_ASAP7_75t_SL g1076 ( 
.A1(n_1065),
.A2(n_106),
.B(n_109),
.C(n_110),
.Y(n_1076)
);

AOI31xp33_ASAP7_75t_L g1077 ( 
.A1(n_1061),
.A2(n_946),
.A3(n_920),
.B(n_114),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_1073),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1070),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_1077),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_1074),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_1071),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1075),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1069),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1076),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1072),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1073),
.Y(n_1087)
);

OA22x2_ASAP7_75t_L g1088 ( 
.A1(n_1073),
.A2(n_920),
.B1(n_923),
.B2(n_115),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1073),
.Y(n_1089)
);

INVxp33_ASAP7_75t_SL g1090 ( 
.A(n_1070),
.Y(n_1090)
);

OAI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1078),
.A2(n_111),
.B1(n_112),
.B2(n_116),
.Y(n_1091)
);

OAI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_1082),
.A2(n_1084),
.B1(n_1089),
.B2(n_1087),
.C(n_1081),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_1082),
.B(n_1080),
.Y(n_1093)
);

AOI221x1_ASAP7_75t_L g1094 ( 
.A1(n_1079),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.C(n_120),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_SL g1095 ( 
.A(n_1086),
.B(n_1085),
.C(n_1083),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_1090),
.A2(n_121),
.B(n_123),
.Y(n_1096)
);

AOI322xp5_ASAP7_75t_L g1097 ( 
.A1(n_1088),
.A2(n_125),
.A3(n_126),
.B1(n_127),
.B2(n_128),
.C1(n_129),
.C2(n_130),
.Y(n_1097)
);

OA22x2_ASAP7_75t_L g1098 ( 
.A1(n_1078),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_1092),
.A2(n_136),
.B1(n_137),
.B2(n_143),
.C(n_144),
.Y(n_1099)
);

AND4x1_ASAP7_75t_L g1100 ( 
.A(n_1094),
.B(n_145),
.C(n_146),
.D(n_147),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_1093),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_1095),
.B(n_149),
.C(n_150),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1091),
.A2(n_151),
.B(n_153),
.C(n_155),
.Y(n_1103)
);

NOR3xp33_ASAP7_75t_L g1104 ( 
.A(n_1098),
.B(n_1096),
.C(n_1097),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1101),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1104),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_1102),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1106),
.A2(n_1103),
.B(n_1100),
.Y(n_1108)
);

OR3x1_ASAP7_75t_L g1109 ( 
.A(n_1108),
.B(n_1107),
.C(n_1099),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_L g1110 ( 
.A(n_1109),
.B(n_1105),
.C(n_165),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_1109),
.B(n_162),
.Y(n_1111)
);

OAI222xp33_ASAP7_75t_L g1112 ( 
.A1(n_1111),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.C1(n_170),
.C2(n_171),
.Y(n_1112)
);

OAI322xp33_ASAP7_75t_L g1113 ( 
.A1(n_1110),
.A2(n_173),
.A3(n_174),
.B1(n_175),
.B2(n_177),
.C1(n_178),
.C2(n_180),
.Y(n_1113)
);

XNOR2xp5_ASAP7_75t_L g1114 ( 
.A(n_1111),
.B(n_187),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_1114),
.B(n_188),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1112),
.A2(n_189),
.B(n_190),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1116),
.A2(n_1115),
.B(n_1113),
.C(n_193),
.Y(n_1117)
);

AOI211xp5_ASAP7_75t_L g1118 ( 
.A1(n_1117),
.A2(n_191),
.B(n_192),
.C(n_194),
.Y(n_1118)
);


endmodule