module fake_aes_7655_n_923 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_923);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_923;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_922;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_921;
wire n_543;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_195;
wire n_165;
wire n_285;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_916;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_29), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_71), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_3), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_10), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_22), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_62), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_14), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_57), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_107), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_53), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_26), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_29), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_30), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_15), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_65), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_28), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_0), .Y(n_132) );
INVx2_ASAP7_75t_SL g133 ( .A(n_38), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_58), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_1), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_32), .Y(n_137) );
BUFx10_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_54), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_100), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_11), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_81), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_16), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_38), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_52), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_99), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_34), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_12), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g149 ( .A(n_27), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_25), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_72), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_45), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_33), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_88), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_25), .Y(n_155) );
INVx4_ASAP7_75t_R g156 ( .A(n_68), .Y(n_156) );
INVx5_ASAP7_75t_L g157 ( .A(n_139), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_139), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_119), .B(n_0), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_118), .B(n_133), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_139), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_113), .B(n_1), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_118), .B(n_133), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_119), .B(n_2), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_119), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_136), .Y(n_168) );
BUFx12f_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g172 ( .A(n_120), .B(n_44), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_115), .Y(n_173) );
INVx5_ASAP7_75t_L g174 ( .A(n_138), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_135), .Y(n_175) );
BUFx12f_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_135), .B(n_2), .Y(n_177) );
INVx5_ASAP7_75t_L g178 ( .A(n_118), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_133), .B(n_3), .Y(n_179) );
NOR2xp33_ASAP7_75t_SL g180 ( .A(n_124), .B(n_46), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_170), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_163), .A2(n_113), .B1(n_149), .B2(n_128), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_164), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_163), .A2(n_128), .B1(n_149), .B2(n_114), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_174), .B(n_122), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_164), .Y(n_186) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_160), .B(n_115), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_164), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_174), .B(n_117), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_163), .A2(n_141), .B1(n_132), .B2(n_121), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_163), .A2(n_155), .B1(n_129), .B2(n_153), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_174), .B(n_169), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_169), .A2(n_127), .B1(n_143), .B2(n_144), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g194 ( .A1(n_169), .A2(n_155), .B1(n_129), .B2(n_125), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_169), .A2(n_137), .B1(n_126), .B2(n_153), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_174), .B(n_122), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_169), .A2(n_131), .B1(n_147), .B2(n_148), .Y(n_197) );
AO22x2_ASAP7_75t_L g198 ( .A1(n_177), .A2(n_131), .B1(n_147), .B2(n_150), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_174), .B(n_148), .Y(n_199) );
AO22x2_ASAP7_75t_L g200 ( .A1(n_177), .A2(n_150), .B1(n_154), .B2(n_140), .Y(n_200) );
OAI22xp33_ASAP7_75t_SL g201 ( .A1(n_180), .A2(n_116), .B1(n_123), .B2(n_130), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_176), .A2(n_116), .B1(n_154), .B2(n_123), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_176), .A2(n_145), .B1(n_134), .B2(n_140), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_160), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_160), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_174), .A2(n_145), .B1(n_134), .B2(n_130), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_176), .A2(n_152), .B1(n_151), .B2(n_146), .Y(n_207) );
OAI22xp33_ASAP7_75t_SL g208 ( .A1(n_180), .A2(n_142), .B1(n_5), .B2(n_6), .Y(n_208) );
OAI22xp33_ASAP7_75t_SL g209 ( .A1(n_180), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_176), .A2(n_160), .B1(n_165), .B2(n_177), .Y(n_210) );
OAI22xp5_ASAP7_75t_SL g211 ( .A1(n_176), .A2(n_179), .B1(n_161), .B2(n_160), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g212 ( .A1(n_173), .A2(n_174), .B1(n_179), .B2(n_161), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_170), .Y(n_213) );
INVxp67_ASAP7_75t_SL g214 ( .A(n_173), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_160), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_174), .B(n_4), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_173), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_160), .Y(n_219) );
OAI22xp33_ASAP7_75t_SL g220 ( .A1(n_172), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_174), .B(n_12), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_167), .B(n_13), .Y(n_222) );
OAI22xp33_ASAP7_75t_SL g223 ( .A1(n_172), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_223) );
AO22x2_ASAP7_75t_L g224 ( .A1(n_177), .A2(n_156), .B1(n_17), .B2(n_18), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_174), .B(n_16), .Y(n_225) );
OA22x2_ASAP7_75t_L g226 ( .A1(n_165), .A2(n_177), .B1(n_168), .B2(n_158), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_165), .A2(n_156), .B1(n_18), .B2(n_19), .Y(n_227) );
AO22x2_ASAP7_75t_L g228 ( .A1(n_177), .A2(n_17), .B1(n_19), .B2(n_20), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_174), .B(n_20), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_214), .Y(n_230) );
XOR2xp5_ASAP7_75t_L g231 ( .A(n_194), .B(n_165), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_205), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_214), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_205), .Y(n_234) );
XOR2x2_ASAP7_75t_L g235 ( .A(n_184), .B(n_161), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_205), .Y(n_236) );
XNOR2xp5_ASAP7_75t_L g237 ( .A(n_191), .B(n_167), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_226), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_204), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_192), .Y(n_240) );
INVxp67_ASAP7_75t_L g241 ( .A(n_183), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_186), .B(n_174), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_188), .B(n_167), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_198), .B(n_174), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_226), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_215), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_192), .B(n_167), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_198), .B(n_167), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_193), .B(n_167), .Y(n_249) );
AND2x2_ASAP7_75t_SL g250 ( .A(n_187), .B(n_177), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_189), .B(n_167), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_216), .Y(n_252) );
INVxp67_ASAP7_75t_SL g253 ( .A(n_210), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_219), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_181), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_181), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_207), .B(n_179), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_195), .B(n_177), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_198), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_185), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_185), .Y(n_261) );
NOR2xp33_ASAP7_75t_SL g262 ( .A(n_182), .B(n_172), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_200), .Y(n_263) );
NAND2xp33_ASAP7_75t_SL g264 ( .A(n_211), .B(n_165), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_200), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_200), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_196), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_187), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_190), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_213), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_212), .B(n_178), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_199), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_224), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_224), .B(n_165), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_182), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_202), .B(n_165), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_228), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
XOR2xp5_ASAP7_75t_L g282 ( .A(n_191), .B(n_165), .Y(n_282) );
INVxp33_ASAP7_75t_L g283 ( .A(n_197), .Y(n_283) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_222), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_228), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_217), .Y(n_286) );
INVxp67_ASAP7_75t_L g287 ( .A(n_203), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_221), .Y(n_288) );
INVx4_ASAP7_75t_SL g289 ( .A(n_225), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_206), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_209), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_220), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_223), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_212), .B(n_178), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_232), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_250), .B(n_227), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_232), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_234), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_234), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_250), .B(n_166), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_250), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_241), .B(n_166), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_240), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_283), .B(n_201), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_236), .Y(n_306) );
INVx3_ASAP7_75t_SL g307 ( .A(n_268), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_257), .B(n_208), .Y(n_308) );
INVx4_ASAP7_75t_L g309 ( .A(n_244), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_236), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_230), .B(n_178), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_230), .B(n_178), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_282), .B(n_178), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_255), .Y(n_315) );
BUFx4_ASAP7_75t_SL g316 ( .A(n_273), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_282), .B(n_268), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_233), .B(n_178), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_246), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_275), .B(n_166), .Y(n_320) );
AND2x2_ASAP7_75t_SL g321 ( .A(n_275), .B(n_166), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_233), .B(n_178), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_253), .B(n_166), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_237), .B(n_166), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_255), .Y(n_325) );
OR2x4_ASAP7_75t_L g326 ( .A(n_258), .B(n_158), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_238), .B(n_178), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_238), .B(n_178), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_237), .B(n_166), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_256), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_245), .B(n_290), .Y(n_332) );
INVxp67_ASAP7_75t_L g333 ( .A(n_244), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_287), .B(n_178), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_240), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_246), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_279), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_291), .B(n_178), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_291), .B(n_166), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_292), .B(n_175), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_252), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_256), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_245), .B(n_178), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_252), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_290), .B(n_178), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_292), .B(n_175), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_293), .B(n_175), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_298), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_298), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_298), .Y(n_352) );
NOR2xp33_ASAP7_75t_SL g353 ( .A(n_309), .B(n_263), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_308), .B(n_276), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_319), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_319), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_298), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_319), .Y(n_358) );
NAND2xp33_ASAP7_75t_L g359 ( .A(n_298), .B(n_265), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_309), .B(n_265), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_298), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_337), .B(n_293), .Y(n_362) );
OR2x6_ASAP7_75t_L g363 ( .A(n_309), .B(n_266), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_298), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_337), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_298), .Y(n_366) );
AND2x6_ASAP7_75t_L g367 ( .A(n_302), .B(n_266), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_298), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_315), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_301), .B(n_273), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_308), .B(n_269), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_301), .B(n_274), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_298), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_337), .B(n_274), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_301), .B(n_259), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_298), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_309), .B(n_231), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_309), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_298), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_337), .B(n_254), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_310), .Y(n_382) );
BUFx8_ASAP7_75t_L g383 ( .A(n_369), .Y(n_383) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_351), .Y(n_384) );
BUFx6f_ASAP7_75t_SL g385 ( .A(n_360), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_354), .A2(n_308), .B1(n_296), .B2(n_264), .Y(n_386) );
BUFx12f_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_369), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_351), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_351), .Y(n_390) );
NAND2x1p5_ASAP7_75t_L g391 ( .A(n_351), .B(n_310), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
BUFx2_ASAP7_75t_R g393 ( .A(n_378), .Y(n_393) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
INVx5_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_349), .B(n_309), .Y(n_396) );
BUFx4_ASAP7_75t_SL g397 ( .A(n_379), .Y(n_397) );
BUFx12f_ASAP7_75t_L g398 ( .A(n_379), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_379), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_354), .B(n_342), .Y(n_400) );
BUFx6f_ASAP7_75t_SL g401 ( .A(n_360), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_357), .Y(n_402) );
BUFx5_ASAP7_75t_L g403 ( .A(n_367), .Y(n_403) );
BUFx8_ASAP7_75t_L g404 ( .A(n_367), .Y(n_404) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_351), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_353), .B(n_280), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_349), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_357), .Y(n_408) );
INVx2_ASAP7_75t_SL g409 ( .A(n_352), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_352), .Y(n_410) );
BUFx4f_ASAP7_75t_SL g411 ( .A(n_370), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_372), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_395), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_386), .A2(n_372), .B1(n_262), .B2(n_296), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_396), .B(n_370), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_407), .Y(n_416) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_411), .A2(n_353), .B1(n_378), .B2(n_309), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_400), .B(n_349), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_407), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_391), .Y(n_420) );
OAI22xp5_ASAP7_75t_SL g421 ( .A1(n_412), .A2(n_378), .B1(n_231), .B2(n_360), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_411), .A2(n_326), .B1(n_363), .B2(n_360), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_391), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_386), .A2(n_296), .B1(n_302), .B2(n_314), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_383), .A2(n_296), .B1(n_302), .B2(n_314), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_400), .B(n_355), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_397), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_387), .A2(n_326), .B1(n_363), .B2(n_360), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_383), .A2(n_302), .B1(n_314), .B2(n_305), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_383), .A2(n_302), .B1(n_398), .B2(n_387), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_397), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_390), .A2(n_359), .B(n_370), .Y(n_432) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_406), .A2(n_305), .B(n_281), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_395), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g437 ( .A1(n_393), .A2(n_281), .B(n_280), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_383), .A2(n_314), .B1(n_305), .B2(n_321), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_385), .A2(n_326), .B1(n_360), .B2(n_363), .Y(n_439) );
CKINVDCx6p67_ASAP7_75t_R g440 ( .A(n_387), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_396), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_396), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_402), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_402), .Y(n_444) );
CKINVDCx11_ASAP7_75t_R g445 ( .A(n_398), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_384), .Y(n_446) );
CKINVDCx11_ASAP7_75t_R g447 ( .A(n_398), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_395), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_383), .A2(n_314), .B1(n_321), .B2(n_330), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_395), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_404), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_385), .A2(n_367), .B1(n_317), .B2(n_360), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_385), .A2(n_321), .B1(n_330), .B2(n_324), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_384), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_388), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_388), .B(n_370), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_385), .A2(n_321), .B1(n_330), .B2(n_324), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_404), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_439), .A2(n_385), .B1(n_401), .B2(n_393), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_421), .A2(n_401), .B1(n_404), .B2(n_367), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_450), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_456), .B(n_366), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_416), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_416), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_443), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_419), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_419), .Y(n_467) );
INVx4_ASAP7_75t_L g468 ( .A(n_458), .Y(n_468) );
INVx4_ASAP7_75t_L g469 ( .A(n_458), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_421), .A2(n_401), .B1(n_404), .B2(n_367), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_456), .B(n_366), .Y(n_471) );
CKINVDCx11_ASAP7_75t_R g472 ( .A(n_445), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_439), .A2(n_417), .B1(n_452), .B2(n_449), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_441), .B(n_371), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_413), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_420), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_414), .A2(n_401), .B1(n_404), .B2(n_367), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_446), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_427), .B(n_403), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_428), .A2(n_401), .B1(n_367), .B2(n_321), .Y(n_480) );
BUFx12f_ASAP7_75t_L g481 ( .A(n_447), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_438), .A2(n_367), .B1(n_321), .B2(n_388), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_441), .B(n_371), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_420), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_423), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_452), .A2(n_363), .B1(n_326), .B2(n_399), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_434), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_446), .Y(n_489) );
OAI222xp33_ASAP7_75t_L g490 ( .A1(n_451), .A2(n_363), .B1(n_399), .B2(n_218), .C1(n_285), .C2(n_406), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_422), .A2(n_363), .B1(n_326), .B2(n_399), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_434), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_453), .A2(n_367), .B1(n_330), .B2(n_324), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_457), .A2(n_367), .B1(n_324), .B2(n_363), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_458), .A2(n_367), .B1(n_317), .B2(n_403), .Y(n_495) );
NOR2x1_ASAP7_75t_R g496 ( .A(n_431), .B(n_403), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_442), .B(n_371), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_443), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g499 ( .A1(n_427), .A2(n_218), .B1(n_235), .B2(n_285), .C1(n_317), .C2(n_373), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_435), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_424), .A2(n_317), .B1(n_403), .B2(n_373), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_442), .B(n_373), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g503 ( .A1(n_451), .A2(n_403), .B1(n_395), .B2(n_317), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_437), .A2(n_403), .B1(n_376), .B2(n_348), .Y(n_504) );
BUFx4f_ASAP7_75t_SL g505 ( .A(n_440), .Y(n_505) );
OAI21xp5_ASAP7_75t_SL g506 ( .A1(n_430), .A2(n_333), .B(n_316), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_437), .A2(n_403), .B1(n_376), .B2(n_348), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_435), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_418), .A2(n_326), .B1(n_381), .B2(n_358), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_429), .A2(n_403), .B1(n_376), .B2(n_348), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_440), .A2(n_358), .B1(n_355), .B2(n_381), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_446), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_425), .A2(n_358), .B1(n_355), .B2(n_365), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_450), .A2(n_403), .B1(n_395), .B2(n_408), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_433), .A2(n_348), .B(n_362), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_415), .B(n_408), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_455), .A2(n_403), .B1(n_348), .B2(n_341), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_455), .A2(n_403), .B1(n_347), .B2(n_341), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_454), .Y(n_519) );
BUFx4f_ASAP7_75t_SL g520 ( .A(n_450), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g521 ( .A1(n_450), .A2(n_418), .B1(n_426), .B2(n_444), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_413), .A2(n_403), .B1(n_395), .B2(n_362), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_426), .A2(n_365), .B1(n_356), .B2(n_333), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_413), .B(n_395), .Y(n_524) );
OAI21xp5_ASAP7_75t_SL g525 ( .A1(n_413), .A2(n_333), .B(n_316), .Y(n_525) );
INVx5_ASAP7_75t_SL g526 ( .A(n_413), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_454), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_413), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_436), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_454), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_444), .A2(n_356), .B1(n_375), .B2(n_342), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_415), .A2(n_375), .B1(n_345), .B2(n_342), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_433), .A2(n_347), .B1(n_341), .B2(n_235), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_484), .Y(n_535) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_459), .A2(n_448), .B1(n_436), .B2(n_410), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_473), .A2(n_347), .B1(n_341), .B2(n_448), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_486), .A2(n_347), .B1(n_448), .B2(n_436), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g539 ( .A1(n_499), .A2(n_249), .B1(n_168), .B2(n_158), .C(n_171), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_511), .A2(n_175), .B(n_432), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_460), .A2(n_448), .B1(n_436), .B2(n_432), .Y(n_541) );
OAI221xp5_ASAP7_75t_SL g542 ( .A1(n_499), .A2(n_171), .B1(n_168), .B2(n_340), .C(n_332), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_459), .A2(n_448), .B1(n_436), .B2(n_340), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_491), .A2(n_448), .B1(n_436), .B2(n_340), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_482), .A2(n_340), .B1(n_338), .B2(n_310), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_463), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_480), .A2(n_310), .B1(n_338), .B2(n_342), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_470), .A2(n_310), .B1(n_338), .B2(n_345), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_506), .A2(n_525), .B1(n_468), .B2(n_469), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_509), .A2(n_310), .B1(n_338), .B2(n_345), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_506), .A2(n_409), .B1(n_390), .B2(n_389), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_509), .A2(n_310), .B1(n_338), .B2(n_345), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_494), .A2(n_310), .B1(n_338), .B2(n_320), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_465), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_525), .B(n_162), .C(n_171), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_477), .A2(n_310), .B1(n_338), .B2(n_320), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_463), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_493), .A2(n_310), .B1(n_338), .B2(n_320), .Y(n_558) );
INVx4_ASAP7_75t_L g559 ( .A(n_468), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_501), .A2(n_310), .B1(n_338), .B2(n_320), .Y(n_560) );
AOI22xp33_ASAP7_75t_SL g561 ( .A1(n_468), .A2(n_410), .B1(n_389), .B2(n_390), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_510), .A2(n_310), .B1(n_338), .B2(n_301), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_469), .A2(n_338), .B1(n_323), .B2(n_335), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_469), .A2(n_323), .B1(n_335), .B2(n_389), .Y(n_564) );
AOI222xp33_ASAP7_75t_L g565 ( .A1(n_505), .A2(n_332), .B1(n_277), .B2(n_159), .C1(n_339), .C2(n_323), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_503), .A2(n_409), .B1(n_389), .B2(n_364), .Y(n_566) );
OAI22xp5_ASAP7_75t_SL g567 ( .A1(n_481), .A2(n_316), .B1(n_394), .B2(n_384), .Y(n_567) );
AOI222xp33_ASAP7_75t_L g568 ( .A1(n_481), .A2(n_332), .B1(n_159), .B2(n_339), .C1(n_323), .C2(n_175), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_464), .B(n_159), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_495), .A2(n_335), .B1(n_159), .B2(n_336), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_513), .A2(n_159), .B1(n_336), .B2(n_359), .Y(n_571) );
NAND3xp33_ASAP7_75t_SL g572 ( .A(n_514), .B(n_248), .C(n_21), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_520), .A2(n_405), .B1(n_394), .B2(n_384), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_464), .B(n_159), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_504), .A2(n_368), .B1(n_374), .B2(n_361), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_507), .A2(n_159), .B1(n_336), .B2(n_327), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_523), .A2(n_334), .B1(n_339), .B2(n_336), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_521), .A2(n_336), .B1(n_327), .B2(n_304), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_467), .Y(n_579) );
OAI22xp33_ASAP7_75t_SL g580 ( .A1(n_484), .A2(n_368), .B1(n_374), .B2(n_350), .Y(n_580) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_519), .A2(n_346), .B(n_350), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_533), .A2(n_350), .B1(n_361), .B2(n_382), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_521), .A2(n_327), .B1(n_304), .B2(n_334), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_515), .A2(n_327), .B1(n_304), .B2(n_334), .Y(n_584) );
OA21x2_ASAP7_75t_L g585 ( .A1(n_519), .A2(n_346), .B(n_361), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_485), .A2(n_382), .B1(n_394), .B2(n_384), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_467), .B(n_384), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_516), .B(n_384), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_515), .A2(n_327), .B1(n_304), .B2(n_405), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_462), .B(n_384), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_485), .A2(n_327), .B1(n_304), .B2(n_405), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_522), .A2(n_382), .B1(n_394), .B2(n_405), .Y(n_592) );
AOI211xp5_ASAP7_75t_L g593 ( .A1(n_490), .A2(n_307), .B(n_294), .C(n_248), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_517), .A2(n_327), .B1(n_304), .B2(n_405), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g595 ( .A1(n_518), .A2(n_382), .B1(n_394), .B2(n_405), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_532), .A2(n_327), .B1(n_304), .B2(n_405), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_474), .A2(n_304), .B1(n_405), .B2(n_394), .Y(n_597) );
OAI221xp5_ASAP7_75t_L g598 ( .A1(n_461), .A2(n_272), .B1(n_267), .B2(n_260), .C(n_261), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_531), .A2(n_339), .B1(n_311), .B2(n_306), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_476), .A2(n_382), .B1(n_394), .B2(n_392), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_483), .A2(n_339), .B1(n_392), .B2(n_289), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_497), .A2(n_392), .B1(n_289), .B2(n_162), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_502), .A2(n_392), .B1(n_289), .B2(n_162), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_462), .A2(n_306), .B1(n_311), .B2(n_300), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_476), .A2(n_392), .B1(n_289), .B2(n_162), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_487), .A2(n_392), .B1(n_289), .B2(n_162), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_498), .B(n_162), .C(n_157), .Y(n_607) );
NAND2x1_ASAP7_75t_L g608 ( .A(n_487), .B(n_392), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_488), .A2(n_162), .B1(n_377), .B2(n_352), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_461), .A2(n_380), .B1(n_377), .B2(n_352), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_488), .A2(n_380), .B1(n_377), .B2(n_352), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_471), .A2(n_311), .B1(n_306), .B2(n_299), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_492), .A2(n_162), .B1(n_377), .B2(n_352), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g614 ( .A1(n_472), .A2(n_162), .B1(n_288), .B2(n_157), .C1(n_278), .C2(n_170), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_479), .A2(n_272), .B1(n_267), .B2(n_260), .C(n_261), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_471), .B(n_21), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_492), .A2(n_380), .B1(n_377), .B2(n_352), .Y(n_617) );
OAI211xp5_ASAP7_75t_SL g618 ( .A1(n_500), .A2(n_278), .B(n_288), .C(n_346), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_500), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_508), .A2(n_162), .B1(n_377), .B2(n_352), .Y(n_620) );
OAI222xp33_ASAP7_75t_L g621 ( .A1(n_508), .A2(n_157), .B1(n_286), .B2(n_24), .C1(n_26), .C2(n_27), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_526), .A2(n_380), .B1(n_377), .B2(n_307), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_466), .B(n_162), .Y(n_623) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_496), .A2(n_466), .B1(n_528), .B2(n_524), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_526), .A2(n_380), .B1(n_377), .B2(n_307), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_527), .B(n_22), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_475), .A2(n_162), .B1(n_380), .B2(n_299), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_475), .A2(n_380), .B1(n_299), .B2(n_300), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_475), .A2(n_380), .B1(n_299), .B2(n_300), .Y(n_629) );
OR2x6_ASAP7_75t_SL g630 ( .A(n_496), .B(n_23), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_527), .B(n_23), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_526), .B(n_24), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_526), .B(n_28), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_528), .A2(n_299), .B1(n_300), .B2(n_279), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_554), .B(n_478), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_590), .B(n_489), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_590), .B(n_489), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_546), .B(n_512), .Y(n_638) );
OA211x2_ASAP7_75t_L g639 ( .A1(n_630), .A2(n_30), .B(n_31), .C(n_32), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_559), .B(n_529), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_546), .B(n_512), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_555), .B(n_170), .C(n_530), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_572), .A2(n_537), .B1(n_614), .B2(n_538), .Y(n_643) );
OAI221xp5_ASAP7_75t_SL g644 ( .A1(n_593), .A2(n_530), .B1(n_271), .B2(n_306), .C(n_311), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_593), .B(n_243), .C(n_303), .D(n_34), .Y(n_645) );
AOI21xp33_ASAP7_75t_L g646 ( .A1(n_632), .A2(n_529), .B(n_170), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_630), .A2(n_529), .B1(n_307), .B2(n_157), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_588), .B(n_529), .Y(n_648) );
OAI221xp5_ASAP7_75t_SL g649 ( .A1(n_543), .A2(n_300), .B1(n_303), .B2(n_254), .C(n_239), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_555), .B(n_170), .C(n_157), .Y(n_650) );
AND2x2_ASAP7_75t_SL g651 ( .A(n_559), .B(n_170), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_559), .B(n_31), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_633), .A2(n_170), .B(n_35), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_557), .B(n_33), .Y(n_654) );
NAND4xp25_ASAP7_75t_L g655 ( .A(n_542), .B(n_303), .C(n_36), .D(n_37), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_534), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_549), .B(n_170), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_619), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_579), .B(n_36), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_544), .A2(n_170), .B1(n_279), .B2(n_157), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g661 ( .A(n_616), .B(n_303), .C(n_39), .D(n_40), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_534), .B(n_37), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_587), .B(n_39), .Y(n_663) );
NAND2xp33_ASAP7_75t_SL g664 ( .A(n_567), .B(n_307), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_604), .B(n_40), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_604), .B(n_41), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_607), .B(n_157), .C(n_279), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_621), .B(n_284), .C(n_344), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_581), .B(n_41), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_612), .B(n_42), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_612), .B(n_42), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_581), .B(n_43), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_581), .B(n_43), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_535), .B(n_157), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_536), .A2(n_325), .B(n_343), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_623), .B(n_157), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_581), .B(n_157), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_585), .B(n_157), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_623), .B(n_157), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_585), .B(n_157), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_626), .B(n_295), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_551), .A2(n_297), .B1(n_295), .B2(n_240), .Y(n_682) );
OAI21xp5_ASAP7_75t_SL g683 ( .A1(n_624), .A2(n_297), .B(n_295), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_607), .B(n_297), .C(n_295), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_631), .B(n_295), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_569), .B(n_297), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_583), .B(n_297), .C(n_343), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_585), .B(n_47), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_578), .B(n_343), .C(n_331), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g690 ( .A(n_541), .B(n_48), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_567), .A2(n_540), .B1(n_565), .B2(n_618), .Y(n_691) );
NAND4xp25_ASAP7_75t_L g692 ( .A(n_568), .B(n_251), .C(n_344), .D(n_329), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_539), .A2(n_307), .B1(n_239), .B2(n_344), .C(n_329), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_585), .B(n_49), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_574), .B(n_343), .C(n_331), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_568), .A2(n_343), .B1(n_331), .B2(n_315), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_608), .B(n_50), .Y(n_697) );
OA21x2_ASAP7_75t_L g698 ( .A1(n_592), .A2(n_328), .B(n_329), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_561), .B(n_331), .C(n_325), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_615), .B(n_328), .C(n_313), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_598), .B(n_51), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_608), .B(n_55), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g703 ( .A1(n_580), .A2(n_328), .B(n_325), .C(n_315), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_550), .B(n_325), .C(n_315), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_599), .B(n_325), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_599), .B(n_315), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_552), .B(n_322), .C(n_318), .Y(n_707) );
OAI22xp33_ASAP7_75t_L g708 ( .A1(n_577), .A2(n_322), .B1(n_318), .B2(n_313), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_586), .B(n_56), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_577), .B(n_59), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_582), .B(n_60), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_573), .B(n_61), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_600), .B(n_63), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_597), .B(n_64), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g715 ( .A1(n_584), .A2(n_322), .B1(n_318), .B2(n_313), .C(n_312), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_610), .B(n_66), .Y(n_716) );
OAI221xp5_ASAP7_75t_SL g717 ( .A1(n_565), .A2(n_312), .B1(n_247), .B2(n_70), .C(n_74), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_548), .B(n_312), .C(n_242), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_611), .B(n_67), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_617), .B(n_69), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_564), .A2(n_240), .B1(n_76), .B2(n_77), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_566), .B(n_75), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_595), .B(n_78), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g724 ( .A1(n_563), .A2(n_79), .B(n_80), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_589), .B(n_82), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_591), .B(n_83), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_545), .B(n_84), .Y(n_727) );
NAND3xp33_ASAP7_75t_SL g728 ( .A(n_556), .B(n_87), .C(n_89), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_628), .B(n_90), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_596), .B(n_91), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_622), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_629), .B(n_95), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_575), .B(n_96), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_609), .B(n_97), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_625), .B(n_98), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_613), .B(n_101), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_645), .A2(n_639), .B1(n_691), .B2(n_652), .Y(n_737) );
OAI211xp5_ASAP7_75t_SL g738 ( .A1(n_643), .A2(n_562), .B(n_553), .C(n_547), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_658), .B(n_620), .Y(n_739) );
NOR3xp33_ASAP7_75t_SL g740 ( .A(n_647), .B(n_560), .C(n_558), .Y(n_740) );
AO21x2_ASAP7_75t_L g741 ( .A1(n_654), .A2(n_606), .B(n_605), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_635), .B(n_601), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_661), .B(n_594), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_703), .B(n_603), .C(n_602), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_638), .Y(n_745) );
NAND4xp75_ASAP7_75t_L g746 ( .A(n_651), .B(n_576), .C(n_571), .D(n_634), .Y(n_746) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_657), .B(n_627), .C(n_570), .Y(n_747) );
NOR3xp33_ASAP7_75t_L g748 ( .A(n_655), .B(n_102), .C(n_103), .Y(n_748) );
XOR2x2_ASAP7_75t_L g749 ( .A(n_651), .B(n_104), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_641), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_636), .B(n_105), .Y(n_751) );
OAI211xp5_ASAP7_75t_SL g752 ( .A1(n_657), .A2(n_106), .B(n_108), .C(n_109), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_674), .B(n_110), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_648), .B(n_111), .Y(n_754) );
NOR3xp33_ASAP7_75t_L g755 ( .A(n_717), .B(n_112), .C(n_270), .Y(n_755) );
OR2x2_ASAP7_75t_L g756 ( .A(n_656), .B(n_648), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_669), .B(n_672), .Y(n_757) );
NAND4xp75_ASAP7_75t_L g758 ( .A(n_640), .B(n_735), .C(n_672), .D(n_673), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_690), .B(n_640), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_663), .B(n_665), .Y(n_760) );
AND2x4_ASAP7_75t_L g761 ( .A(n_669), .B(n_673), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_683), .B(n_642), .C(n_684), .Y(n_762) );
NOR3xp33_ASAP7_75t_SL g763 ( .A(n_644), .B(n_724), .C(n_664), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_663), .B(n_662), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g765 ( .A1(n_688), .A2(n_694), .B1(n_662), .B2(n_698), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_667), .A2(n_692), .B1(n_701), .B2(n_653), .Y(n_766) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_677), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_700), .A2(n_668), .B1(n_735), .B2(n_646), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_666), .B(n_671), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_708), .A2(n_670), .B1(n_664), .B2(n_675), .Y(n_770) );
NOR3xp33_ASAP7_75t_L g771 ( .A(n_659), .B(n_728), .C(n_693), .Y(n_771) );
INVx2_ASAP7_75t_SL g772 ( .A(n_712), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_678), .B(n_680), .Y(n_773) );
INVxp67_ASAP7_75t_R g774 ( .A(n_712), .Y(n_774) );
NAND3xp33_ASAP7_75t_L g775 ( .A(n_699), .B(n_682), .C(n_650), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_697), .B(n_702), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_649), .B(n_710), .Y(n_777) );
NAND3xp33_ASAP7_75t_L g778 ( .A(n_722), .B(n_731), .C(n_711), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_709), .B(n_716), .Y(n_779) );
OR2x2_ASAP7_75t_L g780 ( .A(n_681), .B(n_685), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_686), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_698), .Y(n_782) );
NAND4xp75_ASAP7_75t_L g783 ( .A(n_716), .B(n_698), .C(n_733), .D(n_709), .Y(n_783) );
NAND4xp75_ASAP7_75t_L g784 ( .A(n_729), .B(n_732), .C(n_723), .D(n_713), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_695), .A2(n_725), .B1(n_707), .B2(n_729), .Y(n_785) );
AND2x6_ASAP7_75t_L g786 ( .A(n_719), .B(n_720), .Y(n_786) );
AOI211xp5_ASAP7_75t_L g787 ( .A1(n_721), .A2(n_687), .B(n_689), .C(n_723), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_715), .B(n_676), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_719), .B(n_720), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g790 ( .A(n_713), .B(n_704), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_705), .Y(n_791) );
AOI22xp33_ASAP7_75t_SL g792 ( .A1(n_732), .A2(n_706), .B1(n_736), .B2(n_734), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_660), .A2(n_679), .B1(n_696), .B2(n_718), .C(n_725), .Y(n_793) );
AND2x2_ASAP7_75t_SL g794 ( .A(n_736), .B(n_714), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_730), .B(n_726), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_727), .A2(n_645), .B1(n_639), .B2(n_691), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_636), .B(n_637), .Y(n_797) );
NAND3xp33_ASAP7_75t_L g798 ( .A(n_658), .B(n_703), .C(n_554), .Y(n_798) );
NOR3xp33_ASAP7_75t_L g799 ( .A(n_661), .B(n_652), .C(n_645), .Y(n_799) );
NAND4xp25_ASAP7_75t_L g800 ( .A(n_639), .B(n_691), .C(n_643), .D(n_645), .Y(n_800) );
OA211x2_ASAP7_75t_L g801 ( .A1(n_657), .A2(n_640), .B(n_652), .C(n_735), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_635), .B(n_658), .Y(n_802) );
NAND4xp25_ASAP7_75t_L g803 ( .A(n_639), .B(n_691), .C(n_643), .D(n_645), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_658), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_658), .B(n_554), .Y(n_805) );
INVx4_ASAP7_75t_L g806 ( .A(n_786), .Y(n_806) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_756), .Y(n_807) );
XNOR2xp5_ASAP7_75t_L g808 ( .A(n_800), .B(n_803), .Y(n_808) );
NAND4xp75_ASAP7_75t_SL g809 ( .A(n_743), .B(n_777), .C(n_801), .D(n_779), .Y(n_809) );
BUFx2_ASAP7_75t_L g810 ( .A(n_767), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_745), .B(n_750), .Y(n_811) );
NAND4xp75_ASAP7_75t_SL g812 ( .A(n_749), .B(n_763), .C(n_795), .D(n_788), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g813 ( .A(n_765), .B(n_792), .Y(n_813) );
NAND4xp75_ASAP7_75t_L g814 ( .A(n_737), .B(n_796), .C(n_794), .D(n_759), .Y(n_814) );
INVx4_ASAP7_75t_L g815 ( .A(n_786), .Y(n_815) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_748), .B(n_799), .C(n_746), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_804), .Y(n_817) );
OR2x2_ASAP7_75t_L g818 ( .A(n_802), .B(n_805), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_805), .B(n_760), .Y(n_819) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_784), .B(n_764), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_799), .A2(n_748), .B1(n_774), .B2(n_786), .Y(n_821) );
NAND4xp75_ASAP7_75t_L g822 ( .A(n_770), .B(n_740), .C(n_769), .D(n_790), .Y(n_822) );
NOR4xp25_ASAP7_75t_L g823 ( .A(n_738), .B(n_768), .C(n_798), .D(n_766), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_757), .Y(n_824) );
INVx1_ASAP7_75t_SL g825 ( .A(n_751), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_761), .B(n_765), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_782), .Y(n_827) );
NAND4xp75_ASAP7_75t_L g828 ( .A(n_740), .B(n_789), .C(n_793), .D(n_772), .Y(n_828) );
NAND4xp75_ASAP7_75t_L g829 ( .A(n_793), .B(n_754), .C(n_739), .D(n_742), .Y(n_829) );
OR2x2_ASAP7_75t_L g830 ( .A(n_757), .B(n_780), .Y(n_830) );
XOR2x2_ASAP7_75t_L g831 ( .A(n_758), .B(n_783), .Y(n_831) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_773), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_781), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_791), .B(n_742), .Y(n_834) );
BUFx3_ASAP7_75t_L g835 ( .A(n_786), .Y(n_835) );
NAND4xp75_ASAP7_75t_SL g836 ( .A(n_776), .B(n_753), .C(n_755), .D(n_786), .Y(n_836) );
NAND4xp75_ASAP7_75t_L g837 ( .A(n_739), .B(n_778), .C(n_771), .D(n_755), .Y(n_837) );
BUFx12f_ASAP7_75t_L g838 ( .A(n_752), .Y(n_838) );
NAND4xp75_ASAP7_75t_L g839 ( .A(n_771), .B(n_792), .C(n_787), .D(n_762), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_741), .Y(n_840) );
NAND4xp75_ASAP7_75t_L g841 ( .A(n_775), .B(n_738), .C(n_744), .D(n_752), .Y(n_841) );
NOR4xp25_ASAP7_75t_L g842 ( .A(n_785), .B(n_800), .C(n_803), .D(n_645), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_741), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_747), .B(n_797), .Y(n_844) );
XNOR2x2_ASAP7_75t_L g845 ( .A(n_839), .B(n_808), .Y(n_845) );
XOR2x2_ASAP7_75t_L g846 ( .A(n_808), .B(n_812), .Y(n_846) );
OR2x2_ASAP7_75t_L g847 ( .A(n_834), .B(n_824), .Y(n_847) );
XNOR2xp5_ASAP7_75t_L g848 ( .A(n_831), .B(n_809), .Y(n_848) );
XNOR2x1_ASAP7_75t_L g849 ( .A(n_839), .B(n_822), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_811), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_811), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_817), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_817), .Y(n_853) );
XOR2x2_ASAP7_75t_L g854 ( .A(n_812), .B(n_809), .Y(n_854) );
INVx1_ASAP7_75t_SL g855 ( .A(n_810), .Y(n_855) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_810), .Y(n_856) );
INVx2_ASAP7_75t_SL g857 ( .A(n_835), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_827), .Y(n_858) );
CKINVDCx16_ASAP7_75t_R g859 ( .A(n_806), .Y(n_859) );
NOR2x1_ASAP7_75t_L g860 ( .A(n_814), .B(n_828), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_806), .A2(n_815), .B1(n_821), .B2(n_835), .Y(n_861) );
OR2x2_ASAP7_75t_L g862 ( .A(n_834), .B(n_830), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_833), .Y(n_863) );
INVxp67_ASAP7_75t_L g864 ( .A(n_814), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_833), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_830), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_826), .B(n_844), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_844), .B(n_840), .Y(n_868) );
OR2x2_ASAP7_75t_L g869 ( .A(n_807), .B(n_824), .Y(n_869) );
XNOR2x1_ASAP7_75t_L g870 ( .A(n_822), .B(n_828), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_832), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_818), .Y(n_872) );
XNOR2x1_ASAP7_75t_L g873 ( .A(n_831), .B(n_841), .Y(n_873) );
AO22x2_ASAP7_75t_L g874 ( .A1(n_873), .A2(n_829), .B1(n_840), .B2(n_813), .Y(n_874) );
INVx2_ASAP7_75t_SL g875 ( .A(n_859), .Y(n_875) );
OA22x2_ASAP7_75t_L g876 ( .A1(n_848), .A2(n_821), .B1(n_820), .B2(n_806), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_870), .A2(n_806), .B1(n_815), .B2(n_835), .Y(n_877) );
OA22x2_ASAP7_75t_L g878 ( .A1(n_864), .A2(n_820), .B1(n_815), .B2(n_826), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_856), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g880 ( .A1(n_849), .A2(n_816), .B1(n_831), .B2(n_829), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_862), .Y(n_881) );
NOR2x1_ASAP7_75t_R g882 ( .A(n_845), .B(n_838), .Y(n_882) );
OA22x2_ASAP7_75t_L g883 ( .A1(n_861), .A2(n_815), .B1(n_843), .B2(n_842), .Y(n_883) );
INVx5_ASAP7_75t_L g884 ( .A(n_854), .Y(n_884) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_873), .B(n_841), .Y(n_885) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_857), .A2(n_838), .B1(n_825), .B2(n_807), .Y(n_886) );
AOI22xp5_ASAP7_75t_SL g887 ( .A1(n_857), .A2(n_819), .B1(n_836), .B2(n_825), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_849), .A2(n_816), .B1(n_842), .B2(n_837), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_871), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_880), .A2(n_870), .B1(n_860), .B2(n_867), .Y(n_890) );
HB1xp67_ASAP7_75t_L g891 ( .A(n_879), .Y(n_891) );
CKINVDCx14_ASAP7_75t_R g892 ( .A(n_884), .Y(n_892) );
INVx2_ASAP7_75t_SL g893 ( .A(n_875), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_881), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_889), .Y(n_895) );
BUFx2_ASAP7_75t_L g896 ( .A(n_882), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_883), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_877), .Y(n_898) );
AO22x2_ASAP7_75t_L g899 ( .A1(n_893), .A2(n_845), .B1(n_855), .B2(n_874), .Y(n_899) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_890), .A2(n_888), .B1(n_885), .B2(n_876), .Y(n_900) );
AOI221xp5_ASAP7_75t_L g901 ( .A1(n_898), .A2(n_874), .B1(n_823), .B2(n_884), .C(n_886), .Y(n_901) );
AND4x1_ASAP7_75t_L g902 ( .A(n_898), .B(n_823), .C(n_846), .D(n_854), .Y(n_902) );
OA22x2_ASAP7_75t_L g903 ( .A1(n_896), .A2(n_846), .B1(n_878), .B2(n_867), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_899), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_903), .A2(n_896), .B1(n_893), .B2(n_892), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g906 ( .A1(n_900), .A2(n_897), .B1(n_894), .B2(n_837), .Y(n_906) );
NOR2x1_ASAP7_75t_L g907 ( .A(n_904), .B(n_897), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_905), .A2(n_901), .B1(n_894), .B2(n_891), .Y(n_908) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_906), .Y(n_909) );
INVxp67_ASAP7_75t_L g910 ( .A(n_907), .Y(n_910) );
INVx1_ASAP7_75t_SL g911 ( .A(n_908), .Y(n_911) );
NOR4xp25_ASAP7_75t_L g912 ( .A(n_911), .B(n_909), .C(n_902), .D(n_895), .Y(n_912) );
NOR4xp25_ASAP7_75t_L g913 ( .A(n_910), .B(n_868), .C(n_843), .D(n_851), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_912), .Y(n_914) );
INVx1_ASAP7_75t_SL g915 ( .A(n_913), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_914), .A2(n_887), .B1(n_856), .B2(n_872), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_916), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_917), .A2(n_914), .B1(n_915), .B2(n_866), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_918), .Y(n_919) );
AOI22xp5_ASAP7_75t_SL g920 ( .A1(n_919), .A2(n_850), .B1(n_843), .B2(n_865), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_920), .Y(n_921) );
AOI221x1_ASAP7_75t_L g922 ( .A1(n_921), .A2(n_863), .B1(n_853), .B2(n_852), .C(n_858), .Y(n_922) );
AOI211xp5_ASAP7_75t_L g923 ( .A1(n_922), .A2(n_847), .B(n_818), .C(n_869), .Y(n_923) );
endmodule