module real_aes_7125_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g457 ( .A1(n_0), .A2(n_158), .B(n_458), .C(n_461), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_1), .B(n_452), .Y(n_462) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g120 ( .A(n_2), .Y(n_120) );
INVx1_ASAP7_75t_L g156 ( .A(n_3), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_4), .B(n_159), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_5), .A2(n_447), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_6), .A2(n_181), .B(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_7), .A2(n_38), .B1(n_146), .B2(n_204), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_8), .A2(n_9), .B1(n_709), .B2(n_710), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_8), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_9), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_10), .B(n_181), .Y(n_189) );
AND2x6_ASAP7_75t_L g161 ( .A(n_11), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_12), .A2(n_161), .B(n_438), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_13), .B(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_13), .B(n_39), .Y(n_121) );
INVx1_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
INVx1_ASAP7_75t_L g137 ( .A(n_15), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_16), .B(n_142), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_17), .B(n_159), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_18), .B(n_133), .Y(n_191) );
AO32x2_ASAP7_75t_L g242 ( .A1(n_19), .A2(n_132), .A3(n_175), .B1(n_181), .B2(n_243), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_20), .A2(n_30), .B1(n_123), .B2(n_730), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_20), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_21), .B(n_146), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_22), .B(n_133), .Y(n_163) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_23), .A2(n_56), .B1(n_146), .B2(n_204), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g206 ( .A1(n_24), .A2(n_81), .B1(n_142), .B2(n_146), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_25), .B(n_146), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_26), .A2(n_175), .B(n_438), .C(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_27), .A2(n_175), .B(n_438), .C(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_28), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_29), .B(n_177), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_30), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_30), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_31), .A2(n_447), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_32), .B(n_177), .Y(n_219) );
INVx2_ASAP7_75t_L g144 ( .A(n_33), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_34), .A2(n_444), .B(n_487), .C(n_488), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_35), .B(n_146), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_36), .B(n_177), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_37), .B(n_226), .Y(n_532) );
INVx1_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_40), .B(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_41), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_42), .A2(n_103), .B1(n_114), .B2(n_738), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_43), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_44), .B(n_159), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_45), .B(n_447), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_46), .A2(n_444), .B(n_487), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_47), .B(n_146), .Y(n_184) );
INVx1_ASAP7_75t_L g459 ( .A(n_48), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_49), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_50), .A2(n_90), .B1(n_204), .B2(n_205), .Y(n_203) );
INVx1_ASAP7_75t_L g512 ( .A(n_51), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_52), .B(n_146), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_53), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_54), .B(n_447), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_55), .B(n_154), .Y(n_188) );
AOI22xp33_ASAP7_75t_SL g195 ( .A1(n_57), .A2(n_61), .B1(n_142), .B2(n_146), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_58), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_59), .B(n_146), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_60), .B(n_146), .Y(n_223) );
INVx1_ASAP7_75t_L g162 ( .A(n_62), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_63), .B(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_64), .B(n_452), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_65), .A2(n_148), .B(n_154), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_66), .B(n_146), .Y(n_157) );
INVx1_ASAP7_75t_L g136 ( .A(n_67), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_68), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_69), .B(n_159), .Y(n_490) );
AO32x2_ASAP7_75t_L g201 ( .A1(n_70), .A2(n_175), .A3(n_181), .B1(n_202), .B2(n_207), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_71), .B(n_160), .Y(n_503) );
INVx1_ASAP7_75t_L g171 ( .A(n_72), .Y(n_171) );
INVx1_ASAP7_75t_L g214 ( .A(n_73), .Y(n_214) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_74), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_75), .B(n_471), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g437 ( .A1(n_76), .A2(n_438), .B(n_440), .C(n_444), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_77), .B(n_142), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_78), .Y(n_521) );
INVx1_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_80), .B(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_82), .B(n_204), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_83), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_84), .B(n_142), .Y(n_218) );
INVx2_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_86), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_87), .B(n_174), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_88), .B(n_142), .Y(n_185) );
INVx2_ASAP7_75t_L g110 ( .A(n_89), .Y(n_110) );
OR2x2_ASAP7_75t_L g118 ( .A(n_89), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g726 ( .A(n_89), .B(n_718), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_91), .A2(n_101), .B1(n_142), .B2(n_143), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_92), .B(n_447), .Y(n_485) );
INVx1_ASAP7_75t_L g489 ( .A(n_93), .Y(n_489) );
INVxp67_ASAP7_75t_L g524 ( .A(n_94), .Y(n_524) );
XNOR2xp5_ASAP7_75t_L g727 ( .A(n_95), .B(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_96), .B(n_142), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_97), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g441 ( .A(n_98), .Y(n_441) );
INVx1_ASAP7_75t_L g499 ( .A(n_99), .Y(n_499) );
AND2x2_ASAP7_75t_L g514 ( .A(n_100), .B(n_177), .Y(n_514) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx12_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g739 ( .A(n_106), .Y(n_739) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
OR2x2_ASAP7_75t_L g429 ( .A(n_110), .B(n_119), .Y(n_429) );
NOR2x2_ASAP7_75t_L g717 ( .A(n_110), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO221x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_720), .B1(n_723), .B2(n_732), .C(n_734), .Y(n_114) );
OAI222xp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_708), .B1(n_711), .B2(n_715), .C1(n_716), .C2(n_719), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B1(n_428), .B2(n_430), .Y(n_116) );
INVx2_ASAP7_75t_L g713 ( .A(n_117), .Y(n_713) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g718 ( .A(n_119), .Y(n_718) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_122), .A2(n_430), .B1(n_713), .B2(n_714), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_124), .A2(n_125), .B1(n_729), .B2(n_731), .Y(n_728) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR5x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_319), .C(n_377), .D(n_413), .E(n_420), .Y(n_125) );
NAND3xp33_ASAP7_75t_SL g126 ( .A(n_127), .B(n_265), .C(n_289), .Y(n_126) );
AOI221xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_197), .B1(n_231), .B2(n_236), .C(n_246), .Y(n_127) );
OAI21xp5_ASAP7_75t_SL g399 ( .A1(n_128), .A2(n_400), .B(n_402), .Y(n_399) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_178), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g389 ( .A(n_129), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_164), .Y(n_129) );
INVx2_ASAP7_75t_L g235 ( .A(n_130), .Y(n_235) );
AND2x2_ASAP7_75t_L g248 ( .A(n_130), .B(n_180), .Y(n_248) );
AND2x2_ASAP7_75t_L g302 ( .A(n_130), .B(n_179), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_130), .B(n_165), .Y(n_317) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_163), .Y(n_130) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_131), .A2(n_166), .B(n_176), .Y(n_165) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_132), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_133), .Y(n_181) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_134), .B(n_135), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_152), .B(n_161), .Y(n_138) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B(n_145), .C(n_148), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_141), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_141), .A2(n_532), .B(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
INVx1_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
INVx3_ASAP7_75t_L g213 ( .A(n_146), .Y(n_213) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_146), .Y(n_443) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g204 ( .A(n_147), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
AND2x6_ASAP7_75t_L g438 ( .A(n_147), .B(n_439), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_148), .A2(n_441), .B(n_442), .C(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_149), .A2(n_217), .B(n_218), .Y(n_216) );
INVx4_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g471 ( .A(n_150), .Y(n_471) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g160 ( .A(n_151), .Y(n_160) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
INVx1_ASAP7_75t_L g226 ( .A(n_151), .Y(n_226) );
INVx1_ASAP7_75t_L g439 ( .A(n_151), .Y(n_439) );
AND2x2_ASAP7_75t_L g448 ( .A(n_151), .B(n_155), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_156), .B(n_157), .C(n_158), .Y(n_152) );
O2A1O1Ixp5_ASAP7_75t_L g170 ( .A1(n_153), .A2(n_171), .B(n_172), .C(n_173), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_153), .A2(n_470), .B(n_472), .Y(n_469) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_158), .A2(n_187), .B(n_188), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_158), .A2(n_174), .B1(n_194), .B2(n_195), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_158), .A2(n_174), .B1(n_244), .B2(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_159), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_159), .A2(n_184), .B(n_185), .Y(n_183) );
O2A1O1Ixp5_ASAP7_75t_SL g212 ( .A1(n_159), .A2(n_213), .B(n_214), .C(n_215), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_159), .B(n_524), .Y(n_523) );
INVx5_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g202 ( .A1(n_160), .A2(n_174), .B1(n_203), .B2(n_206), .Y(n_202) );
BUFx3_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_161), .A2(n_183), .B(n_186), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_161), .A2(n_212), .B(n_216), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_161), .A2(n_222), .B(n_227), .Y(n_221) );
INVx4_ASAP7_75t_SL g445 ( .A(n_161), .Y(n_445) );
AND2x4_ASAP7_75t_L g447 ( .A(n_161), .B(n_448), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_161), .B(n_448), .Y(n_500) );
AND2x2_ASAP7_75t_L g335 ( .A(n_164), .B(n_276), .Y(n_335) );
AND2x2_ASAP7_75t_L g368 ( .A(n_164), .B(n_180), .Y(n_368) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OR2x2_ASAP7_75t_L g275 ( .A(n_165), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g288 ( .A(n_165), .B(n_180), .Y(n_288) );
AND2x2_ASAP7_75t_L g295 ( .A(n_165), .B(n_276), .Y(n_295) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_165), .Y(n_304) );
AND2x2_ASAP7_75t_L g311 ( .A(n_165), .B(n_179), .Y(n_311) );
INVx1_ASAP7_75t_L g342 ( .A(n_165), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_175), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_173), .A2(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g460 ( .A(n_174), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_175), .B(n_193), .C(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g207 ( .A(n_177), .Y(n_207) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_177), .A2(n_211), .B(n_219), .Y(n_210) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_177), .A2(n_221), .B(n_230), .Y(n_220) );
INVx1_ASAP7_75t_L g477 ( .A(n_177), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_177), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_177), .A2(n_509), .B(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g318 ( .A(n_178), .Y(n_318) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_190), .Y(n_178) );
INVx2_ASAP7_75t_L g274 ( .A(n_179), .Y(n_274) );
AND2x2_ASAP7_75t_L g296 ( .A(n_179), .B(n_235), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_179), .B(n_342), .Y(n_347) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_180), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g419 ( .A(n_180), .B(n_383), .Y(n_419) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_189), .Y(n_180) );
INVx4_ASAP7_75t_L g196 ( .A(n_181), .Y(n_196) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_181), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_181), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g233 ( .A(n_190), .Y(n_233) );
INVx3_ASAP7_75t_L g334 ( .A(n_190), .Y(n_334) );
OR2x2_ASAP7_75t_L g364 ( .A(n_190), .B(n_365), .Y(n_364) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_190), .B(n_274), .Y(n_390) );
AND2x4_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g277 ( .A(n_191), .Y(n_277) );
AO21x1_ASAP7_75t_L g276 ( .A1(n_193), .A2(n_196), .B(n_277), .Y(n_276) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_196), .A2(n_436), .B(n_449), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_196), .B(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g452 ( .A(n_196), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_196), .B(n_493), .Y(n_492) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_196), .A2(n_498), .B(n_505), .Y(n_497) );
AOI33xp33_ASAP7_75t_L g410 ( .A1(n_197), .A2(n_248), .A3(n_262), .B1(n_334), .B2(n_411), .B3(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_208), .Y(n_198) );
OR2x2_ASAP7_75t_L g263 ( .A(n_199), .B(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_199), .B(n_260), .Y(n_322) );
OR2x2_ASAP7_75t_L g375 ( .A(n_199), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g301 ( .A(n_200), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g326 ( .A(n_200), .B(n_208), .Y(n_326) );
AND2x2_ASAP7_75t_L g393 ( .A(n_200), .B(n_238), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_200), .A2(n_293), .B(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g240 ( .A(n_201), .Y(n_240) );
INVx1_ASAP7_75t_L g253 ( .A(n_201), .Y(n_253) );
AND2x2_ASAP7_75t_L g272 ( .A(n_201), .B(n_242), .Y(n_272) );
AND2x2_ASAP7_75t_L g321 ( .A(n_201), .B(n_241), .Y(n_321) );
INVx2_ASAP7_75t_L g461 ( .A(n_205), .Y(n_461) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_205), .Y(n_491) );
INVx1_ASAP7_75t_L g474 ( .A(n_207), .Y(n_474) );
INVx2_ASAP7_75t_SL g363 ( .A(n_208), .Y(n_363) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
INVx2_ASAP7_75t_L g283 ( .A(n_209), .Y(n_283) );
INVx1_ASAP7_75t_L g414 ( .A(n_209), .Y(n_414) );
AND2x2_ASAP7_75t_L g427 ( .A(n_209), .B(n_308), .Y(n_427) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g254 ( .A(n_210), .Y(n_254) );
OR2x2_ASAP7_75t_L g260 ( .A(n_210), .B(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_210), .Y(n_271) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_220), .Y(n_238) );
AND2x2_ASAP7_75t_L g255 ( .A(n_220), .B(n_241), .Y(n_255) );
INVx1_ASAP7_75t_L g261 ( .A(n_220), .Y(n_261) );
INVx1_ASAP7_75t_L g268 ( .A(n_220), .Y(n_268) );
AND2x2_ASAP7_75t_L g293 ( .A(n_220), .B(n_242), .Y(n_293) );
INVx2_ASAP7_75t_L g309 ( .A(n_220), .Y(n_309) );
AND2x2_ASAP7_75t_L g402 ( .A(n_220), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_220), .B(n_283), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g257 ( .A(n_233), .Y(n_257) );
INVx1_ASAP7_75t_L g286 ( .A(n_233), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_233), .B(n_317), .Y(n_383) );
INVx1_ASAP7_75t_SL g343 ( .A(n_234), .Y(n_343) );
INVx2_ASAP7_75t_L g264 ( .A(n_235), .Y(n_264) );
AND2x2_ASAP7_75t_L g333 ( .A(n_235), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g349 ( .A(n_235), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
INVx1_ASAP7_75t_L g411 ( .A(n_237), .Y(n_411) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g266 ( .A(n_239), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g369 ( .A(n_239), .B(n_359), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_239), .A2(n_380), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AND2x2_ASAP7_75t_L g282 ( .A(n_240), .B(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g307 ( .A(n_240), .Y(n_307) );
INVx1_ASAP7_75t_L g331 ( .A(n_240), .Y(n_331) );
OR2x2_ASAP7_75t_L g395 ( .A(n_241), .B(n_254), .Y(n_395) );
NOR2xp67_ASAP7_75t_L g403 ( .A(n_241), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g308 ( .A(n_242), .B(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g315 ( .A(n_242), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B1(n_256), .B2(n_258), .Y(n_246) );
OR2x2_ASAP7_75t_L g325 ( .A(n_247), .B(n_275), .Y(n_325) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_248), .A2(n_367), .B1(n_369), .B2(n_370), .C1(n_371), .C2(n_374), .Y(n_366) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g313 ( .A(n_252), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_254), .B(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_254), .Y(n_338) );
AND2x2_ASAP7_75t_L g386 ( .A(n_254), .B(n_255), .Y(n_386) );
INVx1_ASAP7_75t_L g404 ( .A(n_254), .Y(n_404) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g370 ( .A(n_257), .B(n_296), .Y(n_370) );
AND2x2_ASAP7_75t_L g412 ( .A(n_257), .B(n_288), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_259), .B(n_307), .Y(n_394) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_260), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g287 ( .A(n_264), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g355 ( .A(n_264), .Y(n_355) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .B(n_273), .C(n_278), .Y(n_265) );
INVxp67_ASAP7_75t_L g279 ( .A(n_266), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_267), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_267), .B(n_314), .Y(n_409) );
BUFx3_ASAP7_75t_L g373 ( .A(n_268), .Y(n_373) );
INVx1_ASAP7_75t_L g280 ( .A(n_269), .Y(n_280) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g299 ( .A(n_271), .B(n_293), .Y(n_299) );
INVx1_ASAP7_75t_SL g339 ( .A(n_272), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g329 ( .A(n_274), .Y(n_329) );
AND2x2_ASAP7_75t_L g352 ( .A(n_274), .B(n_335), .Y(n_352) );
INVx1_ASAP7_75t_SL g323 ( .A(n_275), .Y(n_323) );
INVx1_ASAP7_75t_L g350 ( .A(n_276), .Y(n_350) );
AOI31xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .A3(n_281), .B(n_284), .Y(n_278) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g371 ( .A(n_282), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g345 ( .A(n_283), .Y(n_345) );
BUFx2_ASAP7_75t_L g359 ( .A(n_283), .Y(n_359) );
AND2x2_ASAP7_75t_L g387 ( .A(n_283), .B(n_308), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g360 ( .A(n_287), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_288), .B(n_355), .Y(n_401) );
AND2x2_ASAP7_75t_L g408 ( .A(n_288), .B(n_334), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_294), .B(n_297), .C(n_312), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_294), .A2(n_321), .B1(n_322), .B2(n_323), .C(n_324), .Y(n_320) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g328 ( .A(n_295), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g365 ( .A(n_296), .Y(n_365) );
OAI32xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_300), .A3(n_303), .B1(n_305), .B2(n_310), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_299), .A2(n_352), .B(n_353), .C(n_356), .Y(n_351) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_307), .A2(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g376 ( .A(n_308), .Y(n_376) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_314), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g362 ( .A(n_314), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g379 ( .A(n_316), .Y(n_379) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND4xp25_ASAP7_75t_SL g319 ( .A(n_320), .B(n_332), .C(n_351), .D(n_366), .Y(n_319) );
AND2x2_ASAP7_75t_L g358 ( .A(n_321), .B(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g380 ( .A(n_321), .B(n_373), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_323), .B(n_355), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_327), .B2(n_330), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_325), .A2(n_376), .B1(n_407), .B2(n_409), .Y(n_406) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_325), .A2(n_414), .B(n_415), .C(n_418), .Y(n_413) );
INVx2_ASAP7_75t_L g384 ( .A(n_326), .Y(n_384) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_328), .A2(n_362), .B1(n_379), .B2(n_380), .C1(n_381), .C2(n_384), .Y(n_378) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_336), .C(n_340), .Y(n_332) );
INVx1_ASAP7_75t_L g398 ( .A(n_333), .Y(n_398) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_337), .A2(n_341), .B1(n_344), .B2(n_346), .Y(n_340) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g367 ( .A(n_349), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g425 ( .A(n_352), .Y(n_425) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B1(n_361), .B2(n_364), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_359), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g416 ( .A(n_364), .Y(n_416) );
INVx1_ASAP7_75t_L g397 ( .A(n_368), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_370), .Y(n_424) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND5xp2_ASAP7_75t_L g377 ( .A(n_378), .B(n_385), .C(n_399), .D(n_405), .E(n_410), .Y(n_377) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_388), .C(n_391), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI31xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .A3(n_395), .B(n_396), .Y(n_391) );
INVx1_ASAP7_75t_L g417 ( .A(n_393), .Y(n_417) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI222xp33_ASAP7_75t_L g420 ( .A1(n_407), .A2(n_409), .B1(n_421), .B2(n_424), .C1(n_425), .C2(n_426), .Y(n_420) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g714 ( .A(n_428), .Y(n_714) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR3x1_ASAP7_75t_L g430 ( .A(n_431), .B(n_616), .C(n_665), .Y(n_430) );
NAND5xp2_ASAP7_75t_L g431 ( .A(n_432), .B(n_550), .C(n_579), .D(n_587), .E(n_602), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_478), .B(n_494), .C(n_534), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_463), .Y(n_433) );
AND2x2_ASAP7_75t_L g545 ( .A(n_434), .B(n_542), .Y(n_545) );
AND2x2_ASAP7_75t_L g578 ( .A(n_434), .B(n_464), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_434), .B(n_482), .Y(n_671) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_451), .Y(n_434) );
INVx2_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
BUFx2_ASAP7_75t_L g645 ( .A(n_435), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_446), .Y(n_436) );
INVx5_ASAP7_75t_L g456 ( .A(n_438), .Y(n_456) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_SL g454 ( .A1(n_445), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_445), .A2(n_456), .B(n_521), .C(n_522), .Y(n_520) );
BUFx2_ASAP7_75t_L g467 ( .A(n_447), .Y(n_467) );
AND2x2_ASAP7_75t_L g463 ( .A(n_451), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g543 ( .A(n_451), .Y(n_543) );
AND2x2_ASAP7_75t_L g629 ( .A(n_451), .B(n_542), .Y(n_629) );
AND2x2_ASAP7_75t_L g684 ( .A(n_451), .B(n_481), .Y(n_684) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_462), .Y(n_451) );
INVx2_ASAP7_75t_L g487 ( .A(n_456), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g601 ( .A(n_463), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_463), .B(n_482), .Y(n_648) );
INVx5_ASAP7_75t_L g542 ( .A(n_464), .Y(n_542) );
AND2x4_ASAP7_75t_L g563 ( .A(n_464), .B(n_543), .Y(n_563) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_464), .Y(n_585) );
AND2x2_ASAP7_75t_L g660 ( .A(n_464), .B(n_645), .Y(n_660) );
AND2x2_ASAP7_75t_L g663 ( .A(n_464), .B(n_483), .Y(n_663) );
OR2x6_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
AOI21xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_468), .B(n_474), .Y(n_465) );
INVx2_ASAP7_75t_L g473 ( .A(n_471), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_473), .A2(n_489), .B(n_490), .C(n_491), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_473), .A2(n_491), .B(n_512), .C(n_513), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_478), .B(n_543), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_478), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
AND2x2_ASAP7_75t_L g568 ( .A(n_480), .B(n_543), .Y(n_568) );
AND2x2_ASAP7_75t_L g586 ( .A(n_480), .B(n_483), .Y(n_586) );
INVx1_ASAP7_75t_L g606 ( .A(n_480), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_480), .B(n_542), .Y(n_651) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_480), .Y(n_693) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_481), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_482), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_482), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_482), .A2(n_538), .B(n_599), .C(n_601), .Y(n_598) );
AND2x2_ASAP7_75t_L g605 ( .A(n_482), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g614 ( .A(n_482), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g618 ( .A(n_482), .B(n_542), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_482), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g633 ( .A(n_482), .B(n_543), .Y(n_633) );
AND2x2_ASAP7_75t_L g683 ( .A(n_482), .B(n_684), .Y(n_683) );
INVx5_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g547 ( .A(n_483), .Y(n_547) );
AND2x2_ASAP7_75t_L g588 ( .A(n_483), .B(n_541), .Y(n_588) );
AND2x2_ASAP7_75t_L g600 ( .A(n_483), .B(n_575), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_483), .B(n_629), .Y(n_647) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_492), .Y(n_483) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_515), .Y(n_494) );
INVx1_ASAP7_75t_L g536 ( .A(n_495), .Y(n_536) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_507), .Y(n_495) );
OR2x2_ASAP7_75t_L g538 ( .A(n_496), .B(n_507), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_496), .B(n_545), .C(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_496), .B(n_517), .Y(n_555) );
OR2x2_ASAP7_75t_L g570 ( .A(n_496), .B(n_558), .Y(n_570) );
AND2x2_ASAP7_75t_L g576 ( .A(n_496), .B(n_526), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_496), .B(n_707), .Y(n_706) );
INVx5_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_497), .B(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g612 ( .A(n_497), .B(n_527), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_497), .B(n_526), .Y(n_640) );
OR2x2_ASAP7_75t_L g643 ( .A(n_497), .B(n_526), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B(n_501), .Y(n_498) );
INVx5_ASAP7_75t_SL g558 ( .A(n_507), .Y(n_558) );
OR2x2_ASAP7_75t_L g564 ( .A(n_507), .B(n_516), .Y(n_564) );
AND2x2_ASAP7_75t_L g580 ( .A(n_507), .B(n_581), .Y(n_580) );
AOI321xp33_ASAP7_75t_L g587 ( .A1(n_507), .A2(n_588), .A3(n_589), .B1(n_590), .B2(n_596), .C(n_598), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_507), .B(n_515), .Y(n_597) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_507), .Y(n_610) );
OR2x2_ASAP7_75t_L g657 ( .A(n_507), .B(n_555), .Y(n_657) );
AND2x2_ASAP7_75t_L g679 ( .A(n_507), .B(n_576), .Y(n_679) );
AND2x2_ASAP7_75t_L g698 ( .A(n_507), .B(n_517), .Y(n_698) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
INVx1_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_526), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_517), .B(n_526), .Y(n_539) );
AND2x2_ASAP7_75t_L g548 ( .A(n_517), .B(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g575 ( .A(n_517), .Y(n_575) );
AND2x2_ASAP7_75t_L g581 ( .A(n_517), .B(n_576), .Y(n_581) );
INVxp67_ASAP7_75t_L g611 ( .A(n_517), .Y(n_611) );
OR2x2_ASAP7_75t_L g653 ( .A(n_517), .B(n_558), .Y(n_653) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_525), .Y(n_517) );
OR2x2_ASAP7_75t_L g535 ( .A(n_526), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_SL g549 ( .A(n_526), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_526), .B(n_538), .Y(n_582) );
AND2x2_ASAP7_75t_L g631 ( .A(n_526), .B(n_575), .Y(n_631) );
AND2x2_ASAP7_75t_L g669 ( .A(n_526), .B(n_558), .Y(n_669) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_527), .B(n_558), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_537), .B(n_540), .C(n_544), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_535), .A2(n_537), .B1(n_662), .B2(n_664), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_537), .A2(n_560), .B1(n_615), .B2(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_SL g689 ( .A(n_538), .Y(n_689) );
INVx1_ASAP7_75t_SL g589 ( .A(n_539), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_541), .B(n_561), .Y(n_591) );
AOI222xp33_ASAP7_75t_L g602 ( .A1(n_541), .A2(n_582), .B1(n_589), .B2(n_603), .C1(n_607), .C2(n_613), .Y(n_602) );
AND2x2_ASAP7_75t_L g692 ( .A(n_541), .B(n_693), .Y(n_692) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g567 ( .A(n_542), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_542), .B(n_562), .Y(n_637) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_542), .Y(n_674) );
AND2x2_ASAP7_75t_L g677 ( .A(n_542), .B(n_586), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_542), .B(n_693), .Y(n_703) );
INVx1_ASAP7_75t_L g594 ( .A(n_543), .Y(n_594) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_543), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_L g685 ( .A1(n_545), .A2(n_686), .B(n_687), .C(n_690), .Y(n_685) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_547), .B(n_609), .C(n_612), .Y(n_608) );
OR2x2_ASAP7_75t_L g636 ( .A(n_547), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_547), .B(n_563), .Y(n_664) );
OR2x2_ASAP7_75t_L g569 ( .A(n_549), .B(n_570), .Y(n_569) );
AOI211xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_553), .B(n_559), .C(n_571), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_552), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g658 ( .A(n_553), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_554), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g572 ( .A(n_557), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_558), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g626 ( .A(n_558), .B(n_576), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_558), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_558), .B(n_575), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_564), .B1(n_565), .B2(n_569), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_561), .B(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_563), .B(n_605), .Y(n_604) );
OAI221xp5_ASAP7_75t_SL g627 ( .A1(n_564), .A2(n_628), .B1(n_630), .B2(n_632), .C(n_634), .Y(n_627) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x2_ASAP7_75t_L g682 ( .A(n_567), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g695 ( .A(n_567), .B(n_684), .Y(n_695) );
INVx1_ASAP7_75t_L g615 ( .A(n_568), .Y(n_615) );
INVx1_ASAP7_75t_L g686 ( .A(n_569), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_570), .A2(n_653), .B(n_676), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B(n_577), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI21xp5_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_582), .B(n_583), .Y(n_579) );
INVx1_ASAP7_75t_L g619 ( .A(n_580), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_581), .A2(n_667), .B1(n_670), .B2(n_672), .C(n_675), .Y(n_666) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_589), .A2(n_679), .B1(n_680), .B2(n_682), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g655 ( .A(n_591), .Y(n_655) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp67_ASAP7_75t_SL g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g659 ( .A(n_595), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g624 ( .A(n_600), .Y(n_624) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_605), .B(n_629), .Y(n_681) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_611), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g697 ( .A(n_612), .B(n_698), .Y(n_697) );
AND2x4_ASAP7_75t_L g704 ( .A(n_612), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI211xp5_ASAP7_75t_SL g616 ( .A1(n_617), .A2(n_619), .B(n_620), .C(n_654), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI211xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B(n_627), .C(n_646), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_SL g707 ( .A(n_631), .Y(n_707) );
AND2x2_ASAP7_75t_L g644 ( .A(n_633), .B(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_638), .B1(n_642), .B2(n_644), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
OR2x2_ASAP7_75t_L g652 ( .A(n_640), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g705 ( .A(n_641), .Y(n_705) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI31xp33_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .A3(n_649), .B(n_652), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B(n_658), .C(n_661), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
CKINVDCx16_ASAP7_75t_R g662 ( .A(n_663), .Y(n_662) );
NAND5xp2_ASAP7_75t_L g665 ( .A(n_666), .B(n_678), .C(n_685), .D(n_699), .E(n_702), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_677), .A2(n_703), .B1(n_704), .B2(n_706), .Y(n_702) );
INVx1_ASAP7_75t_SL g701 ( .A(n_679), .Y(n_701) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_694), .B(n_696), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g715 ( .A(n_708), .Y(n_715) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
BUFx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_SL g733 ( .A(n_721), .Y(n_733) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
BUFx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g737 ( .A(n_726), .Y(n_737) );
INVx1_ASAP7_75t_L g731 ( .A(n_729), .Y(n_731) );
BUFx3_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
endmodule