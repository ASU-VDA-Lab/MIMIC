module fake_jpeg_24940_n_22 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_22);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_22;

wire n_13;
wire n_21;
wire n_10;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;

INVxp67_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_2),
.B(n_6),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_0),
.Y(n_10)
);

OR2x4_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_2),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_0),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_11),
.A2(n_3),
.B1(n_5),
.B2(n_12),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_19),
.B1(n_8),
.B2(n_17),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_5),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_17),
.A2(n_18),
.B1(n_8),
.B2(n_9),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_21),
.Y(n_22)
);


endmodule