module real_jpeg_23653_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_33),
.B1(n_38),
.B2(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_1),
.A2(n_33),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_1),
.A2(n_33),
.B1(n_54),
.B2(n_58),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_9),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_5),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_5),
.A2(n_38),
.B1(n_43),
.B2(n_60),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_60),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_26),
.B1(n_38),
.B2(n_43),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_38),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_7),
.A2(n_46),
.B1(n_54),
.B2(n_58),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_57),
.B(n_70),
.C(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_7),
.A2(n_46),
.B1(n_61),
.B2(n_65),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_7),
.B(n_53),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_7),
.A2(n_58),
.B(n_75),
.C(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_7),
.B(n_24),
.C(n_41),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_7),
.B(n_130),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_7),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_7),
.B(n_44),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_11),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_133),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_131),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_109),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_15),
.B(n_109),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_94),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_81),
.B2(n_82),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_49),
.B2(n_50),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_21),
.B(n_34),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_29),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_22),
.A2(n_93),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_23),
.A2(n_24),
.B1(n_40),
.B2(n_41),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_24),
.B(n_197),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_27),
.B(n_32),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_27),
.B(n_92),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_27),
.A2(n_31),
.B(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_27),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_30),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_30),
.B(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_47),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_35),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_45),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_36),
.B(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_36),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_44),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_37)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_38),
.A2(n_43),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_38),
.B(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_43),
.A2(n_46),
.B(n_76),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_44),
.B(n_153),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_45),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_46),
.A2(n_56),
.B(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_47),
.B(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_71),
.B1(n_72),
.B2(n_80),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_62),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_52),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_54),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_58),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_63),
.Y(n_98)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_77),
.B(n_78),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_73),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_73),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_77),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_79),
.B(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_84),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_84),
.B(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_86),
.B(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_88),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_93),
.B(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_104),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_107),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_115),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_110),
.A2(n_111),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_114),
.Y(n_230)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_125),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_117),
.A2(n_118),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_129),
.B(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_231),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_225),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_163),
.B(n_224),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_154),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_137),
.B(n_154),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.C(n_149),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_138),
.B(n_222),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_139),
.B(n_157),
.C(n_158),
.Y(n_226)
);

FAx1_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.CI(n_143),
.CON(n_139),
.SN(n_139)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_145),
.B(n_149),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_146),
.A2(n_148),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_146),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_148),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_219),
.B(n_223),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_207),
.B(n_218),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_186),
.B(n_206),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_167),
.B(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_170),
.B1(n_171),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_180),
.B2(n_185),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_179),
.C(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_194),
.B(n_205),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_201),
.B(n_204),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);


endmodule