module fake_jpeg_24582_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_27),
.B1(n_25),
.B2(n_16),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_53),
.B1(n_17),
.B2(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_13),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_52),
.Y(n_56)
);

AO22x1_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_16),
.B1(n_27),
.B2(n_28),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_24),
.B(n_22),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_16),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_28),
.B(n_30),
.C(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_37),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_18),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_20),
.B1(n_16),
.B2(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_60),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_43),
.B1(n_22),
.B2(n_39),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_38),
.C(n_32),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_66),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_32),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_67),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_65),
.B(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_30),
.Y(n_67)
);

OAI22x1_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_68),
.A2(n_14),
.B1(n_49),
.B2(n_7),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_54),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_77),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_48),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_69),
.C(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_47),
.B1(n_51),
.B2(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_64),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_47),
.B1(n_51),
.B2(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_87),
.B(n_89),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_96),
.B1(n_77),
.B2(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_56),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_97),
.B(n_78),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_59),
.B1(n_70),
.B2(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_66),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_65),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_104),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_74),
.B(n_64),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_79),
.B(n_83),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_82),
.B1(n_75),
.B2(n_84),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_97),
.C(n_95),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_113),
.C(n_101),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_72),
.C(n_91),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_92),
.C(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_116),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_117),
.C(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_102),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_106),
.A3(n_105),
.B1(n_108),
.B2(n_61),
.C1(n_80),
.C2(n_73),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_73),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_9),
.B(n_10),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_122),
.C(n_11),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_6),
.Y(n_125)
);


endmodule