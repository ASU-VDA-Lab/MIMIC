module real_jpeg_25569_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_244;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_30),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_30),
.B1(n_48),
.B2(n_49),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_2),
.A2(n_30),
.B1(n_54),
.B2(n_55),
.Y(n_180)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_64),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_64),
.Y(n_125)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_7),
.A2(n_9),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_57),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_33),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_9),
.A2(n_33),
.B1(n_54),
.B2(n_55),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_9),
.B(n_22),
.C(n_25),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_21),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_49),
.C(n_61),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_9),
.B(n_51),
.C(n_54),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_9),
.B(n_11),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_9),
.B(n_74),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_9),
.B(n_79),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_11),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_11),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_114),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_113),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_98),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_15),
.B(n_98),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_70),
.C(n_80),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_16),
.A2(n_17),
.B1(n_70),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_18),
.B(n_42),
.C(n_58),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_18),
.A2(n_19),
.B1(n_103),
.B2(n_112),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_18),
.B(n_131),
.C(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_18),
.A2(n_19),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_18),
.A2(n_19),
.B1(n_154),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_19),
.B(n_145),
.C(n_154),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_27),
.B(n_31),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_36),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_21),
.A2(n_32),
.B1(n_36),
.B2(n_109),
.Y(n_108)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_26),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_23),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_23),
.A2(n_25),
.B1(n_60),
.B2(n_61),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_25),
.B(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_35),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_58),
.B2(n_69),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_41),
.A2(n_42),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_56),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_44),
.B(n_93),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_53),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_46),
.A2(n_74),
.B1(n_93),
.B2(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

OA22x2_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_49),
.B(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_73),
.B(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_53),
.A2(n_92),
.B(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_54),
.B(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_65),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_65),
.B(n_78),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_59),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_66),
.B1(n_79),
.B2(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_68),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_68),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_71),
.B(n_76),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_70),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_76),
.A2(n_108),
.B1(n_111),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_76),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_76),
.B(n_193),
.C(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_76),
.A2(n_183),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_76),
.B(n_108),
.C(n_173),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_134),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B(n_94),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_94),
.B1(n_95),
.B2(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_81),
.A2(n_91),
.B1(n_120),
.B2(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_83),
.B(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_89),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_91),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_108),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_123),
.C(n_131),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_111),
.B1(n_131),
.B2(n_132),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_136),
.B(n_275),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_133),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_117),
.B(n_133),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_122),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_121),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_124),
.A2(n_128),
.B1(n_129),
.B2(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_124),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_128),
.A2(n_129),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_128),
.A2(n_129),
.B1(n_206),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_129),
.B(n_200),
.C(n_206),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_129),
.B(n_178),
.C(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_131),
.A2(n_132),
.B1(n_169),
.B2(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_131),
.A2(n_132),
.B1(n_152),
.B2(n_166),
.Y(n_243)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_132),
.B(n_152),
.C(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_159),
.B(n_274),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_157),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_139),
.B(n_157),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_140),
.B(n_142),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_144),
.B(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_145),
.A2(n_146),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_152),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_150),
.A2(n_180),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_152),
.A2(n_166),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_152),
.B(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_154),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_269),
.B(n_273),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_196),
.B(n_255),
.C(n_268),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_185),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_162),
.B(n_185),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_172),
.B2(n_184),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_165),
.B(n_171),
.C(n_184),
.Y(n_256)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_182),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_177),
.A2(n_178),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_229),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.C(n_192),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_187),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_192),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_195),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_193),
.B(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_195),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_254),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_215),
.B(n_253),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_212),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_199),
.B(n_212),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_200),
.A2(n_201),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_205),
.B(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_246),
.B(n_252),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_240),
.B(n_245),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_232),
.B(n_239),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_224),
.B(n_231),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_221),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_228),
.B(n_230),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_234),
.Y(n_239)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_248),
.Y(n_252)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_264),
.B2(n_265),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_265),
.C(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);


endmodule