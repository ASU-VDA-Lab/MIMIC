module fake_jpeg_24229_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_17),
.B1(n_16),
.B2(n_29),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_58),
.Y(n_65)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_33),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_32),
.B(n_31),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_18),
.B1(n_27),
.B2(n_32),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_18),
.B1(n_27),
.B2(n_31),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_31),
.B1(n_22),
.B2(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_22),
.B1(n_25),
.B2(n_28),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_52),
.A3(n_41),
.B1(n_51),
.B2(n_48),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_R g100 ( 
.A(n_63),
.B(n_77),
.Y(n_100)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_28),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_34),
.C(n_49),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_45),
.C(n_50),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_74),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_16),
.B1(n_19),
.B2(n_24),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_69),
.B1(n_67),
.B2(n_70),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_73),
.Y(n_91)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_79),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_15),
.C(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_39),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_50),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_90),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_93),
.B1(n_64),
.B2(n_21),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_20),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_46),
.B1(n_43),
.B2(n_55),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_43),
.B1(n_56),
.B2(n_19),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_40),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_62),
.B(n_20),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_38),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_30),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_45),
.C(n_35),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_40),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_35),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_73),
.B1(n_82),
.B2(n_80),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_118),
.B1(n_125),
.B2(n_92),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_128),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_30),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_123),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_29),
.B1(n_23),
.B2(n_24),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_79),
.B(n_75),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_103),
.B(n_102),
.Y(n_131)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_129),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_127),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_30),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_74),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_108),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_96),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_30),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_99),
.Y(n_135)
);

AOI21x1_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_29),
.B(n_61),
.Y(n_161)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_94),
.B(n_90),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_95),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_95),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_142),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_105),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_2),
.C(n_3),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_107),
.C(n_88),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_149),
.C(n_1),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_30),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_106),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_148),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_86),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_87),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_89),
.B1(n_109),
.B2(n_21),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_142),
.B1(n_131),
.B2(n_146),
.Y(n_163)
);

OAI322xp33_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_117),
.A3(n_113),
.B1(n_127),
.B2(n_126),
.C1(n_121),
.C2(n_123),
.Y(n_151)
);

AOI321xp33_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_144),
.A3(n_134),
.B1(n_133),
.B2(n_7),
.C(n_8),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_117),
.B1(n_111),
.B2(n_114),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_150),
.B1(n_134),
.B2(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_162),
.C(n_164),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_165),
.C(n_146),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_145),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_2),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_3),
.C(n_4),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_136),
.Y(n_167)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_132),
.C(n_141),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_175),
.C(n_176),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_173),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_160),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_4),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_4),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_164),
.C(n_152),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_183),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_159),
.B(n_157),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_8),
.B(n_10),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_158),
.C(n_163),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_170),
.C(n_176),
.Y(n_187)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_5),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_191),
.C(n_179),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_157),
.B1(n_172),
.B2(n_158),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_10),
.C(n_12),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_166),
.B1(n_170),
.B2(n_7),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_189),
.A2(n_192),
.B1(n_14),
.B2(n_11),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_181),
.B(n_11),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_189),
.Y(n_200)
);

AOI21x1_ASAP7_75t_SL g201 ( 
.A1(n_195),
.A2(n_197),
.B(n_13),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_186),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_196),
.A2(n_190),
.B(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_198),
.B(n_13),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_200),
.C(n_196),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_13),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_203),
.Y(n_206)
);


endmodule