module real_jpeg_4997_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_1),
.A2(n_83),
.B1(n_85),
.B2(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_1),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_1),
.A2(n_55),
.B1(n_88),
.B2(n_224),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_1),
.A2(n_88),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_1),
.A2(n_88),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_2),
.Y(n_150)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_2),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_3),
.A2(n_167),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_54),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_4),
.A2(n_54),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_4),
.A2(n_54),
.B1(n_258),
.B2(n_261),
.Y(n_257)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_6),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_6),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_6),
.Y(n_189)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_6),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_6),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_7),
.A2(n_85),
.B1(n_91),
.B2(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_7),
.A2(n_95),
.B1(n_209),
.B2(n_253),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_7),
.A2(n_95),
.B1(n_308),
.B2(n_310),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_8),
.A2(n_46),
.B1(n_110),
.B2(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_8),
.B(n_98),
.C(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_8),
.B(n_74),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_8),
.B(n_162),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_8),
.B(n_197),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_8),
.B(n_83),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_9),
.Y(n_140)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_11),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_12),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_12),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_12),
.A2(n_115),
.B1(n_173),
.B2(n_187),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_13),
.A2(n_153),
.B1(n_158),
.B2(n_161),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_13),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_13),
.A2(n_161),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_14),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_14),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_15),
.A2(n_102),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_15),
.Y(n_208)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_233),
.B1(n_234),
.B2(n_350),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_18),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_232),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_191),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_20),
.B(n_191),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_129),
.C(n_175),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_21),
.B(n_347),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_61),
.B2(n_128),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_22),
.B(n_62),
.C(n_96),
.Y(n_215)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_51),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_24),
.B(n_53),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_33),
.B(n_46),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_33)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_34),
.A2(n_47),
.A3(n_133),
.B1(n_136),
.B2(n_138),
.Y(n_132)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_38),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_38),
.Y(n_183)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_47),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_46),
.A2(n_145),
.B(n_255),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_SL g314 ( 
.A1(n_46),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_60),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_60),
.Y(n_226)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_96),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g184 ( 
.A(n_63),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_74),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_64)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_65),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_68),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_73),
.Y(n_315)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_74)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_76),
.Y(n_201)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_78),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_78),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_78),
.Y(n_268)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_82),
.A2(n_89),
.B(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_89),
.B(n_179),
.Y(n_231)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_94),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_109),
.B(n_116),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_97),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_97),
.A2(n_116),
.B(n_265),
.Y(n_264)
);

AOI22x1_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_104),
.B2(n_106),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_103),
.Y(n_261)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_109),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_114),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_117),
.B(n_197),
.Y(n_244)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_119),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_123),
.B1(n_125),
.B2(n_127),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_121),
.Y(n_195)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_127),
.Y(n_247)
);

INVx5_ASAP7_75t_SL g311 ( 
.A(n_127),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_129),
.A2(n_130),
.B1(n_175),
.B2(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_143),
.B2(n_144),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_132),
.B(n_143),
.Y(n_219)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_151),
.B1(n_162),
.B2(n_165),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_145),
.A2(n_252),
.B(n_255),
.Y(n_251)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_152),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_146),
.A2(n_166),
.B1(n_206),
.B2(n_211),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_146),
.B(n_257),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_146),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_147),
.Y(n_256)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_160),
.Y(n_254)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_174),
.Y(n_285)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_175),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_185),
.C(n_190),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_176),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_184),
.A2(n_231),
.B(n_314),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_185),
.B(n_190),
.Y(n_341)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_186),
.Y(n_320)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_218),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_205),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_195),
.A2(n_241),
.B(n_244),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_195),
.A2(n_196),
.B1(n_265),
.B2(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_195),
.A2(n_244),
.B(n_307),
.Y(n_338)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_SL g325 ( 
.A(n_201),
.Y(n_325)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_210),
.Y(n_283)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_228),
.B2(n_229),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_226),
.B(n_227),
.Y(n_222)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_344),
.B(n_349),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_333),
.B(n_343),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_301),
.B(n_332),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_271),
.B(n_300),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_250),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_250),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_240),
.A2(n_245),
.B1(n_246),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_240),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g330 ( 
.A(n_242),
.B(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_262),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_263),
.C(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_252),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_269),
.B2(n_270),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_291),
.B(n_299),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_278),
.B(n_290),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_289),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_289),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_286),
.B(n_288),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_297),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_303),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_318),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_312),
.B2(n_313),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_312),
.C(n_318),
.Y(n_334)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI32xp33_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_323),
.A3(n_325),
.B1(n_326),
.B2(n_330),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_322),
.Y(n_339)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_334),
.B(n_335),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_340),
.B2(n_342),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_339),
.C(n_342),
.Y(n_345)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_345),
.B(n_346),
.Y(n_349)
);


endmodule