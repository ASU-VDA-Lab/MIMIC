module real_aes_4601_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_87;
wire n_171;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g351 ( .A(n_0), .B(n_283), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_1), .A2(n_20), .B1(n_178), .B2(n_183), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_2), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_SL g287 ( .A1(n_3), .A2(n_249), .B(n_288), .C(n_290), .Y(n_287) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_4), .A2(n_65), .B1(n_248), .B2(n_254), .Y(n_356) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_5), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_6), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_7), .A2(n_55), .B1(n_252), .B2(n_254), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_8), .Y(n_84) );
INVx1_ASAP7_75t_L g117 ( .A(n_9), .Y(n_117) );
INVxp67_ASAP7_75t_L g130 ( .A(n_9), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_9), .B(n_58), .Y(n_137) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_10), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_11), .A2(n_46), .B1(n_246), .B2(n_248), .Y(n_245) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_11), .Y(n_637) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_12), .A2(n_56), .B(n_262), .Y(n_261) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_12), .A2(n_56), .B(n_262), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_13), .B(n_102), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_14), .A2(n_30), .B1(n_194), .B2(n_197), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_15), .Y(n_380) );
BUFx3_ASAP7_75t_L g221 ( .A(n_16), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g294 ( .A1(n_17), .A2(n_295), .B(n_296), .C(n_298), .Y(n_294) );
OAI22xp33_ASAP7_75t_SL g354 ( .A1(n_18), .A2(n_33), .B1(n_248), .B2(n_274), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_19), .A2(n_25), .B1(n_274), .B2(n_278), .Y(n_343) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_21), .Y(n_102) );
O2A1O1Ixp5_ASAP7_75t_L g310 ( .A1(n_22), .A2(n_249), .B(n_311), .C(n_313), .Y(n_310) );
AO22x1_ASAP7_75t_L g120 ( .A1(n_23), .A2(n_54), .B1(n_121), .B2(n_132), .Y(n_120) );
INVx1_ASAP7_75t_L g103 ( .A(n_24), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_24), .B(n_57), .Y(n_127) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_26), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_27), .A2(n_68), .B1(n_146), .B2(n_151), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_28), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_29), .B(n_328), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_31), .Y(n_292) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_32), .Y(n_210) );
INVx1_ASAP7_75t_L g262 ( .A(n_34), .Y(n_262) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_35), .Y(n_232) );
AND2x4_ASAP7_75t_L g258 ( .A(n_35), .B(n_230), .Y(n_258) );
AND2x4_ASAP7_75t_L g301 ( .A(n_35), .B(n_230), .Y(n_301) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_36), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g92 ( .A1(n_37), .A2(n_93), .B(n_120), .Y(n_92) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_38), .A2(n_45), .B1(n_188), .B2(n_190), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_39), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_40), .Y(n_320) );
INVx2_ASAP7_75t_L g279 ( .A(n_41), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g381 ( .A1(n_42), .A2(n_249), .B(n_382), .C(n_383), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_43), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g156 ( .A1(n_44), .A2(n_53), .B1(n_157), .B2(n_161), .Y(n_156) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_46), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_47), .A2(n_62), .B1(n_289), .B2(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_48), .B(n_259), .Y(n_367) );
OA22x2_ASAP7_75t_L g107 ( .A1(n_49), .A2(n_58), .B1(n_102), .B2(n_106), .Y(n_107) );
INVx1_ASAP7_75t_L g144 ( .A(n_49), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_50), .Y(n_366) );
NAND2xp33_ASAP7_75t_R g263 ( .A(n_51), .B(n_264), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_51), .A2(n_77), .B1(n_328), .B2(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_52), .A2(n_69), .B1(n_166), .B2(n_174), .Y(n_165) );
INVx1_ASAP7_75t_L g119 ( .A(n_57), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_57), .B(n_141), .Y(n_140) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_57), .Y(n_224) );
OAI21xp33_ASAP7_75t_L g155 ( .A1(n_58), .A2(n_64), .B(n_131), .Y(n_155) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_59), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_60), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_61), .Y(n_275) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_63), .A2(n_88), .B1(n_89), .B2(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_63), .Y(n_629) );
INVx1_ASAP7_75t_L g105 ( .A(n_64), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_64), .B(n_74), .Y(n_138) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_66), .Y(n_247) );
BUFx5_ASAP7_75t_L g248 ( .A(n_66), .Y(n_248) );
INVx1_ASAP7_75t_L g253 ( .A(n_66), .Y(n_253) );
INVx2_ASAP7_75t_L g303 ( .A(n_67), .Y(n_303) );
INVx2_ASAP7_75t_L g386 ( .A(n_70), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_71), .Y(n_297) );
INVx2_ASAP7_75t_SL g230 ( .A(n_72), .Y(n_230) );
INVx1_ASAP7_75t_L g318 ( .A(n_73), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_74), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g323 ( .A(n_75), .Y(n_323) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_76), .Y(n_85) );
OAI21xp33_ASAP7_75t_SL g378 ( .A1(n_76), .A2(n_248), .B(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_SL g281 ( .A(n_77), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_77), .B(n_328), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_216), .B1(n_233), .B2(n_615), .C(n_622), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_201), .Y(n_79) );
AOI22xp33_ASAP7_75t_SL g80 ( .A1(n_81), .A2(n_82), .B1(n_88), .B2(n_89), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_82) );
INVx1_ASAP7_75t_L g86 ( .A(n_83), .Y(n_86) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_84), .A2(n_248), .B1(n_274), .B2(n_275), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_85), .Y(n_87) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_88), .A2(n_89), .B1(n_624), .B2(n_625), .Y(n_623) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
NOR2x1_ASAP7_75t_L g90 ( .A(n_91), .B(n_164), .Y(n_90) );
NAND3xp33_ASAP7_75t_L g91 ( .A(n_92), .B(n_145), .C(n_156), .Y(n_91) );
INVx2_ASAP7_75t_SL g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_108), .Y(n_98) );
AND2x2_ASAP7_75t_L g163 ( .A(n_99), .B(n_160), .Y(n_163) );
AND2x2_ASAP7_75t_L g180 ( .A(n_99), .B(n_181), .Y(n_180) );
AND2x4_ASAP7_75t_L g185 ( .A(n_99), .B(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g99 ( .A(n_100), .B(n_107), .Y(n_99) );
INVx1_ASAP7_75t_L g150 ( .A(n_100), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_101), .B(n_104), .Y(n_100) );
NAND2xp33_ASAP7_75t_L g101 ( .A(n_102), .B(n_103), .Y(n_101) );
INVx2_ASAP7_75t_L g106 ( .A(n_102), .Y(n_106) );
INVx3_ASAP7_75t_L g112 ( .A(n_102), .Y(n_112) );
NAND2xp33_ASAP7_75t_L g118 ( .A(n_102), .B(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_102), .Y(n_126) );
INVx1_ASAP7_75t_L g131 ( .A(n_102), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_103), .B(n_144), .Y(n_143) );
INVxp67_ASAP7_75t_L g225 ( .A(n_103), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OAI21xp5_ASAP7_75t_L g129 ( .A1(n_105), .A2(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_L g128 ( .A(n_107), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g149 ( .A(n_107), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g170 ( .A(n_107), .Y(n_170) );
AND2x4_ASAP7_75t_L g148 ( .A(n_108), .B(n_149), .Y(n_148) );
AND2x4_ASAP7_75t_L g153 ( .A(n_108), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g192 ( .A(n_108), .B(n_169), .Y(n_192) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_114), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g124 ( .A(n_110), .B(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g160 ( .A(n_110), .B(n_114), .Y(n_160) );
OR2x2_ASAP7_75t_L g172 ( .A(n_110), .B(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g181 ( .A(n_110), .B(n_182), .Y(n_181) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_112), .B(n_117), .Y(n_116) );
INVxp67_ASAP7_75t_L g141 ( .A(n_112), .Y(n_141) );
NAND3xp33_ASAP7_75t_L g139 ( .A(n_113), .B(n_140), .C(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g173 ( .A(n_115), .Y(n_173) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_118), .Y(n_115) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx5_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_128), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g135 ( .A(n_126), .Y(n_135) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_127), .Y(n_222) );
INVx2_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_139), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_141), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g154 ( .A(n_142), .B(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_144), .Y(n_226) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g159 ( .A(n_149), .B(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g169 ( .A(n_150), .B(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g176 ( .A(n_154), .B(n_171), .Y(n_176) );
AND2x4_ASAP7_75t_L g200 ( .A(n_154), .B(n_181), .Y(n_200) );
BUFx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g189 ( .A(n_160), .B(n_169), .Y(n_189) );
BUFx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND4xp25_ASAP7_75t_SL g164 ( .A(n_165), .B(n_177), .C(n_187), .D(n_193), .Y(n_164) );
BUFx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_171), .Y(n_168) );
AND2x4_ASAP7_75t_L g196 ( .A(n_169), .B(n_181), .Y(n_196) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g186 ( .A(n_172), .Y(n_186) );
INVx1_ASAP7_75t_L g182 ( .A(n_173), .Y(n_182) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
BUFx12f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx12f_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx12f_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx5_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx8_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B1(n_214), .B2(n_215), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_202), .Y(n_214) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_203), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B1(n_212), .B2(n_213), .Y(n_203) );
INVx1_ASAP7_75t_L g212 ( .A(n_204), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_205), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B1(n_208), .B2(n_211), .Y(n_205) );
CKINVDCx16_ASAP7_75t_R g211 ( .A(n_206), .Y(n_211) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
XOR2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
BUFx10_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_227), .Y(n_218) );
INVxp67_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g627 ( .A(n_220), .B(n_227), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .C(n_226), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_231), .Y(n_227) );
OR2x2_ASAP7_75t_L g631 ( .A(n_228), .B(n_232), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_228), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_228), .B(n_231), .Y(n_635) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_235), .B(n_512), .Y(n_234) );
NOR3xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_423), .C(n_471), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_368), .Y(n_236) );
OAI21xp33_ASAP7_75t_SL g237 ( .A1(n_238), .A2(n_304), .B(n_335), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_238), .A2(n_583), .B(n_585), .Y(n_582) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_265), .Y(n_239) );
OR2x2_ASAP7_75t_L g510 ( .A(n_240), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_240), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g391 ( .A(n_242), .Y(n_391) );
INVx2_ASAP7_75t_L g422 ( .A(n_242), .Y(n_422) );
AND2x2_ASAP7_75t_L g443 ( .A(n_242), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g562 ( .A(n_242), .B(n_267), .Y(n_562) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_263), .Y(n_242) );
AND2x2_ASAP7_75t_L g463 ( .A(n_243), .B(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_256), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_249), .B1(n_251), .B2(n_255), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_246), .A2(n_277), .B1(n_278), .B2(n_279), .Y(n_276) );
INVx1_ASAP7_75t_L g295 ( .A(n_246), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_246), .A2(n_248), .B1(n_365), .B2(n_366), .Y(n_364) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g254 ( .A(n_247), .Y(n_254) );
INVx6_ASAP7_75t_L g274 ( .A(n_247), .Y(n_274) );
INVx3_ASAP7_75t_L g312 ( .A(n_247), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_248), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_248), .B(n_320), .Y(n_319) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_248), .A2(n_274), .B1(n_362), .B2(n_363), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_248), .B(n_380), .Y(n_379) );
OAI22xp33_ASAP7_75t_L g272 ( .A1(n_249), .A2(n_255), .B1(n_273), .B2(n_276), .Y(n_272) );
INVx1_ASAP7_75t_L g334 ( .A(n_249), .Y(n_334) );
OAI221xp5_ASAP7_75t_L g360 ( .A1(n_249), .A2(n_258), .B1(n_298), .B2(n_361), .C(n_364), .Y(n_360) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx4_ASAP7_75t_L g255 ( .A(n_250), .Y(n_255) );
INVx3_ASAP7_75t_L g298 ( .A(n_250), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_250), .B(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_250), .Y(n_342) );
INVx1_ASAP7_75t_L g346 ( .A(n_250), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_250), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g289 ( .A(n_252), .Y(n_289) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g278 ( .A(n_253), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_255), .A2(n_316), .B1(n_317), .B2(n_319), .Y(n_315) );
INVx2_ASAP7_75t_L g331 ( .A(n_255), .Y(n_331) );
NOR2xp67_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_258), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_258), .B(n_284), .Y(n_357) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
BUFx3_ASAP7_75t_L g321 ( .A(n_260), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_260), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx4_ASAP7_75t_L g284 ( .A(n_261), .Y(n_284) );
BUFx3_ASAP7_75t_L g409 ( .A(n_261), .Y(n_409) );
BUFx3_ASAP7_75t_L g271 ( .A(n_264), .Y(n_271) );
INVx1_ASAP7_75t_L g324 ( .A(n_264), .Y(n_324) );
INVx1_ASAP7_75t_L g376 ( .A(n_264), .Y(n_376) );
INVx2_ASAP7_75t_L g466 ( .A(n_264), .Y(n_466) );
INVx2_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_266), .B(n_395), .Y(n_515) );
AND2x2_ASAP7_75t_L g602 ( .A(n_266), .B(n_546), .Y(n_602) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_285), .Y(n_266) );
INVx1_ASAP7_75t_L g419 ( .A(n_267), .Y(n_419) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_272), .B(n_280), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x2_ASAP7_75t_L g616 ( .A(n_269), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_270), .B(n_301), .Y(n_340) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g332 ( .A(n_273), .Y(n_332) );
INVx2_ASAP7_75t_L g291 ( .A(n_274), .Y(n_291) );
INVx2_ASAP7_75t_SL g345 ( .A(n_274), .Y(n_345) );
INVx1_ASAP7_75t_L g333 ( .A(n_276), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_278), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_278), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g359 ( .A(n_282), .Y(n_359) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_SL g299 ( .A(n_283), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_SL g302 ( .A(n_284), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g328 ( .A(n_284), .Y(n_328) );
OR2x2_ASAP7_75t_L g325 ( .A(n_285), .B(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_285), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_285), .B(n_308), .Y(n_400) );
INVx2_ASAP7_75t_L g421 ( .A(n_285), .Y(n_421) );
INVx1_ASAP7_75t_L g460 ( .A(n_285), .Y(n_460) );
INVx1_ASAP7_75t_L g501 ( .A(n_285), .Y(n_501) );
AND2x2_ASAP7_75t_L g536 ( .A(n_285), .B(n_326), .Y(n_536) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_285), .Y(n_591) );
AO31x2_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_293), .A3(n_299), .B(n_302), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_295), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_298), .A2(n_356), .B(n_357), .Y(n_355) );
NOR3xp33_ASAP7_75t_L g309 ( .A(n_300), .B(n_310), .C(n_315), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_300), .A2(n_331), .B1(n_332), .B2(n_333), .C(n_334), .Y(n_330) );
INVx4_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g375 ( .A(n_301), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_325), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g390 ( .A(n_308), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g429 ( .A(n_308), .B(n_421), .Y(n_429) );
INVx2_ASAP7_75t_L g444 ( .A(n_308), .Y(n_444) );
INVx2_ASAP7_75t_L g470 ( .A(n_308), .Y(n_470) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_321), .B(n_322), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g316 ( .A(n_312), .Y(n_316) );
INVx1_ASAP7_75t_L g382 ( .A(n_312), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_321), .B(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_325), .Y(n_426) );
OR2x2_ASAP7_75t_L g441 ( .A(n_325), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g518 ( .A(n_325), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_326), .B(n_470), .Y(n_469) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_326), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_326), .B(n_526), .Y(n_552) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g462 ( .A(n_329), .B(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_331), .A2(n_378), .B(n_381), .Y(n_377) );
AOI322xp5_ASAP7_75t_L g544 ( .A1(n_335), .A2(n_484), .A3(n_522), .B1(n_545), .B2(n_547), .C1(n_548), .C2(n_549), .Y(n_544) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_348), .Y(n_335) );
AND2x2_ASAP7_75t_L g549 ( .A(n_336), .B(n_529), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_336), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g600 ( .A(n_336), .B(n_492), .Y(n_600) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_337), .B(n_397), .Y(n_415) );
AND2x2_ASAP7_75t_L g476 ( .A(n_337), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_337), .B(n_438), .Y(n_520) );
AND2x4_ASAP7_75t_L g557 ( .A(n_337), .B(n_348), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_337), .B(n_479), .Y(n_598) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g387 ( .A(n_338), .B(n_358), .Y(n_387) );
INVx1_ASAP7_75t_L g436 ( .A(n_338), .Y(n_436) );
AND2x2_ASAP7_75t_L g580 ( .A(n_338), .B(n_413), .Y(n_580) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g398 ( .A(n_339), .Y(n_398) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B(n_347), .Y(n_339) );
INVx1_ASAP7_75t_L g407 ( .A(n_341), .Y(n_407) );
OA22x2_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_344), .B2(n_346), .Y(n_341) );
INVx4_ASAP7_75t_L g621 ( .A(n_342), .Y(n_621) );
INVx1_ASAP7_75t_L g410 ( .A(n_347), .Y(n_410) );
INVx1_ASAP7_75t_SL g505 ( .A(n_348), .Y(n_505) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_358), .Y(n_348) );
AND2x2_ASAP7_75t_L g397 ( .A(n_349), .B(n_373), .Y(n_397) );
INVx1_ASAP7_75t_L g438 ( .A(n_349), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_349), .B(n_372), .Y(n_614) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g413 ( .A(n_350), .Y(n_413) );
INVx1_ASAP7_75t_L g455 ( .A(n_350), .Y(n_455) );
AND2x2_ASAP7_75t_L g479 ( .A(n_350), .B(n_358), .Y(n_479) );
AND2x2_ASAP7_75t_L g529 ( .A(n_350), .B(n_373), .Y(n_529) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_350), .Y(n_533) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
OR2x2_ASAP7_75t_L g405 ( .A(n_358), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g435 ( .A(n_358), .B(n_436), .Y(n_435) );
OA21x2_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B(n_367), .Y(n_358) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_359), .A2(n_360), .B(n_367), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_388), .B1(n_395), .B2(n_399), .C(n_401), .Y(n_368) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_387), .Y(n_370) );
AND2x2_ASAP7_75t_L g575 ( .A(n_371), .B(n_435), .Y(n_575) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g589 ( .A(n_372), .B(n_470), .Y(n_589) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g412 ( .A(n_373), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g433 ( .A(n_373), .Y(n_433) );
AND2x2_ASAP7_75t_L g456 ( .A(n_373), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g478 ( .A(n_373), .Y(n_478) );
BUFx2_ASAP7_75t_L g566 ( .A(n_373), .Y(n_566) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI21x1_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_385), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_387), .A2(n_411), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g578 ( .A(n_387), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_388), .A2(n_425), .B1(n_430), .B2(n_437), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
OR2x2_ASAP7_75t_L g486 ( .A(n_389), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g517 ( .A(n_390), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g535 ( .A(n_390), .B(n_536), .Y(n_535) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g609 ( .A(n_394), .B(n_525), .Y(n_609) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR2xp33_ASAP7_75t_SL g521 ( .A(n_396), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x2_ASAP7_75t_L g497 ( .A(n_398), .B(n_478), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_398), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g584 ( .A(n_398), .Y(n_584) );
OR2x2_ASAP7_75t_L g613 ( .A(n_398), .B(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g581 ( .A(n_399), .B(n_562), .Y(n_581) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_414), .B(n_416), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_411), .Y(n_403) );
AND2x2_ASAP7_75t_L g437 ( .A(n_404), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g539 ( .A(n_404), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g448 ( .A(n_406), .B(n_449), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_410), .Y(n_406) );
INVx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g492 ( .A(n_413), .B(n_449), .Y(n_492) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_414), .A2(n_499), .B(n_611), .Y(n_610) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g592 ( .A(n_418), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g467 ( .A(n_420), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g551 ( .A(n_420), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g488 ( .A(n_421), .Y(n_488) );
INVx1_ASAP7_75t_L g527 ( .A(n_422), .Y(n_527) );
AND2x4_ASAP7_75t_L g546 ( .A(n_422), .B(n_470), .Y(n_546) );
INVx1_ASAP7_75t_SL g593 ( .A(n_422), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_439), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g561 ( .A(n_429), .B(n_562), .Y(n_561) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g446 ( .A(n_432), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g545 ( .A(n_432), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_433), .B(n_457), .Y(n_607) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_437), .B(n_458), .Y(n_493) );
AND2x2_ASAP7_75t_L g484 ( .A(n_438), .B(n_448), .Y(n_484) );
AOI222xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_445), .B1(n_451), .B2(n_453), .C1(n_458), .C2(n_467), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g490 ( .A1(n_441), .A2(n_491), .B(n_493), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g558 ( .A1(n_441), .A2(n_559), .B1(n_560), .B2(n_563), .C(n_567), .Y(n_558) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx2_ASAP7_75t_L g473 ( .A(n_443), .Y(n_473) );
AND2x2_ASAP7_75t_L g502 ( .A(n_444), .B(n_462), .Y(n_502) );
INVx1_ASAP7_75t_L g526 ( .A(n_444), .Y(n_526) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_444), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_445), .A2(n_539), .B(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g569 ( .A(n_448), .B(n_540), .Y(n_569) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g457 ( .A(n_450), .Y(n_457) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_456), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_456), .Y(n_483) );
INVx2_ASAP7_75t_L g534 ( .A(n_457), .Y(n_534) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
OR2x2_ASAP7_75t_L g590 ( .A(n_461), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g556 ( .A(n_462), .Y(n_556) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_467), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g511 ( .A(n_469), .B(n_488), .Y(n_511) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_480), .C(n_489), .D(n_494), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_473), .A2(n_568), .B(n_569), .C(n_570), .Y(n_567) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g508 ( .A(n_478), .Y(n_508) );
INVx1_ASAP7_75t_L g540 ( .A(n_478), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_484), .B(n_485), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVxp33_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_492), .B(n_566), .Y(n_571) );
AND2x4_ASAP7_75t_L g583 ( .A(n_492), .B(n_584), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g594 ( .A(n_492), .B(n_507), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B1(n_503), .B2(n_509), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2x1p5_ASAP7_75t_SL g499 ( .A(n_500), .B(n_502), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g568 ( .A(n_501), .Y(n_568) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_502), .Y(n_548) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
OR2x2_ASAP7_75t_L g559 ( .A(n_506), .B(n_532), .Y(n_559) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g547 ( .A(n_511), .Y(n_547) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_572), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_537), .C(n_558), .Y(n_513) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .C(n_528), .Y(n_514) );
AOI22x1_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_519), .B1(n_521), .B2(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
OAI21xp33_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_530), .B(n_535), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .Y(n_530) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVxp67_ASAP7_75t_L g606 ( .A(n_533), .Y(n_606) );
INVx1_ASAP7_75t_L g586 ( .A(n_534), .Y(n_586) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_536), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_544), .C(n_550), .Y(n_537) );
INVx1_ASAP7_75t_L g579 ( .A(n_540), .Y(n_579) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_553), .B(n_557), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_551), .A2(n_569), .B1(n_604), .B2(n_608), .Y(n_603) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVxp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_595), .C(n_610), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_582), .Y(n_573) );
OAI31xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .A3(n_580), .B(n_581), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_592), .B2(n_594), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_599), .B(n_601), .C(n_603), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OA21x2_ASAP7_75t_L g633 ( .A1(n_617), .A2(n_634), .B(n_635), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
CKINVDCx16_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI222xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B1(n_628), .B2(n_630), .C1(n_632), .C2(n_636), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_624), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
endmodule