module fake_jpeg_8045_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_44),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_16),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_23),
.B1(n_30),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_29),
.B1(n_33),
.B2(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_61),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_31),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_0),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_68),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_86),
.Y(n_106)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_98),
.B1(n_58),
.B2(n_67),
.Y(n_111)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_78),
.A2(n_90),
.B1(n_28),
.B2(n_64),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_41),
.B1(n_42),
.B2(n_46),
.Y(n_81)
);

AOI211xp5_ASAP7_75t_SL g120 ( 
.A1(n_81),
.A2(n_57),
.B(n_61),
.C(n_59),
.Y(n_120)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_90),
.Y(n_123)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_0),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_88),
.C(n_73),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_99),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_97),
.Y(n_124)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_74),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_104),
.B(n_128),
.Y(n_154)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_115),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_58),
.B1(n_63),
.B2(n_51),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_53),
.B1(n_18),
.B2(n_82),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

OR2x6_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_59),
.Y(n_112)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_113),
.B(n_120),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_30),
.B1(n_55),
.B2(n_50),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_122),
.B1(n_97),
.B2(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_55),
.B1(n_51),
.B2(n_53),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_69),
.B1(n_28),
.B2(n_96),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_92),
.B(n_41),
.CI(n_42),
.CON(n_128),
.SN(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_129),
.A2(n_144),
.B(n_22),
.C(n_34),
.Y(n_189)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_133),
.B(n_136),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_137),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_120),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_92),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_72),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_151),
.C(n_22),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_142),
.B(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_125),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_55),
.B(n_81),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_81),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_81),
.B1(n_75),
.B2(n_76),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_88),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_147),
.B(n_152),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_100),
.B1(n_121),
.B2(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_32),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_156),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_39),
.C(n_93),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_20),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_102),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_173),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_166),
.A2(n_167),
.B1(n_189),
.B2(n_2),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_100),
.B1(n_107),
.B2(n_110),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_143),
.B1(n_150),
.B2(n_142),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_172),
.B1(n_175),
.B2(n_178),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_107),
.B1(n_117),
.B2(n_118),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_1),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_22),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_179),
.C(n_182),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_117),
.B1(n_80),
.B2(n_71),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_20),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_5),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_91),
.B1(n_32),
.B2(n_20),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_32),
.B1(n_21),
.B2(n_36),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_184),
.B1(n_188),
.B2(n_3),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_34),
.C(n_22),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_34),
.B(n_22),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_186),
.B(n_4),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_21),
.B1(n_36),
.B2(n_34),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_136),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_12),
.C(n_14),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_34),
.B(n_21),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_140),
.A2(n_157),
.B1(n_141),
.B2(n_155),
.Y(n_188)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_198),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_11),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_194),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_131),
.B1(n_17),
.B2(n_145),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_1),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_197),
.B(n_200),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_1),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_138),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_199),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_202),
.A2(n_186),
.B1(n_183),
.B2(n_173),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_16),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_206),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_204),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_205),
.B(n_208),
.Y(n_234)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_213),
.B1(n_193),
.B2(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_210),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_165),
.B(n_10),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_5),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_6),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_212),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_165),
.B(n_179),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_218),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_161),
.B(n_10),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_166),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_219),
.B(n_220),
.Y(n_241)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_160),
.C(n_176),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_191),
.B(n_171),
.CI(n_162),
.CON(n_224),
.SN(n_224)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_169),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_193),
.A2(n_171),
.B1(n_169),
.B2(n_178),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_238),
.B1(n_247),
.B2(n_202),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_173),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_190),
.B1(n_158),
.B2(n_177),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_174),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_177),
.B1(n_181),
.B2(n_184),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_214),
.C(n_221),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_249),
.C(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_227),
.B1(n_236),
.B2(n_237),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_261),
.B1(n_226),
.B2(n_234),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_243),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_196),
.C(n_182),
.Y(n_258)
);

XOR2x2_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_235),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_229),
.B(n_235),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_241),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_263),
.C(n_269),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_227),
.A2(n_207),
.B1(n_194),
.B2(n_200),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_208),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_196),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_223),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_197),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_195),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_200),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_265),
.A2(n_230),
.B1(n_247),
.B2(n_234),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_250),
.B1(n_266),
.B2(n_252),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_228),
.C(n_244),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_285),
.C(n_258),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_237),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_284),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_269),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_225),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_238),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_259),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_263),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_272),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_286),
.C(n_280),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_292),
.B(n_302),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_251),
.B(n_256),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_293),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_294),
.B(n_285),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_273),
.A2(n_254),
.B1(n_261),
.B2(n_246),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_298),
.B1(n_277),
.B2(n_270),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_236),
.B1(n_232),
.B2(n_206),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_SL g300 ( 
.A(n_283),
.B(n_200),
.C(n_239),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_SL g301 ( 
.A(n_279),
.B(n_282),
.C(n_274),
.Y(n_301)
);

NAND4xp25_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_232),
.C(n_204),
.D(n_257),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_306),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_304),
.A2(n_288),
.B1(n_296),
.B2(n_301),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_272),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_271),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_309),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_271),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_313),
.B(n_295),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_284),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_299),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_239),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_15),
.Y(n_330)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_13),
.C(n_14),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_310),
.A2(n_300),
.B1(n_295),
.B2(n_292),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_321),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_320),
.B(n_324),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_314),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_13),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_322),
.A2(n_312),
.B1(n_313),
.B2(n_304),
.Y(n_326)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_303),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_327),
.A2(n_329),
.B(n_331),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_330),
.B(n_13),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

AOI322xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_325),
.A3(n_334),
.B1(n_331),
.B2(n_330),
.C1(n_333),
.C2(n_328),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_323),
.C(n_318),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

AOI221xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_7),
.B(n_9),
.Y(n_341)
);


endmodule