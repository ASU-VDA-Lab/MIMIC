module fake_jpeg_12467_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_44),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_17),
.A2(n_25),
.B(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_5),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g70 ( 
.A(n_15),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_24),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_77),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_1),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_82),
.Y(n_88)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g84 ( 
.A(n_76),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_61),
.B1(n_71),
.B2(n_53),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_91),
.B1(n_49),
.B2(n_52),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_58),
.B1(n_57),
.B2(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_61),
.B1(n_49),
.B2(n_71),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_94),
.B1(n_70),
.B2(n_59),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_65),
.Y(n_96)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_105),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_86),
.B1(n_92),
.B2(n_87),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_110),
.Y(n_117)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_18),
.B(n_40),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_50),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_7),
.Y(n_132)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_56),
.B1(n_62),
.B2(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_46),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_67),
.B1(n_60),
.B2(n_54),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_48),
.B1(n_70),
.B2(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_2),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_4),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_4),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_21),
.C(n_41),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_130),
.B(n_9),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_8),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_139),
.A2(n_143),
.B(n_128),
.C(n_116),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_38),
.C(n_42),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_140),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

AOI321xp33_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_153),
.A3(n_154),
.B1(n_147),
.B2(n_136),
.C(n_134),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_149),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_155),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_141),
.B(n_138),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_161),
.Y(n_162)
);


endmodule