module fake_jpeg_26283_n_66 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_66);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_66;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx6p67_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_37),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

AND2x4_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NOR2xp67_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_14),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_13),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_59)
);

BUFx24_ASAP7_75t_SL g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_40),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_16),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B(n_42),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_49),
.C(n_55),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_58),
.C(n_54),
.Y(n_64)
);

AOI31xp33_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_58),
.A3(n_57),
.B(n_56),
.Y(n_65)
);

FAx1_ASAP7_75t_SL g66 ( 
.A(n_65),
.B(n_41),
.CI(n_52),
.CON(n_66),
.SN(n_66)
);


endmodule