module real_aes_4224_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_393;
wire n_84;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx1_ASAP7_75t_L g427 ( .A(n_0), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_1), .A2(n_12), .B1(n_252), .B2(n_382), .Y(n_390) );
INVx2_ASAP7_75t_L g363 ( .A(n_2), .Y(n_363) );
INVx1_ASAP7_75t_SL g336 ( .A(n_3), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_4), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_5), .B(n_285), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_6), .A2(n_70), .B1(n_130), .B2(n_138), .Y(n_129) );
INVx1_ASAP7_75t_L g109 ( .A(n_7), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_7), .B(n_56), .Y(n_181) );
INVxp67_ASAP7_75t_L g209 ( .A(n_7), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_8), .A2(n_23), .B1(n_142), .B2(n_144), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_9), .A2(n_41), .B1(n_274), .B2(n_276), .Y(n_273) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_10), .A2(n_54), .B(n_283), .Y(n_282) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_10), .A2(n_54), .B(n_283), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_11), .B(n_94), .Y(n_105) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_12), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_13), .B(n_319), .Y(n_402) );
INVx1_ASAP7_75t_SL g186 ( .A(n_14), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_15), .A2(n_64), .B1(n_356), .B2(n_357), .Y(n_355) );
INVx2_ASAP7_75t_L g386 ( .A(n_16), .Y(n_386) );
INVx1_ASAP7_75t_L g191 ( .A(n_17), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_18), .A2(n_20), .B1(n_316), .B2(n_335), .Y(n_391) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_18), .Y(n_685) );
BUFx3_ASAP7_75t_L g234 ( .A(n_19), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_21), .A2(n_49), .B1(n_360), .B2(n_361), .Y(n_359) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_22), .Y(n_223) );
O2A1O1Ixp5_ASAP7_75t_L g379 ( .A1(n_22), .A2(n_256), .B(n_380), .C(n_381), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_24), .Y(n_317) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_26), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g172 ( .A(n_27), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_28), .A2(n_65), .B1(n_288), .B2(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g375 ( .A(n_29), .Y(n_375) );
INVx1_ASAP7_75t_L g95 ( .A(n_30), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_30), .B(n_55), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_31), .B(n_371), .Y(n_422) );
INVx2_ASAP7_75t_L g383 ( .A(n_32), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_33), .Y(n_320) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_34), .Y(n_214) );
INVx2_ASAP7_75t_L g401 ( .A(n_35), .Y(n_401) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_36), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_36), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g341 ( .A(n_37), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_38), .Y(n_217) );
INVx1_ASAP7_75t_L g312 ( .A(n_39), .Y(n_312) );
INVx1_ASAP7_75t_L g283 ( .A(n_40), .Y(n_283) );
INVx1_ASAP7_75t_L g127 ( .A(n_42), .Y(n_127) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_43), .Y(n_245) );
AND2x4_ASAP7_75t_L g259 ( .A(n_43), .B(n_243), .Y(n_259) );
AND2x4_ASAP7_75t_L g306 ( .A(n_43), .B(n_243), .Y(n_306) );
INVx2_ASAP7_75t_L g213 ( .A(n_44), .Y(n_213) );
INVx1_ASAP7_75t_L g346 ( .A(n_45), .Y(n_346) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_46), .Y(n_257) );
INVx1_ASAP7_75t_L g112 ( .A(n_47), .Y(n_112) );
AOI21xp33_ASAP7_75t_SL g166 ( .A1(n_48), .A2(n_167), .B(n_171), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_50), .B(n_338), .Y(n_405) );
OA22x2_ASAP7_75t_L g99 ( .A1(n_51), .A2(n_56), .B1(n_94), .B2(n_98), .Y(n_99) );
INVx1_ASAP7_75t_L g123 ( .A(n_51), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_52), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g153 ( .A(n_53), .Y(n_153) );
INVx1_ASAP7_75t_L g111 ( .A(n_55), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_55), .B(n_121), .Y(n_184) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_55), .Y(n_237) );
OAI21xp33_ASAP7_75t_L g124 ( .A1(n_56), .A2(n_63), .B(n_125), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_57), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_58), .Y(n_373) );
XOR2xp5_ASAP7_75t_L g677 ( .A(n_59), .B(n_83), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_60), .B(n_277), .Y(n_343) );
INVx1_ASAP7_75t_SL g196 ( .A(n_61), .Y(n_196) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_62), .Y(n_81) );
INVx1_ASAP7_75t_L g97 ( .A(n_63), .Y(n_97) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_63), .B(n_75), .Y(n_182) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_66), .Y(n_253) );
BUFx5_ASAP7_75t_L g275 ( .A(n_66), .Y(n_275) );
INVx1_ASAP7_75t_L g303 ( .A(n_66), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_67), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g404 ( .A(n_68), .Y(n_404) );
INVx1_ASAP7_75t_SL g148 ( .A(n_69), .Y(n_148) );
INVx1_ASAP7_75t_L g408 ( .A(n_71), .Y(n_408) );
INVx2_ASAP7_75t_L g325 ( .A(n_72), .Y(n_325) );
INVx2_ASAP7_75t_SL g243 ( .A(n_73), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_74), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_75), .B(n_104), .Y(n_103) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_76), .Y(n_220) );
AO22x2_ASAP7_75t_L g388 ( .A1(n_77), .A2(n_389), .B1(n_393), .B2(n_395), .Y(n_388) );
AO32x2_ASAP7_75t_L g435 ( .A1(n_77), .A2(n_258), .A3(n_384), .B1(n_389), .B2(n_436), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_229), .B1(n_246), .B2(n_260), .C(n_671), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_211), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_82), .B1(n_83), .B2(n_210), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_81), .Y(n_210) );
XOR2xp5_ASAP7_75t_L g672 ( .A(n_82), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_85), .B(n_159), .Y(n_84) );
NOR3xp33_ASAP7_75t_L g85 ( .A(n_86), .B(n_128), .C(n_147), .Y(n_85) );
OAI22xp5_ASAP7_75t_L g86 ( .A1(n_87), .A2(n_112), .B1(n_113), .B2(n_127), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x4_ASAP7_75t_L g90 ( .A(n_91), .B(n_100), .Y(n_90) );
AND2x2_ASAP7_75t_L g143 ( .A(n_91), .B(n_136), .Y(n_143) );
AND2x2_ASAP7_75t_L g165 ( .A(n_91), .B(n_157), .Y(n_165) );
AND2x2_ASAP7_75t_L g199 ( .A(n_91), .B(n_151), .Y(n_199) );
AND2x2_ASAP7_75t_L g91 ( .A(n_92), .B(n_99), .Y(n_91) );
INVx1_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g92 ( .A(n_93), .B(n_96), .Y(n_92) );
NAND2xp33_ASAP7_75t_L g93 ( .A(n_94), .B(n_95), .Y(n_93) );
INVx2_ASAP7_75t_L g98 ( .A(n_94), .Y(n_98) );
INVx3_ASAP7_75t_L g104 ( .A(n_94), .Y(n_104) );
NAND2xp33_ASAP7_75t_L g110 ( .A(n_94), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g125 ( .A(n_94), .Y(n_125) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_94), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_95), .B(n_123), .Y(n_122) );
INVxp67_ASAP7_75t_L g238 ( .A(n_95), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g96 ( .A(n_97), .B(n_98), .Y(n_96) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_97), .A2(n_125), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g135 ( .A(n_99), .Y(n_135) );
AND2x2_ASAP7_75t_L g170 ( .A(n_99), .B(n_134), .Y(n_170) );
AND2x2_ASAP7_75t_L g207 ( .A(n_99), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g126 ( .A(n_101), .Y(n_126) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_106), .Y(n_101) );
AND2x4_ASAP7_75t_L g136 ( .A(n_102), .B(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g151 ( .A(n_102), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g158 ( .A(n_102), .Y(n_158) );
AND2x2_ASAP7_75t_L g204 ( .A(n_102), .B(n_205), .Y(n_204) );
AND2x4_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_104), .B(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g121 ( .A(n_104), .Y(n_121) );
NAND3xp33_ASAP7_75t_L g183 ( .A(n_105), .B(n_120), .C(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g137 ( .A(n_106), .Y(n_137) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g152 ( .A(n_107), .Y(n_152) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx6_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_126), .Y(n_118) );
AND2x4_ASAP7_75t_L g146 ( .A(n_119), .B(n_136), .Y(n_146) );
AND2x4_ASAP7_75t_L g194 ( .A(n_119), .B(n_157), .Y(n_194) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_124), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_123), .Y(n_239) );
AND2x4_ASAP7_75t_L g140 ( .A(n_126), .B(n_133), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_129), .B(n_141), .Y(n_128) );
BUFx12f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx12f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_136), .Y(n_132) );
AND2x4_ASAP7_75t_L g150 ( .A(n_133), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g156 ( .A(n_133), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx8_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B1(n_153), .B2(n_154), .Y(n_147) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g169 ( .A(n_151), .B(n_170), .Y(n_169) );
AND2x4_ASAP7_75t_L g157 ( .A(n_152), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g190 ( .A(n_157), .B(n_170), .Y(n_190) );
NOR3xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_185), .C(n_195), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_161), .B(n_166), .Y(n_160) );
BUFx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_180), .B(n_183), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_179), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B1(n_191), .B2(n_192), .Y(n_185) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_200), .Y(n_195) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx5_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_204), .B(n_207), .Y(n_203) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_206), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_215), .B1(n_227), .B2(n_228), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_212), .Y(n_227) );
XNOR2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_215), .Y(n_228) );
XNOR2xp5_ASAP7_75t_SL g215 ( .A(n_216), .B(n_218), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B1(n_221), .B2(n_226), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g226 ( .A(n_221), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B1(n_224), .B2(n_225), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
BUFx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_240), .Y(n_231) );
INVxp67_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g675 ( .A(n_233), .B(n_240), .Y(n_675) );
AOI211xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_236), .C(n_239), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_244), .Y(n_240) );
OR2x2_ASAP7_75t_L g679 ( .A(n_241), .B(n_245), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_241), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_241), .B(n_244), .Y(n_683) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_258), .Y(n_247) );
OA21x2_ASAP7_75t_L g681 ( .A1(n_248), .A2(n_682), .B(n_683), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_254), .Y(n_248) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_250), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_252), .Y(n_291) );
INVx2_ASAP7_75t_L g377 ( .A(n_252), .Y(n_377) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g277 ( .A(n_253), .Y(n_277) );
INVx2_ASAP7_75t_L g290 ( .A(n_253), .Y(n_290) );
INVx6_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_255), .B(n_305), .Y(n_314) );
INVx4_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_256), .A2(n_390), .B1(n_391), .B2(n_392), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_256), .A2(n_417), .B(n_419), .Y(n_416) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_257), .Y(n_279) );
INVx1_ASAP7_75t_L g293 ( .A(n_257), .Y(n_293) );
INVx3_ASAP7_75t_L g308 ( .A(n_257), .Y(n_308) );
INVx4_ASAP7_75t_L g372 ( .A(n_257), .Y(n_372) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g281 ( .A(n_259), .Y(n_281) );
AND2x2_ASAP7_75t_L g352 ( .A(n_259), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g393 ( .A(n_259), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_569), .Y(n_262) );
NOR2xp33_ASAP7_75t_R g263 ( .A(n_264), .B(n_507), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NOR3xp33_ASAP7_75t_SL g265 ( .A(n_266), .B(n_446), .C(n_482), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_267), .B(n_437), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_347), .B1(n_409), .B2(n_432), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_294), .Y(n_269) );
NAND2x1p5_ASAP7_75t_L g550 ( .A(n_270), .B(n_480), .Y(n_550) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g461 ( .A(n_271), .Y(n_461) );
AND2x2_ASAP7_75t_L g670 ( .A(n_271), .B(n_529), .Y(n_670) );
AND2x2_ASAP7_75t_SL g271 ( .A(n_272), .B(n_286), .Y(n_271) );
NAND2x1p5_ASAP7_75t_L g431 ( .A(n_272), .B(n_286), .Y(n_431) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_278), .B(n_284), .Y(n_272) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
INVx2_ASAP7_75t_L g342 ( .A(n_275), .Y(n_342) );
INVx2_ASAP7_75t_L g420 ( .A(n_275), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_275), .Y(n_424) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g335 ( .A(n_277), .Y(n_335) );
INVx2_ASAP7_75t_L g357 ( .A(n_277), .Y(n_357) );
INVx1_ASAP7_75t_L g418 ( .A(n_277), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_279), .B(n_280), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_279), .A2(n_334), .B(n_336), .C(n_337), .Y(n_333) );
INVx1_ASAP7_75t_L g358 ( .A(n_279), .Y(n_358) );
INVx1_ASAP7_75t_L g392 ( .A(n_279), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g403 ( .A1(n_279), .A2(n_301), .B(n_404), .C(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_280), .B(n_293), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_281), .B(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_281), .B(n_282), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_281), .B(n_282), .Y(n_428) );
BUFx3_ASAP7_75t_L g285 ( .A(n_282), .Y(n_285) );
INVx1_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
INVx1_ASAP7_75t_L g345 ( .A(n_282), .Y(n_345) );
INVx1_ASAP7_75t_L g394 ( .A(n_282), .Y(n_394) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_292), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g310 ( .A(n_290), .Y(n_310) );
AND2x4_ASAP7_75t_L g440 ( .A(n_294), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g669 ( .A(n_294), .B(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_327), .Y(n_294) );
AND2x2_ASAP7_75t_L g429 ( .A(n_295), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g480 ( .A(n_296), .B(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g520 ( .A(n_296), .Y(n_520) );
OR2x2_ASAP7_75t_L g625 ( .A(n_296), .B(n_329), .Y(n_625) );
AO21x2_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_321), .B(n_324), .Y(n_296) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_297), .A2(n_324), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_313), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_304), .B1(n_309), .B2(n_311), .Y(n_298) );
NOR2xp67_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g356 ( .A(n_302), .Y(n_356) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g339 ( .A(n_303), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
NOR3xp33_ASAP7_75t_L g311 ( .A(n_305), .B(n_307), .C(n_312), .Y(n_311) );
AOI221x1_ASAP7_75t_L g366 ( .A1(n_305), .A2(n_367), .B1(n_370), .B2(n_374), .C(n_376), .Y(n_366) );
INVx4_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_307), .A2(n_355), .B1(n_358), .B2(n_359), .Y(n_354) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_308), .A2(n_341), .B(n_342), .C(n_343), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_308), .A2(n_400), .B(n_401), .C(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_318), .B2(n_320), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_318), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g361 ( .A(n_319), .Y(n_361) );
INVx2_ASAP7_75t_L g369 ( .A(n_319), .Y(n_369) );
INVx2_ASAP7_75t_SL g382 ( .A(n_319), .Y(n_382) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx4_ASAP7_75t_L g332 ( .A(n_323), .Y(n_332) );
INVx2_ASAP7_75t_L g364 ( .A(n_323), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g436 ( .A(n_326), .Y(n_436) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g455 ( .A(n_328), .B(n_412), .Y(n_455) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g463 ( .A(n_329), .Y(n_463) );
INVx2_ASAP7_75t_L g481 ( .A(n_329), .Y(n_481) );
AND2x2_ASAP7_75t_L g488 ( .A(n_329), .B(n_457), .Y(n_488) );
INVx1_ASAP7_75t_L g516 ( .A(n_329), .Y(n_516) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_329), .Y(n_602) );
AO31x2_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .A3(n_340), .B(n_344), .Y(n_329) );
INVx2_ASAP7_75t_L g353 ( .A(n_331), .Y(n_353) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g360 ( .A(n_339), .Y(n_360) );
NOR2xp33_ASAP7_75t_SL g344 ( .A(n_345), .B(n_346), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_345), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g347 ( .A(n_348), .B(n_387), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_348), .B(n_541), .Y(n_610) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g506 ( .A(n_349), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_349), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_349), .A2(n_666), .B(n_667), .Y(n_665) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_365), .Y(n_349) );
AND2x2_ASAP7_75t_L g486 ( .A(n_350), .B(n_388), .Y(n_486) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_350), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_350), .B(n_365), .Y(n_548) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g453 ( .A(n_351), .Y(n_453) );
INVx1_ASAP7_75t_L g473 ( .A(n_351), .Y(n_473) );
AOI21x1_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_362), .Y(n_351) );
INVx3_ASAP7_75t_L g380 ( .A(n_360), .Y(n_380) );
INVx1_ASAP7_75t_L g400 ( .A(n_361), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
BUFx3_ASAP7_75t_L g384 ( .A(n_364), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_364), .B(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g414 ( .A(n_364), .Y(n_414) );
AND2x2_ASAP7_75t_L g433 ( .A(n_365), .B(n_396), .Y(n_433) );
INVx1_ASAP7_75t_L g467 ( .A(n_365), .Y(n_467) );
INVx2_ASAP7_75t_L g471 ( .A(n_365), .Y(n_471) );
AND2x2_ASAP7_75t_L g498 ( .A(n_365), .B(n_397), .Y(n_498) );
AO31x2_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_378), .A3(n_384), .B(n_385), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
AND2x2_ASAP7_75t_L g374 ( .A(n_371), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_372), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx2_ASAP7_75t_L g395 ( .A(n_384), .Y(n_395) );
INVx4_ASAP7_75t_L g530 ( .A(n_387), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_387), .B(n_465), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_387), .B(n_547), .Y(n_591) );
AND2x4_ASAP7_75t_L g648 ( .A(n_387), .B(n_470), .Y(n_648) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_396), .Y(n_387) );
AND2x4_ASAP7_75t_L g438 ( .A(n_388), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g543 ( .A(n_388), .Y(n_543) );
INVx1_ASAP7_75t_L g586 ( .A(n_388), .Y(n_586) );
AND2x2_ASAP7_75t_L g472 ( .A(n_396), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx3_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
AND2x4_ASAP7_75t_L g449 ( .A(n_397), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g466 ( .A(n_397), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g542 ( .A(n_397), .Y(n_542) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AO31x2_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .A3(n_406), .B(n_407), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_409), .A2(n_562), .B1(n_565), .B2(n_568), .Y(n_561) );
AND2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_429), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g577 ( .A(n_411), .B(n_515), .Y(n_577) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g442 ( .A(n_412), .Y(n_442) );
AND2x2_ASAP7_75t_L g479 ( .A(n_412), .B(n_431), .Y(n_479) );
INVx2_ASAP7_75t_L g503 ( .A(n_412), .Y(n_503) );
INVx1_ASAP7_75t_L g529 ( .A(n_412), .Y(n_529) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_421), .B(n_428), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g544 ( .A(n_429), .B(n_455), .Y(n_544) );
AND2x2_ASAP7_75t_L g456 ( .A(n_430), .B(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g489 ( .A(n_430), .Y(n_489) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_430), .Y(n_599) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g445 ( .A(n_431), .Y(n_445) );
INVx1_ASAP7_75t_L g567 ( .A(n_431), .Y(n_567) );
AND2x2_ASAP7_75t_L g619 ( .A(n_431), .B(n_503), .Y(n_619) );
NOR2x1_ASAP7_75t_L g557 ( .A(n_432), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AND2x2_ASAP7_75t_L g532 ( .A(n_433), .B(n_452), .Y(n_532) );
AND2x2_ASAP7_75t_L g568 ( .A(n_433), .B(n_476), .Y(n_568) );
OR2x2_ASAP7_75t_L g574 ( .A(n_434), .B(n_575), .Y(n_574) );
BUFx3_ASAP7_75t_L g596 ( .A(n_434), .Y(n_596) );
AND2x4_ASAP7_75t_L g603 ( .A(n_434), .B(n_559), .Y(n_603) );
AND2x2_ASAP7_75t_L g615 ( .A(n_434), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_434), .B(n_466), .Y(n_629) );
AND2x2_ASAP7_75t_L g668 ( .A(n_434), .B(n_477), .Y(n_668) );
BUFx8_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g450 ( .A(n_435), .Y(n_450) );
AND2x2_ASAP7_75t_L g659 ( .A(n_435), .B(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g458 ( .A(n_436), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .C(n_443), .Y(n_437) );
AND2x2_ASAP7_75t_L g494 ( .A(n_438), .B(n_451), .Y(n_494) );
INVx2_ASAP7_75t_L g539 ( .A(n_438), .Y(n_539) );
OAI21xp33_ASAP7_75t_L g552 ( .A1(n_438), .A2(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_438), .B(n_524), .Y(n_634) );
INVx2_ASAP7_75t_SL g505 ( .A(n_439), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_440), .A2(n_496), .B1(n_499), .B2(n_504), .Y(n_495) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g462 ( .A(n_442), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g535 ( .A(n_442), .B(n_457), .Y(n_535) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_444), .B(n_528), .Y(n_579) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g514 ( .A(n_445), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_447), .B(n_468), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_454), .B1(n_459), .B2(n_464), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
AND2x2_ASAP7_75t_L g580 ( .A(n_449), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_449), .B(n_452), .Y(n_650) );
INVx2_ASAP7_75t_L g666 ( .A(n_449), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_450), .B(n_471), .Y(n_564) );
AND2x2_ASAP7_75t_L g637 ( .A(n_450), .B(n_477), .Y(n_637) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx4_ASAP7_75t_L g465 ( .A(n_452), .Y(n_465) );
BUFx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g660 ( .A(n_453), .Y(n_660) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
AND2x2_ASAP7_75t_L g566 ( .A(n_455), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g555 ( .A(n_456), .B(n_462), .Y(n_555) );
AND2x4_ASAP7_75t_L g576 ( .A(n_456), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g460 ( .A(n_457), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g502 ( .A(n_457), .B(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_461), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g662 ( .A(n_462), .Y(n_662) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NAND2x1p5_ASAP7_75t_L g497 ( .A(n_465), .B(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g636 ( .A(n_465), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_466), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g575 ( .A(n_466), .Y(n_575) );
INVx2_ASAP7_75t_L g661 ( .A(n_466), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_474), .B(n_478), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_472), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_470), .B(n_472), .Y(n_667) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_SL g477 ( .A(n_471), .Y(n_477) );
INVx1_ASAP7_75t_L g522 ( .A(n_471), .Y(n_522) );
AND2x2_ASAP7_75t_L g559 ( .A(n_471), .B(n_473), .Y(n_559) );
INVx2_ASAP7_75t_L g476 ( .A(n_473), .Y(n_476) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_473), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_474), .A2(n_532), .B1(n_533), .B2(n_534), .Y(n_531) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
BUFx3_ASAP7_75t_L g553 ( .A(n_476), .Y(n_553) );
OR2x2_ASAP7_75t_L g582 ( .A(n_476), .B(n_481), .Y(n_582) );
AND2x2_ASAP7_75t_L g617 ( .A(n_476), .B(n_541), .Y(n_617) );
INVx1_ASAP7_75t_L g512 ( .A(n_477), .Y(n_512) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g493 ( .A(n_479), .Y(n_493) );
AND2x2_ASAP7_75t_L g533 ( .A(n_479), .B(n_488), .Y(n_533) );
AND2x2_ASAP7_75t_L g584 ( .A(n_479), .B(n_520), .Y(n_584) );
AND2x2_ASAP7_75t_L g601 ( .A(n_479), .B(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g593 ( .A(n_480), .B(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_481), .Y(n_492) );
INVxp67_ASAP7_75t_SL g653 ( .A(n_481), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_487), .B1(n_490), .B2(n_494), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_486), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AND2x2_ASAP7_75t_L g612 ( .A(n_488), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g618 ( .A(n_488), .B(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_493), .B(n_596), .Y(n_595) );
NAND2x1p5_ASAP7_75t_L g605 ( .A(n_496), .B(n_584), .Y(n_605) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g585 ( .A(n_498), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g639 ( .A(n_498), .Y(n_639) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g513 ( .A(n_501), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_502), .Y(n_600) );
OR2x6_ASAP7_75t_L g652 ( .A(n_502), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NOR3x1_ASAP7_75t_L g508 ( .A(n_509), .B(n_536), .C(n_556), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_531), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_513), .B(n_517), .C(n_530), .Y(n_510) );
INVxp67_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x4_ASAP7_75t_L g534 ( .A(n_514), .B(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_515), .Y(n_526) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_523), .C(n_525), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_519), .B(n_619), .Y(n_651) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_520), .B(n_619), .Y(n_646) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g563 ( .A(n_524), .B(n_564), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_525), .A2(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g546 ( .A(n_530), .B(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_534), .A2(n_584), .B1(n_585), .B2(n_587), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .C(n_551), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_544), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g554 ( .A(n_541), .Y(n_554) );
AND2x2_ASAP7_75t_L g558 ( .A(n_541), .B(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_SL g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g616 ( .A(n_548), .Y(n_616) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
INVx1_ASAP7_75t_L g656 ( .A(n_553), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B(n_561), .Y(n_556) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g633 ( .A(n_565), .Y(n_633) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g647 ( .A(n_566), .Y(n_647) );
INVx2_ASAP7_75t_L g613 ( .A(n_567), .Y(n_613) );
NOR2xp33_ASAP7_75t_SL g569 ( .A(n_570), .B(n_643), .Y(n_569) );
NAND4xp75_ASAP7_75t_L g570 ( .A(n_571), .B(n_589), .C(n_606), .D(n_632), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_583), .Y(n_571) );
AOI22xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_576), .B1(n_578), .B2(n_580), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVxp67_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_585), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR3x1_ASAP7_75t_L g589 ( .A(n_590), .B(n_597), .C(n_604), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
OA21x2_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_601), .B(n_603), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVxp67_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
NOR2x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_620), .Y(n_606) );
OAI21xp5_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_611), .B(n_614), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g631 ( .A(n_613), .B(n_625), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_617), .B(n_618), .Y(n_614) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_617), .Y(n_621) );
BUFx3_ASAP7_75t_L g627 ( .A(n_619), .Y(n_627) );
NAND2xp67_ASAP7_75t_L g641 ( .A(n_619), .B(n_642), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B(n_628), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g642 ( .A(n_625), .Y(n_642) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OA21x2_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_635), .Y(n_632) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_640), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR3x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_654), .C(n_663), .Y(n_643) );
AO21x1_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B(n_649), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
AOI21xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B(n_662), .Y(n_654) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI21xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B(n_669), .Y(n_664) );
OAI222xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B1(n_676), .B2(n_678), .C1(n_680), .C2(n_684), .Y(n_671) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
endmodule