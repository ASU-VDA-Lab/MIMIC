module fake_jpeg_2253_n_605 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_605);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_605;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx8_ASAP7_75t_SL g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_56),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_57),
.B(n_62),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_59),
.Y(n_144)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_61),
.B(n_65),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_18),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_70),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_73),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

INVx2_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_75),
.B(n_39),
.Y(n_161)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_43),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g210 ( 
.A(n_78),
.Y(n_210)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_83),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_20),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_87),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_86),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_20),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_112),
.Y(n_157)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_1),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_31),
.B(n_1),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_92),
.Y(n_146)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_94),
.Y(n_199)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_95),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_96),
.Y(n_209)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_97),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_31),
.B(n_1),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_101),
.B(n_103),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_34),
.B(n_2),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_34),
.B(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_104),
.B(n_117),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_105),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_106),
.Y(n_163)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_108),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_37),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_45),
.Y(n_116)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_34),
.B(n_2),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_51),
.B(n_3),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_22),
.B(n_3),
.Y(n_120)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_122),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_40),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_126),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_54),
.B(n_3),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_73),
.A2(n_41),
.B1(n_44),
.B2(n_50),
.Y(n_129)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_129),
.A2(n_132),
.B1(n_141),
.B2(n_152),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_48),
.B1(n_41),
.B2(n_50),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_41),
.B1(n_50),
.B2(n_49),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_78),
.A2(n_41),
.B1(n_50),
.B2(n_49),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_61),
.A2(n_56),
.B(n_22),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_154),
.B(n_12),
.C(n_14),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_58),
.A2(n_49),
.B1(n_47),
.B2(n_44),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_155),
.A2(n_166),
.B1(n_172),
.B2(n_194),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_161),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_71),
.A2(n_49),
.B1(n_47),
.B2(n_44),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_111),
.A2(n_47),
.B1(n_44),
.B2(n_52),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_23),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_175),
.B(n_176),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_67),
.B(n_23),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_75),
.B(n_39),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_177),
.Y(n_263)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_81),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_92),
.Y(n_192)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_100),
.B(n_28),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_216),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_70),
.A2(n_47),
.B1(n_52),
.B2(n_30),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_80),
.A2(n_52),
.B1(n_29),
.B2(n_30),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_196),
.A2(n_198),
.B1(n_213),
.B2(n_4),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_84),
.A2(n_30),
.B1(n_35),
.B2(n_27),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_197),
.A2(n_200),
.B1(n_141),
.B2(n_172),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_127),
.A2(n_29),
.B1(n_35),
.B2(n_27),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_118),
.A2(n_33),
.B1(n_28),
.B2(n_35),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_69),
.A2(n_33),
.B1(n_29),
.B2(n_27),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_203),
.A2(n_204),
.B1(n_220),
.B2(n_15),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_98),
.A2(n_43),
.B1(n_38),
.B2(n_19),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_97),
.Y(n_205)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_206),
.Y(n_224)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_99),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_82),
.A2(n_43),
.B1(n_19),
.B2(n_6),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_95),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_215),
.Y(n_270)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_108),
.Y(n_216)
);

AOI21xp33_ASAP7_75t_SL g217 ( 
.A1(n_68),
.A2(n_19),
.B(n_5),
.Y(n_217)
);

OR2x2_ASAP7_75t_SL g262 ( 
.A(n_217),
.B(n_10),
.Y(n_262)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_76),
.Y(n_218)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_64),
.Y(n_219)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_109),
.A2(n_19),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_161),
.B(n_177),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_222),
.A2(n_242),
.B(n_299),
.C(n_221),
.Y(n_323)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_223),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_130),
.B(n_143),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_226),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_155),
.A2(n_102),
.B1(n_94),
.B2(n_114),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_227),
.A2(n_231),
.B1(n_271),
.B2(n_297),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_145),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_93),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_230),
.B(n_258),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_166),
.A2(n_86),
.B1(n_96),
.B2(n_105),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_149),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_232),
.B(n_234),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_157),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_235),
.Y(n_328)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_124),
.B1(n_115),
.B2(n_89),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_237),
.A2(n_253),
.B1(n_268),
.B2(n_274),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_148),
.A2(n_59),
.B1(n_83),
.B2(n_106),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_238),
.B(n_262),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_144),
.Y(n_240)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_136),
.A2(n_106),
.B(n_66),
.C(n_74),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_77),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_267),
.Y(n_307)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_146),
.Y(n_246)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_251),
.Y(n_330)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_140),
.Y(n_252)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_156),
.A2(n_121),
.B1(n_5),
.B2(n_9),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_170),
.B(n_4),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_254),
.B(n_275),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_255),
.A2(n_260),
.B1(n_223),
.B2(n_265),
.Y(n_351)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_129),
.B(n_16),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_133),
.B(n_4),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_259),
.B(n_264),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_160),
.A2(n_142),
.B1(n_162),
.B2(n_178),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_180),
.B(n_10),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_188),
.Y(n_266)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_169),
.B(n_10),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_186),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_269),
.B(n_272),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_152),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_129),
.B(n_165),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_147),
.B(n_16),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_164),
.B(n_16),
.C(n_181),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_191),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_208),
.B(n_167),
.C(n_209),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_198),
.B(n_197),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_292),
.Y(n_327)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_183),
.Y(n_280)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_135),
.Y(n_281)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_174),
.B1(n_202),
.B2(n_187),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_163),
.B(n_144),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_286),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_167),
.Y(n_284)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_151),
.Y(n_285)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_195),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_135),
.Y(n_287)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_153),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_185),
.B(n_199),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_168),
.Y(n_290)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_290),
.Y(n_352)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_153),
.Y(n_291)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_128),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_168),
.B(n_189),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_300),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_185),
.B(n_132),
.C(n_131),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_273),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_207),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_298),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_213),
.A2(n_194),
.B1(n_196),
.B2(n_137),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_158),
.B(n_173),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_139),
.A2(n_159),
.B1(n_134),
.B2(n_137),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_134),
.B(n_171),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_128),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_301),
.B(n_240),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_279),
.A2(n_138),
.B1(n_150),
.B2(n_159),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_308),
.A2(n_315),
.B1(n_347),
.B2(n_256),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_272),
.A2(n_138),
.B1(n_150),
.B2(n_171),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_282),
.A2(n_221),
.B1(n_202),
.B2(n_174),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_319),
.B(n_294),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_322),
.A2(n_299),
.B1(n_300),
.B2(n_290),
.Y(n_362)
);

OAI21xp33_ASAP7_75t_L g382 ( 
.A1(n_323),
.A2(n_291),
.B(n_285),
.Y(n_382)
);

BUFx24_ASAP7_75t_SL g333 ( 
.A(n_250),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_349),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_242),
.A2(n_295),
.B(n_272),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_339),
.A2(n_340),
.B(n_345),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_258),
.A2(n_245),
.B(n_222),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_344),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_258),
.A2(n_225),
.B(n_278),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_274),
.A2(n_225),
.B1(n_238),
.B2(n_293),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_257),
.B(n_226),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_348),
.B(n_354),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_254),
.B(n_226),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_244),
.B(n_263),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_357),
.Y(n_367)
);

OAI21xp33_ASAP7_75t_SL g380 ( 
.A1(n_351),
.A2(n_266),
.B(n_246),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_275),
.B(n_276),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_353),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_269),
.B(n_230),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_224),
.B(n_228),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_353),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_360),
.B(n_381),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_327),
.A2(n_325),
.B1(n_342),
.B2(n_339),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_361),
.A2(n_354),
.B1(n_337),
.B2(n_356),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_362),
.A2(n_366),
.B1(n_396),
.B2(n_321),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_262),
.B(n_230),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_363),
.A2(n_370),
.B(n_378),
.Y(n_415)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_368),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_347),
.B(n_225),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_310),
.Y(n_371)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_316),
.Y(n_372)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_313),
.B(n_248),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_373),
.B(n_394),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_338),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_SL g437 ( 
.A(n_374),
.B(n_382),
.Y(n_437)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_316),
.Y(n_375)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_375),
.Y(n_422)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_317),
.Y(n_376)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_323),
.A2(n_225),
.B(n_265),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_377),
.A2(n_390),
.B(n_402),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g378 ( 
.A(n_331),
.B(n_277),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_302),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_379),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_380),
.A2(n_393),
.B1(n_326),
.B2(n_302),
.Y(n_406)
);

AO22x1_ASAP7_75t_SL g381 ( 
.A1(n_334),
.A2(n_277),
.B1(n_270),
.B2(n_233),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_335),
.Y(n_384)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_384),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_252),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_387),
.Y(n_424)
);

OA22x2_ASAP7_75t_L g387 ( 
.A1(n_314),
.A2(n_270),
.B1(n_281),
.B2(n_287),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_309),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_388),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_322),
.A2(n_294),
.B1(n_261),
.B2(n_233),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_389),
.A2(n_319),
.B1(n_314),
.B2(n_337),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_340),
.A2(n_284),
.B(n_292),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_391),
.B(n_392),
.Y(n_412)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_315),
.A2(n_241),
.B1(n_229),
.B2(n_239),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_307),
.B(n_224),
.Y(n_394)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_397),
.B(n_401),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_313),
.B(n_343),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_399),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_343),
.B(n_249),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_318),
.B(n_247),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_331),
.A2(n_301),
.B(n_280),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_348),
.B(n_243),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_403),
.B(n_358),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_404),
.A2(n_409),
.B1(n_414),
.B2(n_416),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_406),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_365),
.C(n_398),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_427),
.C(n_436),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_377),
.A2(n_356),
.B1(n_331),
.B2(n_308),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_378),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_366),
.A2(n_356),
.B1(n_334),
.B2(n_329),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_369),
.A2(n_334),
.B1(n_311),
.B2(n_355),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_386),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_417),
.B(n_423),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_369),
.A2(n_360),
.B1(n_395),
.B2(n_370),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_420),
.A2(n_428),
.B1(n_370),
.B2(n_363),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_401),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_387),
.A2(n_355),
.B1(n_321),
.B2(n_312),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_389),
.B1(n_396),
.B2(n_368),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_334),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_429),
.B(n_394),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_385),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_434),
.Y(n_458)
);

AO22x2_ASAP7_75t_SL g433 ( 
.A1(n_362),
.A2(n_332),
.B1(n_305),
.B2(n_324),
.Y(n_433)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_433),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_390),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_365),
.B(n_306),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_364),
.B(n_328),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_440),
.B(n_402),
.C(n_378),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_441),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_442),
.A2(n_446),
.B1(n_460),
.B2(n_461),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_423),
.B(n_372),
.Y(n_443)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_443),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_375),
.Y(n_445)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_445),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_436),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_412),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_449),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_432),
.A2(n_396),
.B(n_381),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_450),
.A2(n_457),
.B(n_463),
.Y(n_483)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_412),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_403),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_454),
.B(n_465),
.C(n_474),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_455),
.B(n_467),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_432),
.A2(n_376),
.B(n_371),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g459 ( 
.A(n_420),
.B(n_381),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_459),
.A2(n_437),
.B(n_421),
.Y(n_481)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_418),
.B(n_383),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_435),
.B(n_367),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_433),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_434),
.A2(n_388),
.B(n_391),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_424),
.A2(n_387),
.B1(n_381),
.B2(n_397),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_464),
.A2(n_466),
.B1(n_469),
.B2(n_470),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_392),
.C(n_326),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_418),
.B(n_424),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_384),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_415),
.A2(n_374),
.B(n_338),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_468),
.A2(n_438),
.B(n_330),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_379),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_410),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_408),
.B(n_387),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_428),
.Y(n_482)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_411),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_472),
.A2(n_430),
.B1(n_426),
.B2(n_419),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_405),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_473),
.A2(n_359),
.B(n_433),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_440),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_475),
.B(n_479),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_415),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_482),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_444),
.A2(n_421),
.B1(n_409),
.B2(n_414),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_485),
.A2(n_488),
.B1(n_482),
.B2(n_481),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_447),
.B(n_416),
.C(n_429),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_486),
.B(n_492),
.C(n_501),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_454),
.B(n_422),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_493),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_444),
.A2(n_446),
.B1(n_459),
.B2(n_464),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_451),
.A2(n_404),
.B1(n_426),
.B2(n_422),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_490),
.A2(n_495),
.B1(n_502),
.B2(n_491),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_411),
.C(n_419),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_430),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_451),
.A2(n_437),
.B1(n_433),
.B2(n_439),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_458),
.A2(n_439),
.B(n_438),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_496),
.A2(n_498),
.B(n_468),
.Y(n_524)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_497),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_499),
.B(n_450),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_448),
.B(n_312),
.C(n_330),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_457),
.A2(n_400),
.B1(n_341),
.B2(n_320),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_441),
.B(n_328),
.C(n_324),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_504),
.C(n_463),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_462),
.B(n_320),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_496),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_506),
.B(n_518),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_480),
.B(n_462),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_507),
.B(n_514),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_508),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_500),
.A2(n_505),
.B1(n_490),
.B2(n_478),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_512),
.A2(n_529),
.B1(n_485),
.B2(n_495),
.Y(n_543)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_476),
.Y(n_515)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_515),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_456),
.Y(n_517)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_489),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_477),
.Y(n_519)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_519),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_479),
.B(n_452),
.C(n_443),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_520),
.B(n_530),
.C(n_503),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_522),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_480),
.B(n_458),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_528),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_524),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_486),
.B(n_473),
.C(n_455),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_499),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_484),
.B(n_456),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_526),
.B(n_449),
.Y(n_532)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_492),
.B(n_445),
.C(n_459),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_531),
.B(n_514),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_532),
.B(n_542),
.Y(n_557)
);

AOI322xp5_ASAP7_75t_SL g534 ( 
.A1(n_517),
.A2(n_469),
.A3(n_467),
.B1(n_475),
.B2(n_461),
.C1(n_466),
.C2(n_453),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_534),
.B(n_548),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_501),
.C(n_487),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_538),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_526),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_493),
.C(n_504),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_539),
.B(n_507),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_527),
.A2(n_483),
.B(n_488),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_543),
.A2(n_508),
.B1(n_512),
.B2(n_530),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_510),
.Y(n_547)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_547),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_547),
.B(n_523),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_551),
.B(n_553),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_541),
.A2(n_527),
.B(n_529),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g567 ( 
.A(n_552),
.B(n_542),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_537),
.B(n_531),
.C(n_539),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_520),
.C(n_513),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_555),
.B(n_562),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_556),
.B(n_561),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_535),
.B(n_516),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_558),
.B(n_564),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_541),
.A2(n_524),
.B(n_509),
.Y(n_559)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_559),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_560),
.A2(n_536),
.B1(n_559),
.B2(n_544),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_521),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_516),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_555),
.Y(n_571)
);

A2O1A1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_532),
.A2(n_522),
.B(n_459),
.C(n_471),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_553),
.B(n_556),
.C(n_550),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_566),
.B(n_571),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_567),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_557),
.A2(n_536),
.B1(n_543),
.B2(n_533),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_573),
.B(n_576),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_SL g575 ( 
.A(n_552),
.B(n_513),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_L g588 ( 
.A(n_575),
.B(n_540),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_565),
.B(n_545),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_557),
.A2(n_540),
.B(n_544),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_577),
.B(n_564),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_567),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_579),
.B(n_587),
.Y(n_593)
);

AOI21xp33_ASAP7_75t_L g590 ( 
.A1(n_580),
.A2(n_572),
.B(n_546),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_560),
.C(n_558),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_583),
.B(n_586),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_569),
.B(n_554),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_585),
.A2(n_498),
.B1(n_502),
.B2(n_453),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_570),
.A2(n_568),
.B1(n_574),
.B2(n_572),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_578),
.B(n_575),
.C(n_573),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g592 ( 
.A1(n_588),
.A2(n_581),
.B(n_585),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_590),
.A2(n_591),
.B(n_581),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_584),
.A2(n_472),
.B(n_470),
.Y(n_591)
);

AO21x2_ASAP7_75t_L g597 ( 
.A1(n_592),
.A2(n_595),
.B(n_579),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_582),
.B(n_400),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_594),
.B(n_400),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_589),
.B(n_593),
.C(n_587),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_596),
.B(n_453),
.C(n_442),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_597),
.B(n_598),
.C(n_599),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_601),
.B(n_460),
.C(n_303),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_602),
.A2(n_600),
.B(n_239),
.Y(n_603)
);

OAI321xp33_ASAP7_75t_L g604 ( 
.A1(n_603),
.A2(n_236),
.A3(n_251),
.B1(n_303),
.B2(n_304),
.C(n_600),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_604),
.B(n_251),
.Y(n_605)
);


endmodule