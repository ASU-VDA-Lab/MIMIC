module fake_netlist_5_2513_n_1834 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1834);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1834;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g178 ( 
.A(n_72),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_43),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_73),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_25),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_56),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_104),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_151),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_87),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_147),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_120),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_62),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_134),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_12),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_108),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_140),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_165),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_136),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_144),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_71),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_79),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_18),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_50),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_39),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_42),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_47),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_25),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_58),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_82),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_56),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_96),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_9),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_6),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_37),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_44),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_4),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_95),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_94),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_34),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_81),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_101),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_102),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_139),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_118),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_97),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_3),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_0),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_9),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_105),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_131),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_35),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_128),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_26),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_163),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_116),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_51),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_112),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_142),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_158),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_77),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_107),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_126),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_88),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_4),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_65),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_143),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_67),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_103),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_170),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_66),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_115),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_172),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_1),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_74),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_100),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_0),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_21),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_83),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_119),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_173),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_154),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_18),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_90),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_109),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_175),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_159),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_93),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_37),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_89),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_54),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_68),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_69),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_17),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_42),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_162),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_156),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_84),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_14),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_6),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_32),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_38),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_122),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_48),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_10),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_50),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_146),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_57),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_123),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_149),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_34),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_168),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_53),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_161),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_135),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_30),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_141),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_129),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_48),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_80),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_59),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_12),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_148),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_58),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_47),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_76),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_64),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_3),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_39),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_55),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_99),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_138),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_106),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_44),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_8),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_40),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_13),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_117),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_111),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_70),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_45),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_35),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_53),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_17),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_41),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_21),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_133),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_150),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_27),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_124),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_1),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_16),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_55),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_52),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_91),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_113),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_169),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_78),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_41),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_85),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_110),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_14),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_61),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_127),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_49),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_330),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_2),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_245),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_209),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_355),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_245),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_219),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_220),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_285),
.B(n_2),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_223),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_182),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_245),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_331),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_199),
.Y(n_372)
);

BUFx2_ASAP7_75t_SL g373 ( 
.A(n_247),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_216),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_349),
.Y(n_375)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_247),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_222),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_224),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_179),
.B(n_5),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_257),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_226),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_317),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_317),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_288),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_227),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_212),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_187),
.B(n_5),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_212),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_232),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_234),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_239),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_204),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_240),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_228),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_206),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_257),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_187),
.B(n_7),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_238),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_257),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g405 ( 
.A(n_187),
.B(n_8),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_242),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_244),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_257),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_248),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_257),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_249),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_269),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_246),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_207),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_250),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_275),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_252),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_218),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_233),
.B(n_11),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_221),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_235),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_281),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_266),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_270),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_288),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_253),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_255),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_292),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_259),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_260),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_294),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_182),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_311),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_322),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_233),
.B(n_11),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_329),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_261),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_286),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_334),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_262),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_291),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_241),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_241),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_303),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_303),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_320),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_293),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_192),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_183),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_194),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_202),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_363),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_180),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_363),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_377),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_362),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_401),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_405),
.B(n_233),
.Y(n_462)
);

XOR2x2_ASAP7_75t_L g463 ( 
.A(n_359),
.B(n_236),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_361),
.B(n_178),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_404),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_371),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_408),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_364),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_379),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_386),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_365),
.B(n_184),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_390),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_392),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_452),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_443),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_376),
.B(n_320),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_R g481 ( 
.A(n_393),
.B(n_263),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_397),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_370),
.B(n_178),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_374),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_444),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_445),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_446),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_369),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_453),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_365),
.B(n_186),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_385),
.B(n_425),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g496 ( 
.A(n_402),
.B(n_189),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_406),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_420),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_450),
.A2(n_213),
.B(n_189),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_387),
.B(n_194),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_366),
.B(n_198),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_407),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_421),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_413),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_424),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_428),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_431),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_366),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_433),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_415),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_436),
.Y(n_514)
);

XNOR2x1_ASAP7_75t_L g515 ( 
.A(n_380),
.B(n_183),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_368),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_417),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_389),
.B(n_213),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_439),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_251),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_426),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_451),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_427),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_429),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_391),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_430),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_395),
.B(n_194),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_449),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_437),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_440),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_380),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_508),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_525),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_496),
.A2(n_360),
.B1(n_367),
.B2(n_432),
.Y(n_536)
);

NOR3xp33_ASAP7_75t_L g537 ( 
.A(n_474),
.B(n_372),
.C(n_383),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_525),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_493),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_493),
.B(n_495),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_251),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_496),
.A2(n_432),
.B1(n_373),
.B2(n_434),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_532),
.A2(n_375),
.B1(n_441),
.B2(n_438),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_394),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_532),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_481),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_467),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_508),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_491),
.B(n_378),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_497),
.Y(n_550)
);

INVx5_ASAP7_75t_L g551 ( 
.A(n_520),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_494),
.B(n_368),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_493),
.B(n_382),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g554 ( 
.A(n_493),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_493),
.B(n_382),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_532),
.B(n_251),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_497),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_503),
.B(n_399),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_532),
.Y(n_559)
);

AO22x2_ASAP7_75t_L g560 ( 
.A1(n_515),
.A2(n_283),
.B1(n_344),
.B2(n_305),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_522),
.B(n_399),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_532),
.B(n_251),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_495),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_467),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_462),
.B(n_251),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_491),
.B(n_384),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_480),
.B(n_396),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_499),
.Y(n_569)
);

BUFx10_ASAP7_75t_L g570 ( 
.A(n_511),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_461),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_456),
.B(n_403),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_501),
.Y(n_574)
);

INVx4_ASAP7_75t_SL g575 ( 
.A(n_520),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_471),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_L g577 ( 
.A(n_520),
.B(n_271),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_499),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_520),
.A2(n_398),
.B1(n_400),
.B2(n_271),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_515),
.A2(n_447),
.B1(n_441),
.B2(n_438),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_500),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_456),
.B(n_403),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_471),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_520),
.A2(n_271),
.B1(n_318),
.B2(n_348),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_462),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_462),
.B(n_409),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_520),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_518),
.B(n_409),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_516),
.B(n_203),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_518),
.B(n_411),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_461),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_462),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_500),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_518),
.B(n_411),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_471),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_471),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_507),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_520),
.B(n_412),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_471),
.B(n_271),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_516),
.Y(n_601)
);

BUFx10_ASAP7_75t_L g602 ( 
.A(n_458),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_507),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_509),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_472),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_465),
.B(n_412),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_515),
.B(n_416),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_473),
.Y(n_608)
);

INVx4_ASAP7_75t_SL g609 ( 
.A(n_471),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_455),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_455),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

AO22x2_ASAP7_75t_L g613 ( 
.A1(n_502),
.A2(n_264),
.B1(n_351),
.B2(n_333),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_502),
.A2(n_422),
.B1(n_416),
.B2(n_447),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_459),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_501),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_518),
.A2(n_271),
.B1(n_318),
.B2(n_319),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_527),
.B(n_225),
.Y(n_618)
);

INVx6_ASAP7_75t_L g619 ( 
.A(n_508),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_465),
.B(n_422),
.Y(n_620)
);

AND2x2_ASAP7_75t_SL g621 ( 
.A(n_454),
.B(n_318),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_509),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_527),
.B(n_318),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_459),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_459),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_487),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_512),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_512),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_508),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_454),
.B(n_180),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_508),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_468),
.B(n_267),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_468),
.B(n_273),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_476),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_464),
.A2(n_318),
.B1(n_229),
.B2(n_289),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_457),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_464),
.B(n_230),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_487),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_464),
.B(n_304),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_464),
.A2(n_290),
.B1(n_302),
.B2(n_312),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_483),
.B(n_304),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_514),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_483),
.B(n_231),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_463),
.B(n_296),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_508),
.Y(n_645)
);

AND2x2_ASAP7_75t_SL g646 ( 
.A(n_457),
.B(n_237),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_514),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_528),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_528),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_510),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_483),
.B(n_254),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_487),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_510),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_510),
.B(n_258),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_L g655 ( 
.A1(n_478),
.A2(n_297),
.B1(n_346),
.B2(n_345),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_487),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_510),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_492),
.B(n_274),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_492),
.B(n_276),
.Y(n_659)
);

INVx5_ASAP7_75t_L g660 ( 
.A(n_479),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_505),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_505),
.B(n_298),
.C(n_337),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_479),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_479),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_484),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_519),
.B(n_265),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_519),
.A2(n_306),
.B1(n_309),
.B2(n_272),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_519),
.B(n_282),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_529),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_463),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_529),
.A2(n_268),
.B1(n_282),
.B2(n_304),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_484),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_484),
.Y(n_673)
);

AND2x2_ASAP7_75t_SL g674 ( 
.A(n_485),
.B(n_282),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_478),
.B(n_282),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_469),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_470),
.Y(n_677)
);

INVx5_ASAP7_75t_L g678 ( 
.A(n_490),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_470),
.Y(n_679)
);

AO22x2_ASAP7_75t_L g680 ( 
.A1(n_463),
.A2(n_489),
.B1(n_488),
.B2(n_486),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_550),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_540),
.B(n_554),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_582),
.B(n_490),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_545),
.B(n_559),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_557),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_564),
.B(n_534),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_569),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_601),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_552),
.B(n_477),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_563),
.A2(n_475),
.B(n_486),
.C(n_488),
.Y(n_690)
);

AOI221xp5_ASAP7_75t_L g691 ( 
.A1(n_560),
.A2(n_313),
.B1(n_335),
.B2(n_217),
.C(n_214),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_549),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_664),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_539),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_664),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_578),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_545),
.B(n_490),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_665),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_584),
.B(n_181),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_585),
.B(n_592),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_564),
.A2(n_489),
.B1(n_300),
.B2(n_217),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_553),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_665),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_551),
.B(n_277),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_585),
.B(n_592),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_588),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_558),
.A2(n_214),
.B(n_210),
.C(n_205),
.Y(n_707)
);

NOR2x1p5_ASAP7_75t_L g708 ( 
.A(n_549),
.B(n_482),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_587),
.B(n_278),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_567),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_676),
.B(n_279),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_539),
.A2(n_651),
.B1(n_643),
.B2(n_637),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_676),
.B(n_280),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_573),
.B(n_498),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_555),
.B(n_284),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_672),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_561),
.B(n_513),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_538),
.B(n_63),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_588),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_607),
.A2(n_316),
.B(n_210),
.C(n_205),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_677),
.B(n_295),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_590),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_621),
.A2(n_299),
.B1(n_332),
.B2(n_341),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_546),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_587),
.B(n_579),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_536),
.A2(n_190),
.B1(n_256),
.B2(n_301),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_567),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_574),
.A2(n_599),
.B(n_562),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_568),
.B(n_485),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_581),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_614),
.B(n_521),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_587),
.B(n_343),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_636),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_568),
.B(n_523),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_679),
.B(n_181),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_644),
.B(n_300),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_593),
.B(n_185),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_630),
.B(n_586),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_651),
.A2(n_313),
.B1(n_316),
.B2(n_314),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_598),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_603),
.B(n_185),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_580),
.B(n_543),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_621),
.B(n_504),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_673),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_590),
.B(n_506),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_673),
.Y(n_746)
);

O2A1O1Ixp5_ASAP7_75t_L g747 ( 
.A1(n_556),
.A2(n_188),
.B(n_357),
.C(n_356),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_604),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_544),
.B(n_517),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_L g750 ( 
.A(n_655),
.B(n_338),
.C(n_342),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_626),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_544),
.B(n_594),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_594),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_606),
.B(n_524),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_620),
.B(n_526),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_587),
.B(n_188),
.Y(n_756)
);

NOR2xp67_ASAP7_75t_L g757 ( 
.A(n_662),
.B(n_190),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_646),
.B(n_530),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_622),
.B(n_75),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_587),
.B(n_191),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_R g761 ( 
.A(n_595),
.B(n_460),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_626),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_638),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_638),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_627),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_628),
.B(n_191),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_642),
.B(n_193),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_651),
.A2(n_314),
.B1(n_308),
.B2(n_327),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_647),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_648),
.B(n_193),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_646),
.B(n_466),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_649),
.B(n_196),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_533),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_L g774 ( 
.A1(n_544),
.A2(n_195),
.B1(n_208),
.B2(n_211),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_650),
.B(n_653),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_652),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_575),
.B(n_196),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_595),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_652),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_674),
.A2(n_357),
.B1(n_356),
.B2(n_354),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_656),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_575),
.B(n_197),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_544),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_657),
.B(n_197),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_637),
.A2(n_323),
.B1(n_327),
.B2(n_328),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_658),
.B(n_354),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_659),
.B(n_353),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_535),
.B(n_353),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_674),
.B(n_350),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_535),
.B(n_350),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_675),
.B(n_310),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_616),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_535),
.B(n_201),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_547),
.B(n_565),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_639),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_656),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_675),
.B(n_618),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_618),
.B(n_310),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_611),
.Y(n_799)
);

OAI221xp5_ASAP7_75t_L g800 ( 
.A1(n_640),
.A2(n_308),
.B1(n_323),
.B2(n_335),
.C(n_328),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_611),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_639),
.B(n_301),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_SL g803 ( 
.A(n_595),
.B(n_347),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_618),
.B(n_167),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_575),
.B(n_200),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_641),
.B(n_200),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_547),
.B(n_326),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_632),
.B(n_326),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_547),
.B(n_325),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_575),
.B(n_201),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_641),
.B(n_307),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_565),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_571),
.B(n_324),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_618),
.A2(n_315),
.B1(n_307),
.B2(n_256),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_602),
.B(n_339),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_666),
.B(n_132),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_542),
.B(n_215),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_616),
.B(n_215),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_613),
.B(n_315),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_589),
.B(n_174),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_637),
.A2(n_287),
.B1(n_243),
.B2(n_19),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_623),
.B(n_171),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_661),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_623),
.B(n_153),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_669),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_666),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_L g827 ( 
.A(n_670),
.B(n_13),
.C(n_15),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_637),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_612),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_612),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_644),
.B(n_22),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_623),
.B(n_137),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_589),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_615),
.Y(n_834)
);

OAI221xp5_ASAP7_75t_L g835 ( 
.A1(n_667),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.C(n_27),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_663),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_556),
.B(n_130),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_826),
.Y(n_838)
);

AOI21xp33_ASAP7_75t_L g839 ( 
.A1(n_789),
.A2(n_589),
.B(n_680),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_694),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_818),
.A2(n_562),
.B(n_654),
.C(n_566),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_738),
.B(n_570),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_689),
.B(n_605),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_728),
.A2(n_541),
.B(n_577),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_836),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_682),
.A2(n_541),
.B(n_577),
.Y(n_846)
);

OAI21xp33_ASAP7_75t_L g847 ( 
.A1(n_701),
.A2(n_560),
.B(n_680),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_702),
.B(n_633),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_816),
.Y(n_849)
);

OAI321xp33_ASAP7_75t_L g850 ( 
.A1(n_835),
.A2(n_589),
.A3(n_671),
.B1(n_617),
.B2(n_560),
.C(n_566),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_818),
.A2(n_654),
.B(n_668),
.C(n_600),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_727),
.B(n_570),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_706),
.B(n_570),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_792),
.A2(n_668),
.B(n_615),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_792),
.A2(n_635),
.B(n_591),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_797),
.A2(n_537),
.B(n_631),
.C(n_663),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_795),
.B(n_623),
.Y(n_857)
);

OAI22xp5_ASAP7_75t_L g858 ( 
.A1(n_706),
.A2(n_613),
.B1(n_680),
.B2(n_631),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_795),
.B(n_623),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_751),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_791),
.A2(n_742),
.B(n_719),
.C(n_722),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_700),
.A2(n_596),
.B(n_548),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_751),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_733),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_705),
.A2(n_533),
.B(n_548),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_L g866 ( 
.A(n_712),
.B(n_643),
.Y(n_866)
);

NOR2x1_ASAP7_75t_L g867 ( 
.A(n_778),
.B(n_576),
.Y(n_867)
);

AO32x1_ASAP7_75t_L g868 ( 
.A1(n_819),
.A2(n_572),
.A3(n_613),
.B1(n_637),
.B2(n_643),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_719),
.A2(n_643),
.B1(n_637),
.B2(n_613),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_686),
.B(n_597),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_722),
.A2(n_643),
.B1(n_619),
.B2(n_583),
.Y(n_871)
);

BUFx4f_ASAP7_75t_L g872 ( 
.A(n_749),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_792),
.A2(n_643),
.B(n_597),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_694),
.A2(n_548),
.B(n_645),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_753),
.B(n_576),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_688),
.Y(n_876)
);

OAI21x1_ASAP7_75t_L g877 ( 
.A1(n_794),
.A2(n_836),
.B(n_775),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_692),
.B(n_608),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_714),
.B(n_608),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_816),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_836),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_753),
.B(n_576),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_762),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_684),
.A2(n_645),
.B(n_629),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_686),
.B(n_624),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_761),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_681),
.B(n_624),
.Y(n_887)
);

O2A1O1Ixp5_ASAP7_75t_L g888 ( 
.A1(n_715),
.A2(n_782),
.B(n_805),
.C(n_810),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_685),
.B(n_610),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_690),
.A2(n_625),
.B(n_610),
.C(n_629),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_752),
.A2(n_625),
.B(n_660),
.C(n_678),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_697),
.A2(n_678),
.B(n_660),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_729),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_752),
.A2(n_619),
.B1(n_625),
.B2(n_634),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_687),
.B(n_619),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_717),
.B(n_634),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_798),
.A2(n_678),
.B(n_634),
.C(n_608),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_816),
.B(n_609),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_773),
.A2(n_609),
.B(n_98),
.Y(n_899)
);

BUFx12f_ASAP7_75t_L g900 ( 
.A(n_708),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_736),
.B(n_602),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_696),
.B(n_609),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_763),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_730),
.B(n_602),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_740),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_821),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_748),
.B(n_28),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_747),
.A2(n_114),
.B(n_86),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_804),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_734),
.B(n_29),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_721),
.A2(n_29),
.B(n_30),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_763),
.Y(n_912)
);

AO21x1_ASAP7_75t_L g913 ( 
.A1(n_837),
.A2(n_31),
.B(n_33),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_740),
.B(n_33),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_765),
.B(n_36),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_710),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_788),
.A2(n_813),
.B(n_790),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_720),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_764),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_769),
.A2(n_60),
.B(n_49),
.C(n_52),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_828),
.A2(n_46),
.B1(n_54),
.B2(n_57),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_776),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_780),
.A2(n_59),
.B1(n_60),
.B2(n_720),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_793),
.A2(n_809),
.B(n_807),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_764),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_796),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_802),
.B(n_806),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_704),
.A2(n_732),
.B(n_709),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_802),
.B(n_806),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_779),
.A2(n_781),
.B(n_812),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_704),
.A2(n_709),
.B(n_711),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_734),
.B(n_808),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_779),
.Y(n_933)
);

NOR3xp33_ASAP7_75t_L g934 ( 
.A(n_743),
.B(n_754),
.C(n_755),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_729),
.A2(n_811),
.B1(n_718),
.B2(n_787),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_693),
.A2(n_829),
.B(n_801),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_713),
.A2(n_786),
.B(n_777),
.Y(n_937)
);

CKINVDCx8_ASAP7_75t_R g938 ( 
.A(n_749),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_693),
.A2(n_716),
.B(n_801),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_781),
.Y(n_940)
);

XOR2xp5_ASAP7_75t_L g941 ( 
.A(n_745),
.B(n_724),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_777),
.A2(n_782),
.B(n_805),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_739),
.A2(n_768),
.B(n_691),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_823),
.Y(n_944)
);

AO21x1_ASAP7_75t_L g945 ( 
.A1(n_837),
.A2(n_718),
.B(n_817),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_811),
.B(n_724),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_817),
.A2(n_699),
.B(n_726),
.C(n_783),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_820),
.B(n_804),
.Y(n_948)
);

CKINVDCx10_ASAP7_75t_R g949 ( 
.A(n_749),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_825),
.B(n_759),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_756),
.A2(n_760),
.B(n_784),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_759),
.B(n_834),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_759),
.B(n_834),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_774),
.B(n_771),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_778),
.B(n_758),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_695),
.B(n_698),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_819),
.B(n_749),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_723),
.A2(n_718),
.B(n_814),
.C(n_757),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_699),
.A2(n_735),
.B(n_800),
.C(n_767),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_803),
.B(n_815),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_833),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_703),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_L g963 ( 
.A(n_785),
.B(n_750),
.C(n_770),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_831),
.B(n_731),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_737),
.B(n_741),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_766),
.B(n_772),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_744),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_744),
.B(n_746),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_799),
.A2(n_830),
.B(n_829),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_820),
.B(n_827),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_820),
.B(n_804),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_822),
.A2(n_824),
.B(n_832),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_820),
.A2(n_797),
.B1(n_789),
.B2(n_738),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_804),
.A2(n_682),
.B(n_554),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_797),
.A2(n_789),
.B1(n_738),
.B2(n_540),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_738),
.B(n_702),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_682),
.A2(n_554),
.B(n_725),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_738),
.B(n_689),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_728),
.A2(n_682),
.B(n_574),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_682),
.A2(n_554),
.B(n_725),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_738),
.B(n_702),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_821),
.A2(n_742),
.B1(n_789),
.B2(n_828),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_818),
.A2(n_728),
.B(n_683),
.C(n_556),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_738),
.B(n_702),
.Y(n_984)
);

OAI21xp33_ASAP7_75t_L g985 ( 
.A1(n_701),
.A2(n_558),
.B(n_552),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_789),
.A2(n_496),
.B1(n_493),
.B2(n_821),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_818),
.A2(n_707),
.B(n_835),
.C(n_563),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_751),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_797),
.A2(n_789),
.B1(n_738),
.B2(n_540),
.Y(n_989)
);

NAND3xp33_ASAP7_75t_SL g990 ( 
.A(n_689),
.B(n_607),
.C(n_580),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_728),
.A2(n_682),
.B(n_574),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_728),
.A2(n_682),
.B(n_574),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_738),
.B(n_702),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_682),
.A2(n_554),
.B(n_725),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_738),
.B(n_689),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_682),
.A2(n_554),
.B(n_725),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_826),
.Y(n_997)
);

OR2x6_ASAP7_75t_SL g998 ( 
.A(n_726),
.B(n_458),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_SL g999 ( 
.A(n_689),
.B(n_607),
.C(n_580),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_682),
.A2(n_554),
.B(n_725),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_728),
.A2(n_682),
.B(n_574),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_L g1002 ( 
.A(n_689),
.B(n_607),
.C(n_558),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_738),
.B(n_702),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_682),
.A2(n_554),
.B(n_725),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_826),
.Y(n_1005)
);

INVx11_ASAP7_75t_L g1006 ( 
.A(n_761),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_728),
.A2(n_682),
.B(n_574),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_930),
.A2(n_877),
.B(n_972),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_936),
.A2(n_939),
.B(n_854),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_936),
.A2(n_939),
.B(n_854),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_978),
.B(n_995),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_946),
.B(n_843),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_976),
.B(n_981),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_864),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_945),
.A2(n_975),
.A3(n_989),
.B(n_861),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_866),
.A2(n_980),
.B(n_977),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_862),
.A2(n_884),
.B(n_865),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_994),
.A2(n_1000),
.B(n_996),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_903),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_927),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_1004),
.A2(n_991),
.B(n_979),
.Y(n_1021)
);

AND2x2_ASAP7_75t_SL g1022 ( 
.A(n_1002),
.B(n_934),
.Y(n_1022)
);

OA21x2_ASAP7_75t_L g1023 ( 
.A1(n_979),
.A2(n_992),
.B(n_991),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_969),
.A2(n_873),
.B(n_874),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_SL g1025 ( 
.A1(n_913),
.A2(n_950),
.B(n_947),
.Y(n_1025)
);

AOI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_985),
.A2(n_982),
.B(n_954),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_984),
.B(n_993),
.Y(n_1027)
);

AO31x2_ASAP7_75t_L g1028 ( 
.A1(n_982),
.A2(n_973),
.A3(n_858),
.B(n_942),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_1003),
.B(n_965),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_849),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_849),
.B(n_880),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_992),
.A2(n_1007),
.B(n_1001),
.Y(n_1032)
);

AND2x2_ASAP7_75t_SL g1033 ( 
.A(n_986),
.B(n_879),
.Y(n_1033)
);

BUFx12f_ASAP7_75t_L g1034 ( 
.A(n_900),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_966),
.B(n_848),
.Y(n_1035)
);

OAI22x1_ASAP7_75t_L g1036 ( 
.A1(n_896),
.A2(n_941),
.B1(n_960),
.B2(n_910),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1001),
.A2(n_1007),
.B(n_952),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_953),
.A2(n_917),
.B(n_924),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_903),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_893),
.B(n_964),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_838),
.Y(n_1041)
);

AOI221xp5_ASAP7_75t_SL g1042 ( 
.A1(n_943),
.A2(n_923),
.B1(n_906),
.B2(n_847),
.C(n_921),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_997),
.Y(n_1043)
);

AND2x6_ASAP7_75t_L g1044 ( 
.A(n_849),
.B(n_880),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_974),
.A2(n_931),
.B(n_937),
.Y(n_1045)
);

AO31x2_ASAP7_75t_L g1046 ( 
.A1(n_891),
.A2(n_856),
.A3(n_951),
.B(n_923),
.Y(n_1046)
);

AOI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_959),
.A2(n_963),
.B(n_929),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1005),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_935),
.B(n_880),
.Y(n_1049)
);

AOI221xp5_ASAP7_75t_L g1050 ( 
.A1(n_990),
.A2(n_999),
.B1(n_906),
.B2(n_839),
.C(n_921),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_983),
.A2(n_888),
.B(n_846),
.Y(n_1051)
);

OAI22x1_ASAP7_75t_L g1052 ( 
.A1(n_970),
.A2(n_842),
.B1(n_914),
.B2(n_961),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_987),
.A2(n_850),
.B(n_958),
.C(n_918),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_898),
.A2(n_909),
.B1(n_948),
.B2(n_971),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_962),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_905),
.B(n_909),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_860),
.Y(n_1057)
);

BUFx4_ASAP7_75t_SL g1058 ( 
.A(n_948),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_SL g1059 ( 
.A1(n_857),
.A2(n_859),
.B(n_902),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_914),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_944),
.B(n_905),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_905),
.B(n_909),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_933),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_844),
.A2(n_855),
.B(n_846),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_852),
.A2(n_904),
.B(n_876),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_840),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_870),
.B(n_907),
.Y(n_1067)
);

CKINVDCx11_ASAP7_75t_R g1068 ( 
.A(n_998),
.Y(n_1068)
);

AOI21x1_ASAP7_75t_L g1069 ( 
.A1(n_928),
.A2(n_968),
.B(n_956),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_870),
.B(n_915),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_901),
.B(n_955),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_922),
.B(n_926),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_909),
.B(n_881),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_885),
.B(n_940),
.Y(n_1074)
);

AOI21x1_ASAP7_75t_L g1075 ( 
.A1(n_875),
.A2(n_882),
.B(n_892),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_878),
.B(n_957),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_845),
.B(n_881),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_863),
.B(n_912),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_932),
.B(n_850),
.Y(n_1079)
);

INVx5_ASAP7_75t_L g1080 ( 
.A(n_840),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_890),
.A2(n_897),
.A3(n_920),
.B(n_911),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_851),
.A2(n_841),
.B(n_898),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_883),
.B(n_919),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_925),
.A2(n_988),
.B(n_967),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_872),
.B(n_853),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_948),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_L g1087 ( 
.A(n_867),
.B(n_895),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_887),
.A2(n_889),
.B(n_899),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_886),
.B(n_894),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_869),
.B(n_871),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_868),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_949),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_908),
.B(n_916),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_938),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_868),
.A2(n_872),
.B(n_1006),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_864),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_864),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_930),
.A2(n_877),
.B(n_936),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_978),
.A2(n_995),
.B(n_982),
.C(n_985),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_903),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_903),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_838),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_840),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1002),
.A2(n_999),
.B(n_990),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_930),
.A2(n_877),
.B(n_936),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_978),
.B(n_727),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_905),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_973),
.B(n_978),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_930),
.A2(n_877),
.B(n_936),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_866),
.A2(n_694),
.B(n_725),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_838),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_978),
.B(n_727),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_978),
.A2(n_995),
.B(n_982),
.C(n_985),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_879),
.B(n_876),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_930),
.A2(n_877),
.B(n_936),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_866),
.A2(n_694),
.B(n_725),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_864),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_870),
.B(n_849),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_866),
.A2(n_694),
.B(n_725),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_864),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_978),
.B(n_995),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_930),
.A2(n_877),
.B(n_936),
.Y(n_1122)
);

O2A1O1Ixp5_ASAP7_75t_L g1123 ( 
.A1(n_978),
.A2(n_995),
.B(n_983),
.C(n_917),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_864),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_SL g1125 ( 
.A1(n_945),
.A2(n_913),
.B(n_950),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_903),
.Y(n_1126)
);

OAI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_978),
.A2(n_995),
.B1(n_982),
.B2(n_906),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_840),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_838),
.Y(n_1129)
);

CKINVDCx14_ASAP7_75t_R g1130 ( 
.A(n_886),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_870),
.B(n_849),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_982),
.A2(n_906),
.B1(n_921),
.B2(n_978),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_866),
.A2(n_694),
.B(n_725),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_870),
.B(n_849),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_930),
.A2(n_877),
.B(n_936),
.Y(n_1135)
);

AND2x6_ASAP7_75t_L g1136 ( 
.A(n_849),
.B(n_880),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_983),
.A2(n_888),
.B(n_975),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_870),
.B(n_849),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_978),
.B(n_995),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_1006),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_864),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_978),
.B(n_995),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_849),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_930),
.A2(n_877),
.B(n_936),
.Y(n_1144)
);

INVx4_ASAP7_75t_L g1145 ( 
.A(n_905),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_961),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_983),
.A2(n_888),
.B(n_975),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_978),
.A2(n_995),
.B1(n_1002),
.B2(n_973),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_978),
.B(n_995),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_978),
.B(n_995),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_978),
.B(n_995),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_931),
.A2(n_937),
.B(n_928),
.Y(n_1152)
);

NOR2x1_ASAP7_75t_R g1153 ( 
.A(n_886),
.B(n_458),
.Y(n_1153)
);

AOI21x1_ASAP7_75t_SL g1154 ( 
.A1(n_927),
.A2(n_929),
.B(n_859),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1130),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1041),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1012),
.B(n_1106),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1080),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_1080),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1112),
.B(n_1139),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1038),
.A2(n_1037),
.B(n_1045),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1060),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1055),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1139),
.B(n_1011),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1121),
.A2(n_1150),
.B1(n_1149),
.B2(n_1151),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1118),
.B(n_1131),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1127),
.A2(n_1132),
.B1(n_1050),
.B2(n_1026),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1043),
.Y(n_1168)
);

O2A1O1Ixp5_ASAP7_75t_SL g1169 ( 
.A1(n_1047),
.A2(n_1108),
.B(n_1137),
.C(n_1147),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1014),
.Y(n_1170)
);

CKINVDCx16_ASAP7_75t_R g1171 ( 
.A(n_1034),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1099),
.A2(n_1113),
.B(n_1148),
.C(n_1104),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1064),
.A2(n_1018),
.B(n_1110),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1118),
.B(n_1131),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1048),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1142),
.A2(n_1127),
.B1(n_1033),
.B2(n_1022),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_1117),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1060),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1141),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1099),
.B(n_1113),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1029),
.B(n_1035),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1071),
.B(n_1076),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1033),
.A2(n_1022),
.B1(n_1071),
.B2(n_1108),
.Y(n_1183)
);

INVx5_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1098),
.A2(n_1115),
.B(n_1105),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1102),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1111),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1013),
.B(n_1027),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1040),
.B(n_1020),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1116),
.A2(n_1119),
.B(n_1133),
.Y(n_1190)
);

BUFx12f_ASAP7_75t_L g1191 ( 
.A(n_1034),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1132),
.B(n_1020),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1129),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1086),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1118),
.B(n_1131),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1079),
.A2(n_1093),
.B1(n_1090),
.B2(n_1023),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1079),
.A2(n_1090),
.B1(n_1036),
.B2(n_1049),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1097),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1080),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1120),
.B(n_1124),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1023),
.A2(n_1082),
.B(n_1123),
.Y(n_1201)
);

AND2x4_ASAP7_75t_SL g1202 ( 
.A(n_1107),
.B(n_1145),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1042),
.B(n_1090),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1134),
.B(n_1138),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1023),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1146),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1123),
.A2(n_1051),
.B(n_1053),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1025),
.A2(n_1067),
.B(n_1070),
.C(n_1072),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1086),
.A2(n_1091),
.B1(n_1063),
.B2(n_1095),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1057),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1094),
.A2(n_1085),
.B1(n_1086),
.B2(n_1130),
.Y(n_1211)
);

AND2x4_ASAP7_75t_L g1212 ( 
.A(n_1134),
.B(n_1138),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1019),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1078),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1134),
.B(n_1138),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1065),
.B(n_1114),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1146),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1019),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1066),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1083),
.Y(n_1220)
);

BUFx4f_ASAP7_75t_L g1221 ( 
.A(n_1086),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1052),
.A2(n_1089),
.B1(n_1094),
.B2(n_1054),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1039),
.Y(n_1223)
);

OR2x6_ASAP7_75t_SL g1224 ( 
.A(n_1140),
.B(n_1061),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1058),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1107),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1068),
.Y(n_1227)
);

CKINVDCx20_ASAP7_75t_R g1228 ( 
.A(n_1068),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1066),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1028),
.B(n_1074),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1145),
.Y(n_1231)
);

AOI21xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1056),
.A2(n_1062),
.B(n_1031),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_L g1233 ( 
.A(n_1153),
.B(n_1031),
.C(n_1062),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1030),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1103),
.Y(n_1235)
);

BUFx12f_ASAP7_75t_L g1236 ( 
.A(n_1030),
.Y(n_1236)
);

INVx5_ASAP7_75t_L g1237 ( 
.A(n_1044),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1028),
.B(n_1100),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1125),
.A2(n_1101),
.B1(n_1126),
.B2(n_1087),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1028),
.B(n_1101),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1024),
.A2(n_1088),
.B(n_1009),
.C(n_1010),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1017),
.A2(n_1008),
.B(n_1144),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1028),
.B(n_1126),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1030),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1092),
.B(n_1056),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_1073),
.B(n_1077),
.C(n_1143),
.Y(n_1246)
);

O2A1O1Ixp5_ASAP7_75t_L g1247 ( 
.A1(n_1152),
.A2(n_1075),
.B(n_1069),
.C(n_1073),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1030),
.B(n_1143),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1008),
.A2(n_1109),
.B(n_1135),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1143),
.B(n_1015),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1084),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1143),
.B(n_1128),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1015),
.B(n_1046),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1015),
.B(n_1046),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1058),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1015),
.B(n_1046),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1046),
.B(n_1081),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1081),
.B(n_1091),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1128),
.B(n_1044),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1044),
.B(n_1136),
.Y(n_1260)
);

O2A1O1Ixp5_ASAP7_75t_SL g1261 ( 
.A1(n_1154),
.A2(n_1059),
.B(n_1081),
.C(n_1122),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1044),
.B(n_1136),
.Y(n_1262)
);

INVx5_ASAP7_75t_SL g1263 ( 
.A(n_1136),
.Y(n_1263)
);

BUFx12f_ASAP7_75t_L g1264 ( 
.A(n_1136),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1136),
.B(n_1081),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_1154),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1059),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1032),
.A2(n_1021),
.B(n_1016),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_1080),
.B(n_909),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1118),
.B(n_1131),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1130),
.Y(n_1271)
);

CKINVDCx11_ASAP7_75t_R g1272 ( 
.A(n_1034),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1014),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1012),
.B(n_1106),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1012),
.B(n_978),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1118),
.B(n_1131),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1032),
.A2(n_1021),
.B(n_1016),
.Y(n_1277)
);

BUFx2_ASAP7_75t_L g1278 ( 
.A(n_1014),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1139),
.B(n_978),
.Y(n_1279)
);

BUFx4f_ASAP7_75t_L g1280 ( 
.A(n_1034),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1014),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1041),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1012),
.B(n_1106),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1041),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1014),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_SL g1286 ( 
.A(n_1096),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1055),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1096),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1012),
.B(n_1106),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1012),
.B(n_1106),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1032),
.A2(n_1021),
.B(n_1016),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1139),
.B(n_995),
.C(n_978),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1041),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1032),
.A2(n_1021),
.B(n_1016),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1014),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1032),
.A2(n_1021),
.B(n_1016),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1139),
.A2(n_978),
.B(n_995),
.C(n_985),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1012),
.B(n_1106),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_1097),
.B(n_1096),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1080),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1118),
.B(n_1131),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1032),
.A2(n_1021),
.B(n_1016),
.Y(n_1302)
);

BUFx2_ASAP7_75t_R g1303 ( 
.A(n_1224),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1167),
.A2(n_1292),
.B1(n_1176),
.B2(n_1279),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1156),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1165),
.B(n_1279),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1168),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1198),
.Y(n_1308)
);

INVx4_ASAP7_75t_L g1309 ( 
.A(n_1184),
.Y(n_1309)
);

AOI21xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1164),
.A2(n_1216),
.B(n_1171),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1210),
.Y(n_1311)
);

NAND2x1p5_ASAP7_75t_L g1312 ( 
.A(n_1184),
.B(n_1237),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1264),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1172),
.B(n_1183),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1197),
.B(n_1203),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1175),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1221),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1186),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1187),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1164),
.A2(n_1188),
.B1(n_1181),
.B2(n_1222),
.Y(n_1320)
);

BUFx8_ASAP7_75t_SL g1321 ( 
.A(n_1191),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1188),
.B(n_1181),
.Y(n_1322)
);

AOI21xp33_ASAP7_75t_L g1323 ( 
.A1(n_1167),
.A2(n_1297),
.B(n_1208),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1184),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1180),
.A2(n_1275),
.B1(n_1192),
.B2(n_1203),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1160),
.B(n_1157),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1182),
.B(n_1192),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1221),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1180),
.A2(n_1227),
.B1(n_1283),
.B2(n_1298),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1196),
.B(n_1240),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1287),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1196),
.A2(n_1290),
.B1(n_1289),
.B2(n_1274),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1211),
.A2(n_1177),
.B1(n_1285),
.B2(n_1206),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1184),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1189),
.B(n_1214),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1201),
.A2(n_1207),
.B(n_1173),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1233),
.A2(n_1211),
.B1(n_1207),
.B2(n_1220),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1193),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1237),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1245),
.A2(n_1281),
.B1(n_1170),
.B2(n_1179),
.Y(n_1340)
);

OAI21xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1169),
.A2(n_1239),
.B(n_1262),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1213),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1273),
.A2(n_1295),
.B1(n_1278),
.B2(n_1299),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1166),
.B(n_1174),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1282),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1253),
.B(n_1254),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1177),
.A2(n_1285),
.B1(n_1206),
.B2(n_1246),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1218),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1284),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1256),
.B(n_1223),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1293),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1237),
.A2(n_1178),
.B1(n_1162),
.B2(n_1239),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1228),
.A2(n_1286),
.B1(n_1263),
.B2(n_1271),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1162),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1178),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1265),
.A2(n_1288),
.B1(n_1232),
.B2(n_1225),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1268),
.A2(n_1302),
.B1(n_1277),
.B2(n_1296),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1200),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1272),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1238),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1265),
.A2(n_1255),
.B1(n_1263),
.B2(n_1217),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1244),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1263),
.A2(n_1262),
.B1(n_1286),
.B2(n_1230),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1238),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1243),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1243),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1258),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1260),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1155),
.A2(n_1280),
.B1(n_1266),
.B2(n_1209),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1259),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1291),
.A2(n_1294),
.B1(n_1230),
.B2(n_1257),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1251),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1267),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1269),
.A2(n_1301),
.B1(n_1276),
.B2(n_1270),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1209),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1236),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1280),
.A2(n_1231),
.B1(n_1226),
.B2(n_1194),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1248),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1269),
.A2(n_1301),
.B1(n_1276),
.B2(n_1270),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1195),
.A2(n_1215),
.B1(n_1204),
.B2(n_1212),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1195),
.A2(n_1215),
.B1(n_1204),
.B2(n_1212),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1248),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1158),
.B(n_1159),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1250),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1234),
.Y(n_1385)
);

CKINVDCx11_ASAP7_75t_R g1386 ( 
.A(n_1252),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1219),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1159),
.B(n_1300),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1202),
.Y(n_1389)
);

BUFx8_ASAP7_75t_L g1390 ( 
.A(n_1252),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1205),
.B(n_1241),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1161),
.B(n_1185),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1247),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1229),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1247),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1235),
.Y(n_1396)
);

INVx4_ASAP7_75t_SL g1397 ( 
.A(n_1199),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1300),
.A2(n_1199),
.B1(n_1190),
.B2(n_1185),
.Y(n_1398)
);

OAI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1261),
.A2(n_995),
.B1(n_978),
.B2(n_803),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1249),
.A2(n_1008),
.B(n_1242),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1249),
.A2(n_1008),
.B(n_1242),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1170),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1156),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1281),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1264),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1156),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1198),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1281),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1163),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1198),
.Y(n_1410)
);

NAND2x1p5_ASAP7_75t_L g1411 ( 
.A(n_1184),
.B(n_1237),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1156),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1292),
.A2(n_995),
.B1(n_978),
.B2(n_1139),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1292),
.A2(n_995),
.B1(n_978),
.B2(n_1139),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1156),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1163),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1156),
.Y(n_1417)
);

AO21x1_ASAP7_75t_L g1418 ( 
.A1(n_1207),
.A2(n_1108),
.B(n_1093),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1156),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1156),
.Y(n_1420)
);

BUFx2_ASAP7_75t_SL g1421 ( 
.A(n_1286),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1156),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1176),
.B(n_1172),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1156),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1249),
.A2(n_1008),
.B(n_1242),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1390),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1372),
.Y(n_1427)
);

AO21x1_ASAP7_75t_SL g1428 ( 
.A1(n_1323),
.A2(n_1375),
.B(n_1337),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1360),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1413),
.A2(n_1414),
.B1(n_1423),
.B2(n_1314),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1308),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1364),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1365),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1326),
.B(n_1306),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1366),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1373),
.Y(n_1436)
);

AO21x1_ASAP7_75t_SL g1437 ( 
.A1(n_1337),
.A2(n_1371),
.B(n_1391),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1390),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1322),
.B(n_1327),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1327),
.B(n_1320),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1350),
.B(n_1384),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1321),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1367),
.Y(n_1443)
);

AO31x2_ASAP7_75t_L g1444 ( 
.A1(n_1418),
.A2(n_1393),
.A3(n_1395),
.B(n_1363),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1391),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1330),
.B(n_1346),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1314),
.B(n_1423),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1400),
.A2(n_1425),
.B(n_1401),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1407),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1371),
.B(n_1315),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1392),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_SL g1452 ( 
.A1(n_1418),
.A2(n_1356),
.B(n_1325),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1392),
.Y(n_1453)
);

BUFx4f_ASAP7_75t_L g1454 ( 
.A(n_1312),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1341),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1354),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1315),
.B(n_1325),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1410),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1355),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1398),
.B(n_1370),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1336),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1396),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1390),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1304),
.A2(n_1329),
.B1(n_1332),
.B2(n_1333),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1305),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1307),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1304),
.B(n_1335),
.Y(n_1467)
);

AOI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1361),
.A2(n_1352),
.B(n_1318),
.Y(n_1468)
);

NAND3x1_ASAP7_75t_L g1469 ( 
.A(n_1316),
.B(n_1403),
.C(n_1422),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1399),
.A2(n_1310),
.B(n_1347),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1370),
.B(n_1324),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1319),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1332),
.B(n_1338),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1345),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1349),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1351),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1312),
.Y(n_1477)
);

AO21x2_ASAP7_75t_L g1478 ( 
.A1(n_1406),
.A2(n_1424),
.B(n_1415),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1412),
.B(n_1417),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1419),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1362),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1420),
.A2(n_1394),
.B(n_1387),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1383),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1311),
.Y(n_1484)
);

AO21x1_ASAP7_75t_SL g1485 ( 
.A1(n_1357),
.A2(n_1378),
.B(n_1382),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1411),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1358),
.B(n_1404),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1342),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1331),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1309),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1348),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1357),
.B(n_1409),
.Y(n_1492)
);

BUFx8_ASAP7_75t_SL g1493 ( 
.A(n_1359),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1408),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1340),
.B(n_1416),
.Y(n_1495)
);

NAND2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1309),
.B(n_1334),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1324),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1334),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1339),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1369),
.B(n_1368),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1383),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1388),
.Y(n_1502)
);

INVxp67_ASAP7_75t_R g1503 ( 
.A(n_1500),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1427),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1439),
.B(n_1343),
.Y(n_1505)
);

INVxp67_ASAP7_75t_SL g1506 ( 
.A(n_1488),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1436),
.Y(n_1507)
);

AOI21xp33_ASAP7_75t_L g1508 ( 
.A1(n_1470),
.A2(n_1377),
.B(n_1339),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1460),
.B(n_1368),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1434),
.B(n_1402),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1481),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1478),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1460),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1457),
.B(n_1385),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1449),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1446),
.B(n_1344),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1446),
.B(n_1344),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1458),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1464),
.A2(n_1353),
.B(n_1381),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1445),
.B(n_1421),
.Y(n_1520)
);

OAI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1430),
.A2(n_1380),
.B1(n_1374),
.B2(n_1379),
.C(n_1328),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1478),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1482),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1457),
.B(n_1397),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1482),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1467),
.B(n_1386),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

NAND2xp33_ASAP7_75t_R g1528 ( 
.A(n_1442),
.B(n_1389),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1451),
.B(n_1376),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1429),
.B(n_1397),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1493),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1451),
.B(n_1376),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1441),
.B(n_1397),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1453),
.B(n_1313),
.Y(n_1534)
);

AOI222xp33_ASAP7_75t_L g1535 ( 
.A1(n_1440),
.A2(n_1447),
.B1(n_1359),
.B2(n_1473),
.C1(n_1494),
.C2(n_1431),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1460),
.B(n_1453),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1441),
.B(n_1397),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1441),
.B(n_1303),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1453),
.B(n_1313),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1460),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1465),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1465),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1450),
.B(n_1447),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1429),
.B(n_1317),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1450),
.B(n_1466),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_1491),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1466),
.B(n_1472),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1426),
.A2(n_1313),
.B1(n_1405),
.B2(n_1328),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1472),
.B(n_1386),
.Y(n_1549)
);

OAI221xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1519),
.A2(n_1455),
.B1(n_1495),
.B2(n_1500),
.C(n_1487),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1543),
.B(n_1473),
.Y(n_1551)
);

OAI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1519),
.A2(n_1455),
.B1(n_1481),
.B2(n_1426),
.C(n_1463),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1515),
.B(n_1459),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1507),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1518),
.B(n_1459),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1535),
.A2(n_1405),
.B(n_1468),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_L g1557 ( 
.A1(n_1535),
.A2(n_1508),
.B(n_1505),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1508),
.B(n_1492),
.C(n_1443),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1468),
.Y(n_1559)
);

AOI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1510),
.A2(n_1452),
.B1(n_1443),
.B2(n_1462),
.C(n_1476),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1538),
.A2(n_1405),
.B(n_1496),
.Y(n_1561)
);

NAND3xp33_ASAP7_75t_L g1562 ( 
.A(n_1520),
.B(n_1492),
.C(n_1497),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1538),
.A2(n_1405),
.B(n_1496),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1536),
.B(n_1437),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1521),
.A2(n_1428),
.B1(n_1452),
.B2(n_1549),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1511),
.B(n_1456),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1548),
.B(n_1501),
.C(n_1317),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1498),
.C(n_1497),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1549),
.A2(n_1496),
.B(n_1477),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1536),
.B(n_1444),
.Y(n_1570)
);

NAND3xp33_ASAP7_75t_L g1571 ( 
.A(n_1529),
.B(n_1498),
.C(n_1501),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1511),
.A2(n_1454),
.B1(n_1438),
.B2(n_1463),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1545),
.B(n_1444),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1514),
.B(n_1456),
.Y(n_1574)
);

AND2x2_ASAP7_75t_SL g1575 ( 
.A(n_1513),
.B(n_1454),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1523),
.A2(n_1461),
.B(n_1448),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1545),
.B(n_1444),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1529),
.B(n_1435),
.C(n_1433),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1513),
.B(n_1444),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1530),
.A2(n_1469),
.B(n_1454),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1530),
.B(n_1502),
.C(n_1483),
.Y(n_1581)
);

NAND4xp25_ASAP7_75t_L g1582 ( 
.A(n_1544),
.B(n_1474),
.C(n_1475),
.D(n_1476),
.Y(n_1582)
);

OAI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1534),
.A2(n_1438),
.B1(n_1463),
.B2(n_1426),
.C(n_1486),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1506),
.B(n_1475),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1524),
.A2(n_1537),
.B(n_1533),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_SL g1586 ( 
.A(n_1531),
.B(n_1532),
.C(n_1534),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1532),
.B(n_1432),
.C(n_1433),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_L g1588 ( 
.A1(n_1524),
.A2(n_1435),
.B(n_1432),
.Y(n_1588)
);

NAND3xp33_ASAP7_75t_L g1589 ( 
.A(n_1539),
.B(n_1499),
.C(n_1480),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1503),
.A2(n_1454),
.B1(n_1438),
.B2(n_1469),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1546),
.B(n_1480),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1544),
.A2(n_1462),
.B1(n_1479),
.B2(n_1489),
.C(n_1484),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1516),
.A2(n_1428),
.B1(n_1485),
.B2(n_1471),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1540),
.B(n_1444),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1509),
.A2(n_1477),
.B1(n_1486),
.B2(n_1490),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1576),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1554),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1559),
.B(n_1512),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1559),
.B(n_1512),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1573),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

INVx2_ASAP7_75t_SL g1602 ( 
.A(n_1570),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1577),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1576),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1579),
.B(n_1594),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1551),
.B(n_1522),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1557),
.A2(n_1516),
.B1(n_1517),
.B2(n_1509),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1584),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1591),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1552),
.A2(n_1517),
.B1(n_1509),
.B2(n_1485),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1564),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1574),
.B(n_1525),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1575),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1527),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1589),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1578),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1587),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1568),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1553),
.B(n_1504),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1580),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1582),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1575),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1597),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1604),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1615),
.B(n_1592),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1615),
.B(n_1560),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1602),
.B(n_1503),
.Y(n_1627)
);

NAND4xp25_ASAP7_75t_L g1628 ( 
.A(n_1620),
.B(n_1550),
.C(n_1558),
.D(n_1556),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1616),
.B(n_1598),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1616),
.B(n_1555),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1603),
.B(n_1585),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1615),
.B(n_1588),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1617),
.B(n_1562),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1597),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1597),
.Y(n_1635)
);

AOI21xp33_ASAP7_75t_SL g1636 ( 
.A1(n_1620),
.A2(n_1528),
.B(n_1583),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1617),
.B(n_1547),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1619),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1613),
.Y(n_1639)
);

OAI33xp33_ASAP7_75t_L g1640 ( 
.A1(n_1617),
.A2(n_1566),
.A3(n_1590),
.B1(n_1572),
.B2(n_1541),
.B3(n_1542),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1616),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1619),
.Y(n_1642)
);

INVxp67_ASAP7_75t_SL g1643 ( 
.A(n_1616),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1603),
.B(n_1569),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1619),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1602),
.B(n_1595),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1602),
.B(n_1593),
.Y(n_1647)
);

NAND2xp33_ASAP7_75t_L g1648 ( 
.A(n_1621),
.B(n_1567),
.Y(n_1648)
);

NOR4xp25_ASAP7_75t_L g1649 ( 
.A(n_1621),
.B(n_1565),
.C(n_1586),
.D(n_1563),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1599),
.B(n_1571),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1596),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1623),
.Y(n_1652)
);

NAND2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1639),
.B(n_1613),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1639),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1623),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1634),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1646),
.B(n_1620),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1634),
.Y(n_1658)
);

INVxp67_ASAP7_75t_SL g1659 ( 
.A(n_1641),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1635),
.Y(n_1660)
);

AOI222xp33_ASAP7_75t_L g1661 ( 
.A1(n_1648),
.A2(n_1621),
.B1(n_1565),
.B2(n_1618),
.C1(n_1610),
.C2(n_1613),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1631),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1626),
.Y(n_1663)
);

OAI33xp33_ASAP7_75t_L g1664 ( 
.A1(n_1626),
.A2(n_1618),
.A3(n_1614),
.B1(n_1612),
.B2(n_1608),
.B3(n_1609),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1651),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1625),
.B(n_1600),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1646),
.B(n_1602),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1631),
.B(n_1605),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1644),
.B(n_1605),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1651),
.Y(n_1670)
);

NOR2x1_ASAP7_75t_L g1671 ( 
.A(n_1628),
.B(n_1613),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1625),
.B(n_1632),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1651),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1641),
.Y(n_1674)
);

NOR2xp67_ASAP7_75t_L g1675 ( 
.A(n_1636),
.B(n_1613),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1644),
.B(n_1605),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1643),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1633),
.B(n_1614),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1632),
.B(n_1608),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1647),
.B(n_1611),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1643),
.B(n_1600),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1649),
.B(n_1613),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1647),
.B(n_1600),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1633),
.B(n_1606),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1647),
.B(n_1627),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1638),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1624),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1636),
.B(n_1321),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1629),
.B(n_1601),
.Y(n_1689)
);

NAND2x1p5_ASAP7_75t_L g1690 ( 
.A(n_1627),
.B(n_1622),
.Y(n_1690)
);

INVxp67_ASAP7_75t_L g1691 ( 
.A(n_1630),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1624),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1629),
.B(n_1606),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1652),
.Y(n_1694)
);

INVx3_ASAP7_75t_L g1695 ( 
.A(n_1653),
.Y(n_1695)
);

BUFx2_ASAP7_75t_SL g1696 ( 
.A(n_1675),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1677),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1652),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1655),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1663),
.B(n_1672),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1675),
.B(n_1638),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1653),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1671),
.A2(n_1628),
.B1(n_1640),
.B2(n_1607),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1677),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1674),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1690),
.B(n_1642),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1678),
.B(n_1666),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1654),
.Y(n_1708)
);

INVx4_ASAP7_75t_L g1709 ( 
.A(n_1653),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1655),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1688),
.B(n_1682),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1656),
.Y(n_1712)
);

NAND3xp33_ASAP7_75t_L g1713 ( 
.A(n_1671),
.B(n_1649),
.C(n_1650),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1665),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1690),
.B(n_1642),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1666),
.B(n_1678),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1690),
.B(n_1645),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1654),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1667),
.B(n_1622),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1657),
.A2(n_1610),
.B1(n_1622),
.B2(n_1650),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1665),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1668),
.B(n_1645),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1665),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1656),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1667),
.B(n_1622),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1674),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1670),
.Y(n_1727)
);

AND3x1_ASAP7_75t_L g1728 ( 
.A(n_1657),
.B(n_1561),
.C(n_1622),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1658),
.Y(n_1729)
);

AOI222xp33_ASAP7_75t_L g1730 ( 
.A1(n_1713),
.A2(n_1664),
.B1(n_1640),
.B2(n_1662),
.C1(n_1659),
.C2(n_1691),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1713),
.A2(n_1661),
.B(n_1662),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1711),
.A2(n_1679),
.B(n_1684),
.C(n_1622),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1709),
.B(n_1708),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1711),
.Y(n_1734)
);

NOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1696),
.B(n_1684),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1703),
.A2(n_1661),
.B1(n_1685),
.B2(n_1668),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1630),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1703),
.A2(n_1685),
.B1(n_1669),
.B2(n_1676),
.Y(n_1738)
);

AOI21xp33_ASAP7_75t_L g1739 ( 
.A1(n_1700),
.A2(n_1686),
.B(n_1693),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1708),
.B(n_1669),
.Y(n_1740)
);

NAND2x1p5_ASAP7_75t_L g1741 ( 
.A(n_1709),
.B(n_1676),
.Y(n_1741)
);

NOR2x1_ASAP7_75t_L g1742 ( 
.A(n_1696),
.B(n_1686),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1705),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1707),
.B(n_1693),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1695),
.Y(n_1746)
);

OR2x6_ASAP7_75t_L g1747 ( 
.A(n_1696),
.B(n_1681),
.Y(n_1747)
);

AOI21xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1720),
.A2(n_1716),
.B(n_1702),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1720),
.A2(n_1680),
.B1(n_1683),
.B2(n_1607),
.Y(n_1749)
);

O2A1O1Ixp5_ASAP7_75t_L g1750 ( 
.A1(n_1709),
.A2(n_1681),
.B(n_1689),
.C(n_1660),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1707),
.B(n_1637),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1719),
.B(n_1725),
.Y(n_1752)
);

OAI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1709),
.A2(n_1718),
.B1(n_1695),
.B2(n_1702),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1726),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1726),
.Y(n_1755)
);

NAND3xp33_ASAP7_75t_SL g1756 ( 
.A(n_1731),
.B(n_1718),
.C(n_1709),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1734),
.B(n_1716),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1752),
.B(n_1728),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1736),
.B(n_1716),
.Y(n_1759)
);

NAND2x1p5_ASAP7_75t_L g1760 ( 
.A(n_1735),
.B(n_1695),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1738),
.A2(n_1725),
.B1(n_1719),
.B2(n_1695),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1743),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1744),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1754),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1741),
.B(n_1728),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1755),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1740),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1733),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1737),
.B(n_1719),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1733),
.B(n_1704),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1742),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1750),
.A2(n_1695),
.B(n_1702),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1745),
.B(n_1748),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1753),
.B(n_1697),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1747),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1756),
.A2(n_1739),
.B1(n_1732),
.B2(n_1751),
.C(n_1749),
.Y(n_1776)
);

XNOR2xp5_ASAP7_75t_L g1777 ( 
.A(n_1767),
.B(n_1749),
.Y(n_1777)
);

OAI21xp33_ASAP7_75t_L g1778 ( 
.A1(n_1759),
.A2(n_1773),
.B(n_1761),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1768),
.B(n_1730),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1775),
.Y(n_1780)
);

OAI21xp33_ASAP7_75t_L g1781 ( 
.A1(n_1774),
.A2(n_1725),
.B(n_1719),
.Y(n_1781)
);

O2A1O1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1771),
.A2(n_1747),
.B(n_1704),
.C(n_1697),
.Y(n_1782)
);

AOI211x1_ASAP7_75t_SL g1783 ( 
.A1(n_1772),
.A2(n_1746),
.B(n_1704),
.C(n_1697),
.Y(n_1783)
);

AOI21xp33_ASAP7_75t_L g1784 ( 
.A1(n_1757),
.A2(n_1747),
.B(n_1697),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1769),
.B(n_1719),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1770),
.B(n_1698),
.C(n_1694),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1762),
.Y(n_1787)
);

A2O1A1Ixp33_ASAP7_75t_L g1788 ( 
.A1(n_1776),
.A2(n_1771),
.B(n_1765),
.C(n_1758),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1780),
.Y(n_1789)
);

NOR3xp33_ASAP7_75t_L g1790 ( 
.A(n_1778),
.B(n_1763),
.C(n_1766),
.Y(n_1790)
);

NAND3xp33_ASAP7_75t_L g1791 ( 
.A(n_1786),
.B(n_1764),
.C(n_1762),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1777),
.B(n_1764),
.Y(n_1792)
);

NAND4xp25_ASAP7_75t_L g1793 ( 
.A(n_1779),
.B(n_1765),
.C(n_1758),
.D(n_1701),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1782),
.B(n_1701),
.C(n_1698),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1784),
.A2(n_1760),
.B(n_1701),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_SL g1796 ( 
.A(n_1783),
.B(n_1760),
.C(n_1715),
.Y(n_1796)
);

NOR2x1_ASAP7_75t_L g1797 ( 
.A(n_1787),
.B(n_1694),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1781),
.A2(n_1760),
.B1(n_1725),
.B2(n_1722),
.Y(n_1798)
);

NOR2x1_ASAP7_75t_L g1799 ( 
.A(n_1785),
.B(n_1699),
.Y(n_1799)
);

NOR2x1_ASAP7_75t_L g1800 ( 
.A(n_1791),
.B(n_1699),
.Y(n_1800)
);

AOI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1796),
.A2(n_1717),
.B(n_1715),
.C(n_1706),
.Y(n_1801)
);

INVxp67_ASAP7_75t_SL g1802 ( 
.A(n_1799),
.Y(n_1802)
);

O2A1O1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1788),
.A2(n_1729),
.B(n_1710),
.C(n_1712),
.Y(n_1803)
);

OAI21xp33_ASAP7_75t_SL g1804 ( 
.A1(n_1798),
.A2(n_1715),
.B(n_1706),
.Y(n_1804)
);

AOI211x1_ASAP7_75t_SL g1805 ( 
.A1(n_1793),
.A2(n_1714),
.B(n_1727),
.C(n_1723),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_SL g1806 ( 
.A(n_1790),
.B(n_1717),
.C(n_1706),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1800),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1802),
.A2(n_1795),
.B(n_1792),
.Y(n_1808)
);

AO22x2_ASAP7_75t_L g1809 ( 
.A1(n_1806),
.A2(n_1789),
.B1(n_1794),
.B2(n_1797),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1804),
.A2(n_1725),
.B1(n_1722),
.B2(n_1717),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1803),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1805),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1801),
.B(n_1722),
.Y(n_1813)
);

NAND4xp25_ASAP7_75t_L g1814 ( 
.A(n_1808),
.B(n_1721),
.C(n_1727),
.D(n_1714),
.Y(n_1814)
);

NAND2x1p5_ASAP7_75t_L g1815 ( 
.A(n_1807),
.B(n_1811),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1813),
.B(n_1680),
.Y(n_1816)
);

CKINVDCx12_ASAP7_75t_R g1817 ( 
.A(n_1809),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1812),
.B(n_1710),
.Y(n_1818)
);

AND3x2_ASAP7_75t_L g1819 ( 
.A(n_1809),
.B(n_1729),
.C(n_1724),
.Y(n_1819)
);

NOR3xp33_ASAP7_75t_L g1820 ( 
.A(n_1818),
.B(n_1810),
.C(n_1724),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1815),
.Y(n_1821)
);

XNOR2xp5_ASAP7_75t_L g1822 ( 
.A(n_1819),
.B(n_1389),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1821),
.Y(n_1823)
);

NAND4xp75_ASAP7_75t_L g1824 ( 
.A(n_1823),
.B(n_1817),
.C(n_1816),
.D(n_1822),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1824),
.Y(n_1825)
);

OAI21x1_ASAP7_75t_L g1826 ( 
.A1(n_1824),
.A2(n_1814),
.B(n_1820),
.Y(n_1826)
);

OAI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1825),
.A2(n_1712),
.B1(n_1723),
.B2(n_1714),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1826),
.Y(n_1828)
);

AOI31xp33_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1826),
.A3(n_1721),
.B(n_1723),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1827),
.B(n_1727),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1829),
.A2(n_1721),
.B(n_1673),
.Y(n_1831)
);

AOI222xp33_ASAP7_75t_L g1832 ( 
.A1(n_1831),
.A2(n_1830),
.B1(n_1721),
.B2(n_1670),
.C1(n_1673),
.C2(n_1687),
.Y(n_1832)
);

AOI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1670),
.B1(n_1673),
.B2(n_1692),
.C(n_1687),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1833),
.A2(n_1692),
.B1(n_1687),
.B2(n_1683),
.Y(n_1834)
);


endmodule