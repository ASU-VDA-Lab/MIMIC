module fake_jpeg_5231_n_98 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_3),
.B(n_6),
.Y(n_14)
);

BUFx12f_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_5),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_17),
.B1(n_22),
.B2(n_12),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_22),
.B1(n_12),
.B2(n_20),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_4),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_16),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_20),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_33),
.B1(n_24),
.B2(n_25),
.Y(n_41)
);

CKINVDCx9p33_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_6),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_15),
.C(n_18),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_35),
.B(n_36),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_17),
.B1(n_22),
.B2(n_12),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_32),
.B1(n_26),
.B2(n_10),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_42),
.B1(n_50),
.B2(n_23),
.Y(n_58)
);

AO22x2_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_16),
.B1(n_19),
.B2(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_48),
.Y(n_54)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_26),
.A2(n_32),
.B1(n_27),
.B2(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_26),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_64),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_67),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_26),
.B1(n_9),
.B2(n_10),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_7),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_45),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_9),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_34),
.C(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_37),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_74),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_53),
.C(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_50),
.B(n_43),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_50),
.C(n_42),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_66),
.B1(n_54),
.B2(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_58),
.B1(n_61),
.B2(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_63),
.B1(n_59),
.B2(n_61),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_72),
.C(n_60),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_69),
.B(n_75),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_55),
.B(n_85),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.C(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_38),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_82),
.A3(n_83),
.B1(n_85),
.B2(n_80),
.C1(n_75),
.C2(n_81),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_82),
.A3(n_88),
.B1(n_60),
.B2(n_55),
.C1(n_38),
.C2(n_41),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_67),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_95),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_92),
.B(n_49),
.Y(n_96)
);

NAND5xp2_ASAP7_75t_SL g98 ( 
.A(n_96),
.B(n_47),
.C(n_51),
.D(n_97),
.E(n_95),
.Y(n_98)
);


endmodule