module fake_jpeg_7154_n_239 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_10),
.B(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_28),
.Y(n_59)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_43),
.Y(n_65)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_25),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_21),
.B1(n_16),
.B2(n_15),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_61),
.B1(n_80),
.B2(n_88),
.Y(n_94)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_28),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_54),
.Y(n_97)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_59),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_15),
.C(n_29),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_87),
.C(n_85),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_43),
.B1(n_44),
.B2(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_67),
.B1(n_76),
.B2(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_14),
.B1(n_29),
.B2(n_27),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_27),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_71),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_35),
.A2(n_30),
.B(n_31),
.C(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_32),
.B(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_37),
.A2(n_18),
.B1(n_25),
.B2(n_30),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_18),
.Y(n_78)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_37),
.A2(n_25),
.B1(n_31),
.B2(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_30),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_0),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_31),
.B1(n_25),
.B2(n_17),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_34),
.B(n_31),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_40),
.A2(n_31),
.B1(n_17),
.B2(n_0),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_40),
.A2(n_26),
.B1(n_7),
.B2(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_26),
.B1(n_6),
.B2(n_2),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_58),
.B1(n_52),
.B2(n_69),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_102),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_26),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_1),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_26),
.C(n_1),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_88),
.C(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_50),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_4),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_73),
.B(n_51),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_120),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_130),
.B1(n_101),
.B2(n_105),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_80),
.Y(n_120)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_57),
.C(n_71),
.Y(n_123)
);

XNOR2x1_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_136),
.Y(n_157)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_134),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_61),
.C(n_56),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_65),
.B(n_26),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_94),
.A2(n_55),
.B1(n_82),
.B2(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_133),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_69),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_141),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_9),
.B(n_4),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_54),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_54),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_138),
.B(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_84),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_97),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_147),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_138),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_159),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_131),
.B1(n_100),
.B2(n_106),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_139),
.B1(n_121),
.B2(n_118),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_161),
.B1(n_130),
.B2(n_134),
.Y(n_171)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_102),
.B1(n_111),
.B2(n_106),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_162),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_77),
.B(n_49),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_126),
.B(n_141),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_97),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_167),
.B(n_127),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_140),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_168),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_68),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_179),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_175),
.B(n_176),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_129),
.B(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_183),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_131),
.B1(n_100),
.B2(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_151),
.B1(n_149),
.B2(n_166),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_93),
.B(n_117),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_188),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_93),
.C(n_104),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_148),
.C(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_117),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_147),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_113),
.B(n_49),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_208)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_157),
.B1(n_164),
.B2(n_161),
.C(n_153),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_201),
.A3(n_182),
.B1(n_193),
.B2(n_200),
.C1(n_181),
.C2(n_198),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_165),
.C(n_153),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_165),
.C(n_153),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_167),
.C(n_156),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_185),
.C(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_196),
.Y(n_206)
);

OAI322xp33_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_167),
.A3(n_164),
.B1(n_152),
.B2(n_154),
.C1(n_155),
.C2(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.Y(n_209)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_198),
.A2(n_176),
.B(n_188),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_206),
.B(n_191),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_212),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_213),
.C(n_195),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_197),
.B(n_180),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_177),
.A3(n_183),
.B1(n_173),
.B2(n_154),
.C1(n_72),
.C2(n_109),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_220),
.B(n_221),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_218),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_192),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_216),
.B1(n_205),
.B2(n_208),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_227),
.B1(n_162),
.B2(n_8),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_200),
.B1(n_196),
.B2(n_177),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_178),
.B1(n_1),
.B2(n_72),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_221),
.A2(n_220),
.B1(n_178),
.B2(n_218),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_230),
.C(n_231),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_224),
.B(n_178),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_232),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_162),
.B(n_8),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_6),
.B(n_9),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_229),
.A2(n_226),
.B(n_222),
.C(n_225),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_222),
.B(n_225),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.C(n_235),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_238),
.B(n_227),
.Y(n_239)
);


endmodule