module fake_aes_9212_n_710 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_710);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_710;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g79 ( .A(n_63), .Y(n_79) );
INVx1_ASAP7_75t_SL g80 ( .A(n_45), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_15), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_50), .Y(n_82) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_71), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_7), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_77), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_57), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_28), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_7), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_24), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_75), .Y(n_91) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
BUFx2_ASAP7_75t_L g93 ( .A(n_47), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_67), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_73), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_13), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_34), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_13), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_49), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_4), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_61), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_46), .Y(n_102) );
INVxp33_ASAP7_75t_L g103 ( .A(n_68), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_66), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_23), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_31), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_37), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_6), .Y(n_108) );
BUFx2_ASAP7_75t_SL g109 ( .A(n_11), .Y(n_109) );
BUFx10_ASAP7_75t_L g110 ( .A(n_18), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_5), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_12), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_56), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_60), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_20), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_59), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_16), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_41), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_74), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_22), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_44), .Y(n_122) );
INVxp33_ASAP7_75t_SL g123 ( .A(n_5), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_17), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_8), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_10), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_27), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_123), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_124), .B(n_0), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_93), .B(n_1), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_84), .B(n_3), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_90), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_103), .B(n_3), .Y(n_135) );
INVx2_ASAP7_75t_SL g136 ( .A(n_110), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_124), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_96), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_79), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_119), .B(n_4), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_79), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_102), .B(n_6), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_87), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_91), .B(n_8), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_94), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_83), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_81), .B(n_9), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_96), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_83), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_97), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_99), .Y(n_157) );
NOR2x1_ASAP7_75t_L g158 ( .A(n_101), .B(n_9), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_126), .B(n_10), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_104), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_83), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_105), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_117), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_118), .B(n_12), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_121), .Y(n_165) );
BUFx12f_ASAP7_75t_L g166 ( .A(n_110), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_92), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_92), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_123), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g170 ( .A(n_82), .B(n_43), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_92), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_136), .B(n_114), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
NOR2xp33_ASAP7_75t_SL g175 ( .A(n_166), .B(n_114), .Y(n_175) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_135), .B(n_107), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_141), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_145), .B(n_118), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_129), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_129), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_139), .B(n_125), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_141), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_151), .A2(n_113), .B1(n_111), .B2(n_98), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_151), .A2(n_100), .B1(n_108), .B2(n_109), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_145), .B(n_95), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_136), .B(n_95), .Y(n_189) );
CKINVDCx12_ASAP7_75t_R g190 ( .A(n_144), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_156), .B(n_106), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_151), .A2(n_92), .B1(n_112), .B2(n_122), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_142), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_146), .B(n_120), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_152), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_146), .B(n_120), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_142), .B(n_82), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_159), .A2(n_112), .B1(n_115), .B2(n_106), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_159), .A2(n_112), .B1(n_115), .B2(n_107), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
INVx5_ASAP7_75t_L g203 ( .A(n_150), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_135), .B(n_86), .Y(n_204) );
BUFx4f_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_149), .B(n_86), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_144), .B(n_85), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_142), .B(n_85), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_149), .B(n_116), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_134), .Y(n_212) );
BUFx4f_ASAP7_75t_L g213 ( .A(n_155), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_147), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_163), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_163), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_155), .B(n_160), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_160), .B(n_80), .Y(n_218) );
OR2x6_ASAP7_75t_L g219 ( .A(n_131), .B(n_112), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_165), .B(n_88), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_137), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_130), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_165), .B(n_88), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g225 ( .A1(n_128), .A2(n_14), .B1(n_17), .B2(n_18), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_150), .Y(n_226) );
OR2x2_ASAP7_75t_L g227 ( .A(n_132), .B(n_157), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_130), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_147), .B(n_21), .Y(n_229) );
INVx5_ASAP7_75t_L g230 ( .A(n_150), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_157), .B(n_25), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_137), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_147), .B(n_26), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g235 ( .A(n_170), .B(n_29), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_162), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_137), .Y(n_237) );
NOR2x2_ASAP7_75t_L g238 ( .A(n_219), .B(n_128), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_237), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_191), .A2(n_148), .B(n_158), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g241 ( .A(n_197), .B(n_169), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_227), .B(n_162), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_215), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_227), .B(n_158), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_213), .B(n_138), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_190), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_205), .A2(n_138), .B1(n_169), .B2(n_171), .Y(n_247) );
NOR2xp33_ASAP7_75t_SL g248 ( .A(n_235), .B(n_130), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_237), .Y(n_249) );
OAI22xp5_ASAP7_75t_SL g250 ( .A1(n_190), .A2(n_168), .B1(n_167), .B2(n_171), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_176), .A2(n_167), .B1(n_168), .B2(n_133), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_213), .B(n_168), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_188), .B(n_167), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_195), .B(n_154), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
AND3x1_ASAP7_75t_L g256 ( .A(n_175), .B(n_154), .C(n_143), .Y(n_256) );
OAI22xp33_ASAP7_75t_L g257 ( .A1(n_197), .A2(n_154), .B1(n_143), .B2(n_140), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_206), .B(n_143), .Y(n_258) );
OR2x6_ASAP7_75t_L g259 ( .A(n_181), .B(n_140), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_216), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_198), .B(n_140), .Y(n_261) );
NOR2x1p5_ASAP7_75t_L g262 ( .A(n_181), .B(n_133), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_176), .A2(n_133), .B1(n_153), .B2(n_150), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_204), .B(n_30), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_204), .B(n_32), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_234), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_236), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_222), .Y(n_269) );
INVx8_ASAP7_75t_L g270 ( .A(n_219), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_189), .B(n_33), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_220), .B(n_161), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_207), .B(n_35), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_214), .Y(n_274) );
NAND2xp33_ASAP7_75t_L g275 ( .A(n_172), .B(n_161), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_218), .B(n_161), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_207), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_172), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_224), .A2(n_161), .B1(n_153), .B2(n_150), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_182), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_205), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_180), .B(n_161), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_182), .Y(n_283) );
NOR3x1_ASAP7_75t_L g284 ( .A(n_184), .B(n_36), .C(n_38), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_192), .B(n_39), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_205), .A2(n_161), .B1(n_153), .B2(n_48), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_186), .A2(n_153), .B1(n_42), .B2(n_51), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_213), .B(n_153), .Y(n_288) );
NAND3xp33_ASAP7_75t_SL g289 ( .A(n_200), .B(n_40), .C(n_52), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_183), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_183), .Y(n_291) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_214), .Y(n_292) );
AOI22xp33_ASAP7_75t_SL g293 ( .A1(n_221), .A2(n_153), .B1(n_54), .B2(n_55), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_174), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g295 ( .A1(n_194), .A2(n_53), .B1(n_58), .B2(n_62), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_221), .B(n_64), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_194), .A2(n_65), .B1(n_69), .B2(n_70), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_214), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_194), .B(n_78), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_196), .B(n_72), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_196), .B(n_76), .Y(n_301) );
BUFx4f_ASAP7_75t_L g302 ( .A(n_219), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_196), .B(n_187), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_174), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_202), .B(n_174), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_202), .B(n_232), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_232), .B(n_173), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_201), .B(n_202), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_SL g309 ( .A1(n_285), .A2(n_231), .B(n_193), .C(n_212), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_305), .A2(n_210), .B(n_199), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_304), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_242), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_259), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_242), .A2(n_225), .B(n_217), .C(n_184), .Y(n_314) );
NOR2x1_ASAP7_75t_L g315 ( .A(n_262), .B(n_219), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_244), .B(n_211), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_264), .A2(n_265), .B1(n_273), .B2(n_244), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_259), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_277), .B(n_241), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_264), .B(n_212), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_265), .A2(n_209), .B1(n_233), .B2(n_229), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_246), .B(n_209), .Y(n_323) );
AOI222xp33_ASAP7_75t_L g324 ( .A1(n_302), .A2(n_228), .B1(n_223), .B2(n_179), .C1(n_185), .C2(n_208), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_259), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_273), .B(n_208), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_278), .A2(n_178), .B1(n_179), .B2(n_185), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_270), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_307), .B(n_178), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_240), .B(n_223), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_240), .B(n_228), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_306), .B(n_203), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_302), .B(n_203), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_305), .A2(n_203), .B(n_230), .Y(n_335) );
O2A1O1Ixp5_ASAP7_75t_L g336 ( .A1(n_308), .A2(n_203), .B(n_230), .C(n_226), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_303), .A2(n_203), .B(n_230), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_270), .B(n_230), .Y(n_338) );
AOI22xp33_ASAP7_75t_SL g339 ( .A1(n_270), .A2(n_230), .B1(n_177), .B2(n_226), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_296), .B(n_177), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_281), .B(n_177), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_L g342 ( .A1(n_306), .A2(n_177), .B(n_226), .C(n_290), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_280), .A2(n_177), .B1(n_226), .B2(n_291), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_245), .B(n_226), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_245), .B(n_247), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_L g346 ( .A1(n_283), .A2(n_294), .B(n_260), .C(n_243), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_301), .A2(n_281), .B1(n_266), .B2(n_267), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_282), .A2(n_253), .B(n_258), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_272), .B(n_301), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_SL g350 ( .A1(n_271), .A2(n_248), .B(n_279), .C(n_295), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_276), .B(n_257), .Y(n_351) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_251), .A2(n_254), .B(n_261), .C(n_298), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_239), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_299), .A2(n_275), .B(n_292), .Y(n_354) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_274), .A2(n_263), .B(n_269), .C(n_268), .Y(n_355) );
BUFx12f_ASAP7_75t_L g356 ( .A(n_239), .Y(n_356) );
INVx4_ASAP7_75t_L g357 ( .A(n_239), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_255), .Y(n_358) );
NAND2x2_ASAP7_75t_L g359 ( .A(n_238), .B(n_284), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_250), .B(n_249), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_293), .A2(n_297), .B1(n_256), .B2(n_287), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_287), .B(n_300), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_312), .Y(n_363) );
NAND3xp33_ASAP7_75t_L g364 ( .A(n_361), .B(n_286), .C(n_248), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_359), .A2(n_289), .B1(n_252), .B2(n_288), .Y(n_365) );
AO32x2_ASAP7_75t_L g366 ( .A1(n_318), .A2(n_347), .A3(n_343), .B1(n_357), .B2(n_327), .Y(n_366) );
AO32x2_ASAP7_75t_L g367 ( .A1(n_357), .A2(n_309), .A3(n_328), .B1(n_350), .B2(n_342), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_321), .A2(n_345), .B1(n_349), .B2(n_351), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_362), .A2(n_344), .B(n_354), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_322), .A2(n_346), .B1(n_326), .B2(n_331), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_314), .B(n_320), .Y(n_371) );
AO31x2_ASAP7_75t_L g372 ( .A1(n_355), .A2(n_352), .A3(n_332), .B(n_348), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_354), .A2(n_348), .B(n_310), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_313), .B(n_325), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_314), .B(n_319), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_310), .A2(n_329), .B(n_333), .Y(n_377) );
AO31x2_ASAP7_75t_L g378 ( .A1(n_360), .A2(n_341), .A3(n_337), .B(n_335), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_316), .A2(n_340), .B(n_337), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_315), .A2(n_339), .B1(n_338), .B2(n_356), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_330), .A2(n_311), .B1(n_334), .B2(n_317), .C(n_335), .Y(n_381) );
A2O1A1Ixp33_ASAP7_75t_L g382 ( .A1(n_336), .A2(n_340), .B(n_317), .C(n_353), .Y(n_382) );
BUFx12f_ASAP7_75t_L g383 ( .A(n_358), .Y(n_383) );
AO31x2_ASAP7_75t_L g384 ( .A1(n_324), .A2(n_361), .A3(n_362), .B(n_355), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_358), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_358), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_353), .A2(n_336), .B(n_342), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_312), .B(n_221), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_336), .A2(n_342), .B(n_343), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_312), .B(n_242), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_318), .A2(n_314), .B(n_312), .C(n_277), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_312), .B(n_242), .Y(n_392) );
NAND2x1p5_ASAP7_75t_L g393 ( .A(n_328), .B(n_181), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_318), .A2(n_205), .B(n_312), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_312), .B(n_328), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_373), .A2(n_364), .B(n_369), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_389), .A2(n_387), .B(n_377), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_364), .A2(n_390), .B(n_392), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_376), .A2(n_388), .B1(n_375), .B2(n_371), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_368), .A2(n_394), .B(n_370), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_368), .B(n_363), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_395), .A2(n_380), .B1(n_374), .B2(n_381), .Y(n_403) );
NOR3xp33_ASAP7_75t_L g404 ( .A(n_391), .B(n_370), .C(n_395), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_379), .B(n_365), .C(n_382), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_384), .A2(n_386), .B(n_385), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_374), .B(n_393), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_378), .Y(n_408) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_366), .A2(n_384), .B(n_367), .C(n_378), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_384), .B(n_372), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_372), .Y(n_412) );
OA21x2_ASAP7_75t_L g413 ( .A1(n_366), .A2(n_367), .B(n_383), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_367), .A2(n_318), .B(n_373), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_366), .B(n_312), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_388), .B(n_312), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_390), .A2(n_392), .B1(n_312), .B2(n_318), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_388), .B(n_312), .Y(n_418) );
AO31x2_ASAP7_75t_L g419 ( .A1(n_373), .A2(n_370), .A3(n_369), .B(n_368), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_371), .B(n_390), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_388), .B(n_312), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_376), .B(n_221), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_373), .A2(n_369), .B(n_364), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_372), .Y(n_424) );
AND2x4_ASAP7_75t_SL g425 ( .A(n_416), .B(n_418), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_406), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_404), .B(n_408), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_408), .B(n_410), .Y(n_428) );
OA21x2_ASAP7_75t_L g429 ( .A1(n_396), .A2(n_409), .B(n_414), .Y(n_429) );
OR2x6_ASAP7_75t_L g430 ( .A(n_400), .B(n_402), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_420), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_410), .B(n_419), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_399), .B(n_402), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_412), .B(n_418), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_422), .A2(n_417), .B1(n_416), .B2(n_421), .C(n_398), .Y(n_436) );
INVx3_ASAP7_75t_L g437 ( .A(n_406), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_412), .B(n_421), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_420), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_401), .B(n_424), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_407), .Y(n_441) );
INVx4_ASAP7_75t_L g442 ( .A(n_413), .Y(n_442) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_397), .A2(n_411), .B(n_405), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_403), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_417), .B(n_405), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_419), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_401), .Y(n_447) );
AOI211xp5_ASAP7_75t_L g448 ( .A1(n_411), .A2(n_415), .B(n_401), .C(n_424), .Y(n_448) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_397), .A2(n_415), .B(n_424), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_406), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_413), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_419), .B(n_413), .Y(n_452) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_423), .A2(n_419), .B(n_413), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_419), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_423), .B(n_420), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_423), .B(n_408), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_402), .Y(n_458) );
AO31x2_ASAP7_75t_L g459 ( .A1(n_409), .A2(n_400), .A3(n_411), .B(n_410), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_402), .B(n_420), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_445), .A2(n_436), .B(n_456), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_441), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_460), .B(n_438), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_447), .Y(n_464) );
INVx4_ASAP7_75t_L g465 ( .A(n_425), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_433), .B(n_457), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_425), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_433), .B(n_457), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_426), .Y(n_469) );
NAND3xp33_ASAP7_75t_SL g470 ( .A(n_436), .B(n_444), .C(n_445), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_428), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_433), .B(n_455), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_428), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_434), .B(n_460), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_447), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_426), .Y(n_476) );
NOR2x1_ASAP7_75t_SL g477 ( .A(n_431), .B(n_439), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_441), .B(n_439), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_433), .B(n_457), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_432), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_433), .B(n_446), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_432), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_440), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_446), .B(n_455), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_435), .B(n_438), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_431), .A2(n_439), .B1(n_425), .B2(n_434), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_431), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_440), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_460), .B(n_438), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_450), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_450), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_446), .B(n_455), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_435), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_452), .B(n_435), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_454), .B(n_427), .Y(n_499) );
BUFx3_ASAP7_75t_L g500 ( .A(n_437), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_452), .B(n_430), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_458), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_452), .B(n_430), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_430), .B(n_453), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_465), .A2(n_434), .B1(n_458), .B2(n_456), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_476), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_496), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_491), .B(n_427), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_497), .B(n_427), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_497), .B(n_466), .Y(n_511) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_470), .B(n_427), .C(n_448), .D(n_442), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_470), .B(n_442), .C(n_427), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_486), .B(n_459), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_465), .B(n_448), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_497), .B(n_459), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_466), .B(n_459), .Y(n_517) );
NOR2xp33_ASAP7_75t_R g518 ( .A(n_462), .B(n_442), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_478), .B(n_442), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_496), .B(n_459), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_467), .Y(n_521) );
OR2x6_ASAP7_75t_L g522 ( .A(n_465), .B(n_430), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_477), .A2(n_430), .B(n_429), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_486), .B(n_459), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_469), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_463), .B(n_459), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_466), .B(n_459), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_492), .Y(n_528) );
INVx2_ASAP7_75t_SL g529 ( .A(n_467), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_468), .B(n_459), .Y(n_530) );
INVx11_ASAP7_75t_L g531 ( .A(n_465), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_492), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_463), .B(n_453), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_468), .B(n_453), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_463), .B(n_453), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_499), .B(n_442), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_502), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_502), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_499), .B(n_430), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_468), .B(n_430), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_493), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_493), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_464), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_479), .B(n_429), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_474), .B(n_451), .Y(n_545) );
BUFx3_ASAP7_75t_L g546 ( .A(n_467), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_479), .B(n_429), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_490), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_479), .B(n_429), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_477), .Y(n_550) );
INVx4_ASAP7_75t_L g551 ( .A(n_489), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_481), .B(n_429), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_489), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_481), .B(n_443), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_475), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_501), .B(n_443), .Y(n_556) );
NAND2xp33_ASAP7_75t_R g557 ( .A(n_487), .B(n_443), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_501), .B(n_449), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_509), .A2(n_488), .B1(n_474), .B2(n_506), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_528), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_511), .B(n_472), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_511), .B(n_489), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_528), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_512), .B(n_461), .C(n_487), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_551), .B(n_499), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_532), .Y(n_566) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_525), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_510), .B(n_472), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_508), .B(n_461), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_532), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_516), .B(n_483), .Y(n_571) );
INVxp33_ASAP7_75t_L g572 ( .A(n_518), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_514), .B(n_482), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_537), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_553), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_537), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_538), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_513), .B(n_488), .C(n_504), .D(n_485), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_516), .B(n_483), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_533), .B(n_482), .Y(n_580) );
NAND2x1_ASAP7_75t_L g581 ( .A(n_551), .B(n_494), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_538), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_535), .B(n_480), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_510), .B(n_472), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_534), .B(n_480), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_534), .B(n_476), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_524), .B(n_484), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_553), .B(n_494), .Y(n_588) );
AOI32xp33_ASAP7_75t_L g589 ( .A1(n_521), .A2(n_501), .A3(n_503), .B1(n_472), .B2(n_504), .Y(n_589) );
NAND4xp25_ASAP7_75t_L g590 ( .A(n_515), .B(n_519), .C(n_523), .D(n_557), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_526), .B(n_469), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_542), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_507), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_517), .B(n_484), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_517), .B(n_485), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_548), .B(n_495), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_531), .A2(n_472), .B1(n_500), .B2(n_473), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_551), .B(n_471), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_558), .B(n_503), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_550), .A2(n_485), .B1(n_495), .B2(n_503), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_541), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_541), .B(n_494), .C(n_487), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_527), .B(n_495), .Y(n_603) );
NAND2x1_ASAP7_75t_L g604 ( .A(n_522), .B(n_494), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_525), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_543), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_555), .Y(n_607) );
AND2x6_ASAP7_75t_L g608 ( .A(n_546), .B(n_504), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_527), .B(n_473), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_530), .B(n_471), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_593), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_606), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_601), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_569), .B(n_520), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_592), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_560), .Y(n_616) );
OAI21xp33_ASAP7_75t_SL g617 ( .A1(n_590), .A2(n_531), .B(n_529), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_563), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_561), .B(n_558), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_575), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_566), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_599), .B(n_540), .Y(n_622) );
INVx3_ASAP7_75t_L g623 ( .A(n_608), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_608), .B(n_539), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_570), .Y(n_625) );
NAND2xp33_ASAP7_75t_L g626 ( .A(n_608), .B(n_529), .Y(n_626) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_581), .B(n_546), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_567), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_571), .B(n_530), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_574), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_576), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_562), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_579), .B(n_549), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_564), .A2(n_522), .B1(n_539), .B2(n_540), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_585), .B(n_549), .Y(n_635) );
NAND2xp33_ASAP7_75t_L g636 ( .A(n_608), .B(n_498), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_590), .B(n_545), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_577), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_586), .B(n_544), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_573), .B(n_554), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_582), .Y(n_641) );
NOR2x1p5_ASAP7_75t_SL g642 ( .A(n_605), .B(n_505), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_607), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_580), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_587), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_583), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_609), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_610), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_637), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_614), .B(n_595), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_613), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_619), .B(n_556), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_637), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_631), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_631), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_622), .B(n_556), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_641), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_611), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_641), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_615), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_646), .B(n_547), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_617), .A2(n_589), .B1(n_578), .B2(n_559), .C(n_600), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_623), .B(n_565), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_616), .Y(n_664) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_623), .A2(n_565), .B1(n_597), .B2(n_598), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_614), .B(n_603), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_624), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_618), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_621), .Y(n_669) );
OAI21xp5_ASAP7_75t_SL g670 ( .A1(n_634), .A2(n_572), .B(n_600), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_612), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_649), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_665), .B(n_627), .Y(n_673) );
XNOR2x1_ASAP7_75t_L g674 ( .A(n_667), .B(n_627), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_650), .B(n_640), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_662), .A2(n_626), .B(n_636), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_651), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_653), .A2(n_644), .B1(n_647), .B2(n_648), .C(n_620), .Y(n_678) );
AOI322xp5_ASAP7_75t_L g679 ( .A1(n_666), .A2(n_634), .A3(n_629), .B1(n_632), .B2(n_626), .C1(n_633), .C2(n_635), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_670), .A2(n_636), .B1(n_628), .B2(n_559), .C(n_604), .Y(n_680) );
AOI322xp5_ASAP7_75t_L g681 ( .A1(n_661), .A2(n_639), .A3(n_624), .B1(n_645), .B2(n_594), .C1(n_584), .C2(n_568), .Y(n_681) );
NAND5xp2_ASAP7_75t_L g682 ( .A(n_658), .B(n_602), .C(n_552), .D(n_547), .E(n_544), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_661), .B(n_643), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_667), .B(n_624), .Y(n_684) );
AOI21xp33_ASAP7_75t_R g685 ( .A1(n_667), .A2(n_630), .B(n_625), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_683), .Y(n_686) );
OAI211xp5_ASAP7_75t_SL g687 ( .A1(n_680), .A2(n_660), .B(n_669), .C(n_668), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_676), .A2(n_663), .B(n_588), .C(n_664), .Y(n_688) );
OAI211xp5_ASAP7_75t_SL g689 ( .A1(n_679), .A2(n_655), .B(n_657), .C(n_659), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_672), .A2(n_673), .B(n_678), .C(n_677), .Y(n_690) );
AND2x4_ASAP7_75t_L g691 ( .A(n_684), .B(n_663), .Y(n_691) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_674), .B(n_663), .Y(n_692) );
AOI31xp33_ASAP7_75t_L g693 ( .A1(n_685), .A2(n_652), .A3(n_656), .B(n_645), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_686), .B(n_681), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_693), .B(n_671), .Y(n_695) );
NAND4xp75_ASAP7_75t_L g696 ( .A(n_692), .B(n_642), .C(n_682), .D(n_652), .Y(n_696) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_687), .B(n_682), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_688), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_694), .Y(n_699) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_698), .Y(n_700) );
NAND5xp2_ASAP7_75t_L g701 ( .A(n_696), .B(n_690), .C(n_697), .D(n_689), .E(n_695), .Y(n_701) );
OR5x1_ASAP7_75t_L g702 ( .A(n_700), .B(n_691), .C(n_675), .D(n_656), .E(n_671), .Y(n_702) );
XNOR2xp5_ASAP7_75t_L g703 ( .A(n_699), .B(n_655), .Y(n_703) );
INVx4_ASAP7_75t_L g704 ( .A(n_702), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_703), .B(n_699), .C(n_701), .Y(n_705) );
OAI22x1_ASAP7_75t_L g706 ( .A1(n_704), .A2(n_654), .B1(n_598), .B2(n_638), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_706), .A2(n_705), .B(n_591), .Y(n_707) );
OAI21xp5_ASAP7_75t_SL g708 ( .A1(n_707), .A2(n_596), .B(n_539), .Y(n_708) );
INVxp33_ASAP7_75t_L g709 ( .A(n_708), .Y(n_709) );
OAI21xp33_ASAP7_75t_L g710 ( .A1(n_709), .A2(n_552), .B(n_536), .Y(n_710) );
endmodule