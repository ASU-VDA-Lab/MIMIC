module fake_jpeg_2845_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_45),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_1),
.C(n_2),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_62),
.C(n_70),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_29),
.B1(n_32),
.B2(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_33),
.B1(n_27),
.B2(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_18),
.B(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_55),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_18),
.B(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_15),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_14),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_1),
.C(n_2),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_1),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_3),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_42),
.B1(n_39),
.B2(n_23),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_23),
.B1(n_36),
.B2(n_28),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_80),
.Y(n_122)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_79),
.Y(n_136)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_84),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_36),
.B1(n_37),
.B2(n_28),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_37),
.B1(n_19),
.B2(n_26),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_109),
.Y(n_128)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

CKINVDCx9p33_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_33),
.B1(n_27),
.B2(n_22),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_20),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_114),
.Y(n_130)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_20),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_34),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_22),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_21),
.B(n_63),
.C(n_64),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_117),
.B(n_123),
.C(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_71),
.B(n_21),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_11),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_12),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_13),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_91),
.A2(n_66),
.B1(n_17),
.B2(n_7),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_143),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_72),
.B(n_3),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_73),
.C(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_4),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_9),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_82),
.Y(n_161)
);

NOR2xp67_ASAP7_75t_R g186 ( 
.A(n_147),
.B(n_82),
.Y(n_186)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_157),
.Y(n_171)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_88),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_159),
.C(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_130),
.B1(n_117),
.B2(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_160),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_87),
.C(n_107),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_92),
.B1(n_113),
.B2(n_75),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_161),
.B(n_167),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_128),
.Y(n_177)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_107),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_104),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_124),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_125),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_184),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_134),
.B1(n_113),
.B2(n_75),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_183),
.B1(n_158),
.B2(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_132),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_132),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_187),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_86),
.B1(n_112),
.B2(n_135),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_116),
.B(n_126),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_185),
.A2(n_186),
.B(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NAND2x1p5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_203),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_180),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_194),
.A2(n_181),
.B(n_155),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_159),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_176),
.C(n_179),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_202),
.B1(n_169),
.B2(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_201),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_157),
.Y(n_199)
);

OAI322xp33_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_177),
.A3(n_186),
.B1(n_181),
.B2(n_185),
.C1(n_155),
.C2(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_146),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_162),
.B1(n_156),
.B2(n_149),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_146),
.A3(n_164),
.B1(n_119),
.B2(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_190),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_139),
.C(n_124),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_191),
.B(n_172),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_216),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_86),
.B1(n_112),
.B2(n_151),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_165),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_116),
.B(n_139),
.C(n_135),
.D(n_101),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_215),
.B(n_203),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_199),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_224),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_197),
.B1(n_195),
.B2(n_192),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_222),
.B1(n_207),
.B2(n_214),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_212),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_208),
.C(n_210),
.Y(n_227)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_230),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_226),
.B(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_231),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_213),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_207),
.B(n_210),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_233),
.B(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_218),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_237),
.Y(n_243)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_229),
.Y(n_237)
);

AOI21x1_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_225),
.B(n_224),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_236),
.B1(n_222),
.B2(n_219),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_239),
.A2(n_238),
.B(n_240),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_244),
.B(n_240),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_247),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_223),
.B(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_243),
.B(n_227),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_230),
.B(n_217),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_251),
.B(n_76),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_124),
.C(n_76),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_101),
.Y(n_253)
);


endmodule