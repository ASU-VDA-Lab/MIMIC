module real_jpeg_9692_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_1),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_48),
.Y(n_116)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_23),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_8),
.A2(n_22),
.B(n_23),
.C(n_59),
.D(n_61),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_76),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g95 ( 
.A1(n_8),
.A2(n_26),
.B(n_50),
.C(n_86),
.D(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_8),
.B(n_26),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_8),
.B(n_60),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_8),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_44),
.B(n_111),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_42),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_11),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_91),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_64),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_17),
.B(n_64),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.C(n_58),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_18),
.A2(n_19),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_31),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.C(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_60)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_27),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_51),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_38),
.B(n_40),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_32),
.A2(n_38),
.B1(n_44),
.B2(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_33),
.B(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_33),
.B(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_38),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_34),
.A2(n_53),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_38),
.A2(n_40),
.B(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_38),
.B(n_123),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_39),
.B(n_41),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_39),
.A2(n_43),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_44),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_45),
.A2(n_46),
.B1(n_58),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_47),
.A2(n_57),
.B(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_55),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_50),
.B(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_57),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_58),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_68),
.B(n_69),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_82),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_81),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_75),
.B1(n_79),
.B2(n_80),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_75),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_84),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_132),
.B(n_138),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_112),
.B(n_131),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_97),
.B1(n_98),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_106),
.C(n_109),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_120),
.B(n_130),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_118),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_125),
.B(n_129),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_133),
.B(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);


endmodule