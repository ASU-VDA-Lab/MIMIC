module fake_jpeg_22916_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_48),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_0),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_27),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_1),
.CON(n_46),
.SN(n_46)
);

OAI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_34),
.B(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_37),
.B1(n_36),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_61),
.B1(n_79),
.B2(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_37),
.B1(n_34),
.B2(n_28),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_53),
.A2(n_84),
.B1(n_85),
.B2(n_47),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_34),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_56),
.A2(n_70),
.B(n_33),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_37),
.B1(n_27),
.B2(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_62),
.B(n_69),
.Y(n_116)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_64),
.Y(n_101)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_32),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_27),
.B1(n_19),
.B2(n_24),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_38),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_30),
.B1(n_26),
.B2(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_38),
.B1(n_26),
.B2(n_30),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_39),
.A2(n_17),
.B1(n_18),
.B2(n_33),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_89),
.B(n_118),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_95),
.Y(n_131)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_25),
.B1(n_22),
.B2(n_35),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_97),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_105),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_24),
.B1(n_35),
.B2(n_43),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_49),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_49),
.B1(n_44),
.B2(n_47),
.Y(n_106)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_1),
.A3(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_56),
.B(n_44),
.CI(n_49),
.CON(n_108),
.SN(n_108)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_72),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_89),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_53),
.A2(n_43),
.B1(n_47),
.B2(n_21),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_59),
.A2(n_33),
.B1(n_18),
.B2(n_17),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_81),
.B1(n_17),
.B2(n_18),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_55),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_39),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_121),
.B(n_21),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_33),
.B1(n_18),
.B2(n_17),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_21),
.B1(n_29),
.B2(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_93),
.B1(n_115),
.B2(n_104),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_134),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_54),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_157),
.C(n_107),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_132),
.B(n_113),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_73),
.CI(n_83),
.CON(n_130),
.SN(n_130)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_130),
.B(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_137),
.Y(n_164)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_88),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_142),
.Y(n_192)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_78),
.B1(n_86),
.B2(n_74),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_149),
.B1(n_152),
.B2(n_155),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_58),
.B1(n_29),
.B2(n_1),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_58),
.Y(n_151)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_90),
.A2(n_29),
.B1(n_1),
.B2(n_3),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_109),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_159),
.B1(n_142),
.B2(n_125),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_108),
.C(n_104),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_7),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_158)
);

XOR2x2_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_11),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_11),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_156),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_108),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_161),
.A2(n_173),
.B(n_176),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_167),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_127),
.B(n_116),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_137),
.B1(n_147),
.B2(n_139),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_171),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_106),
.B1(n_93),
.B2(n_115),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_155),
.B1(n_94),
.B2(n_130),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_172),
.B(n_174),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_132),
.B(n_143),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_177),
.B(n_181),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_129),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_16),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

OA21x2_ASAP7_75t_SL g208 ( 
.A1(n_182),
.A2(n_12),
.B(n_13),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_107),
.C(n_120),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_120),
.C(n_106),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_106),
.C(n_102),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_189),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_134),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_150),
.A2(n_102),
.B(n_94),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_13),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_153),
.B(n_130),
.C(n_158),
.D(n_152),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_196),
.A2(n_204),
.B(n_210),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_197),
.A2(n_205),
.B1(n_163),
.B2(n_180),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_164),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_198),
.B(n_201),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_189),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_211),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_174),
.A2(n_154),
.B1(n_124),
.B2(n_138),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_193),
.A2(n_123),
.B1(n_138),
.B2(n_14),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_175),
.B1(n_181),
.B2(n_160),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_208),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_13),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_220),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_190),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_222),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_175),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_15),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_173),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_234),
.C(n_202),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_214),
.B(n_183),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_228),
.B(n_236),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_176),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_235),
.B1(n_245),
.B2(n_246),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_221),
.A2(n_193),
.B1(n_170),
.B2(n_187),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_237),
.B1(n_241),
.B2(n_242),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_161),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_182),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_211),
.A2(n_169),
.B1(n_194),
.B2(n_161),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_171),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_239),
.B(n_247),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_205),
.A2(n_178),
.B1(n_186),
.B2(n_167),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_227),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_252),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_261),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_207),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_264),
.C(n_265),
.Y(n_270)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_232),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_267),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_209),
.B1(n_207),
.B2(n_217),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_225),
.B1(n_228),
.B2(n_224),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_202),
.C(n_200),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_230),
.C(n_243),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_200),
.C(n_196),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_268),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_241),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_220),
.C(n_199),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_199),
.C(n_204),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_272),
.A2(n_277),
.B(n_282),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_201),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_273),
.B(n_284),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_229),
.CI(n_226),
.CON(n_275),
.SN(n_275)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_233),
.B(n_229),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_278),
.A2(n_280),
.B(n_286),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_229),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_283),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_268),
.B(n_239),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_258),
.B(n_236),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_251),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_287),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_246),
.B(n_249),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_263),
.B1(n_258),
.B2(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_295),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_280),
.B(n_270),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_294),
.A2(n_279),
.B(n_281),
.Y(n_303)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_224),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_250),
.C(n_252),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_271),
.C(n_281),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_225),
.B1(n_253),
.B2(n_245),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_301),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_215),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_309),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_304),
.C(n_300),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_271),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_290),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_275),
.B(n_210),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_292),
.B(n_276),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_318),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_301),
.B(n_288),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_313),
.A2(n_315),
.B(n_308),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_195),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_310),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_319),
.C(n_307),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_292),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_290),
.C(n_293),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_323),
.B(n_317),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_327),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_324),
.A2(n_313),
.B(n_311),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_SL g329 ( 
.A(n_326),
.B(n_321),
.C(n_306),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_309),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_195),
.Y(n_332)
);

AO31x2_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_216),
.A3(n_247),
.B(n_203),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_15),
.C(n_16),
.Y(n_334)
);


endmodule