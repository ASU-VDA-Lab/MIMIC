module real_jpeg_26060_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_36),
.B1(n_93),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_1),
.A2(n_36),
.B1(n_53),
.B2(n_54),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_2),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_78),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_2),
.B(n_54),
.C(n_64),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_31),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_2),
.A2(n_81),
.B1(n_163),
.B2(n_170),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_69),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_69),
.Y(n_153)
);

INVx8_ASAP7_75t_SL g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_8),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_9),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_58),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_12),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_73),
.Y(n_83)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_15),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_126),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_19),
.B(n_87),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_60),
.C(n_74),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_20),
.A2(n_21),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_22),
.B(n_41),
.C(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_23),
.A2(n_37),
.B1(n_39),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_24),
.A2(n_31),
.B1(n_35),
.B2(n_77),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_27),
.A2(n_29),
.A3(n_33),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_29),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g77 ( 
.A(n_28),
.B(n_78),
.CON(n_77),
.SN(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_28),
.A2(n_45),
.B(n_91),
.C(n_94),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_29),
.B(n_44),
.C(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_32),
.A2(n_33),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_33),
.B(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_44),
.A2(n_45),
.B1(n_93),
.B2(n_109),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B(n_56),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_53),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_59),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_51),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_54),
.B1(n_64),
.B2(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_53),
.B(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_59),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_60),
.A2(n_61),
.B1(n_74),
.B2(n_75),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_68),
.B(n_70),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_62),
.A2(n_72),
.B(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_68),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_62),
.A2(n_133),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_62),
.A2(n_132),
.B1(n_133),
.B2(n_143),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_67),
.B(n_78),
.Y(n_168)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_76),
.B(n_80),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_78),
.B(n_171),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_84),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_81),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_81),
.A2(n_160),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_86),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_103),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_102),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_116),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_110),
.B2(n_113),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_137),
.B(n_185),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_128),
.B(n_134),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.C(n_131),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_130),
.B(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_180),
.B(n_184),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_156),
.B(n_179),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_140),
.B(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_144),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_151),
.C(n_152),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_166),
.B(n_178),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_165),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_165),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_173),
.B(n_177),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_181),
.B(n_182),
.Y(n_184)
);


endmodule