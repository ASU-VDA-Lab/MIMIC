module real_jpeg_18375_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_0),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_22),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_2),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_2),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_2),
.A2(n_87),
.B1(n_170),
.B2(n_176),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_2),
.A2(n_87),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_2),
.A2(n_87),
.B1(n_300),
.B2(n_303),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_4),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_5),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_5),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g454 ( 
.A(n_5),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_6),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_6),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_6),
.A2(n_270),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_6),
.A2(n_270),
.B1(n_472),
.B2(n_474),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g528 ( 
.A1(n_6),
.A2(n_270),
.B1(n_529),
.B2(n_534),
.Y(n_528)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_7),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_7),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_7),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_8),
.Y(n_151)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_8),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_8),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_8),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_8),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_8),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_9),
.A2(n_42),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_9),
.A2(n_42),
.B1(n_158),
.B2(n_162),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_9),
.A2(n_42),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_10),
.A2(n_72),
.B1(n_340),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_10),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_10),
.A2(n_370),
.B1(n_398),
.B2(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_10),
.A2(n_370),
.B1(n_462),
.B2(n_467),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_10),
.A2(n_370),
.B1(n_504),
.B2(n_505),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g334 ( 
.A1(n_12),
.A2(n_335),
.A3(n_339),
.B1(n_341),
.B2(n_346),
.Y(n_334)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_12),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_12),
.A2(n_89),
.B1(n_345),
.B2(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_12),
.B(n_27),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_12),
.B(n_119),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_12),
.B(n_513),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_12),
.B(n_138),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_12),
.A2(n_172),
.B1(n_345),
.B2(n_537),
.Y(n_536)
);

OAI32xp33_ASAP7_75t_L g540 ( 
.A1(n_12),
.A2(n_541),
.A3(n_543),
.B1(n_544),
.B2(n_548),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_14),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_14),
.A2(n_77),
.B1(n_191),
.B2(n_195),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_14),
.A2(n_77),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_14),
.A2(n_77),
.B1(n_353),
.B2(n_359),
.Y(n_352)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_15),
.Y(n_140)
);

BUFx4f_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_15),
.Y(n_218)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_15),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_16),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_16),
.A2(n_52),
.B1(n_95),
.B2(n_100),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_16),
.A2(n_52),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_16),
.A2(n_52),
.B1(n_253),
.B2(n_256),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_584),
.Y(n_22)
);

OAI221xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_62),
.B1(n_65),
.B2(n_289),
.C(n_578),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_24),
.B(n_62),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_25),
.B(n_282),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_25),
.B(n_282),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_47),
.Y(n_25)
);

OAI21x1_ASAP7_75t_SL g266 ( 
.A1(n_26),
.A2(n_54),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

OR2x6_ASAP7_75t_L g54 ( 
.A(n_27),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_27),
.B(n_48),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_27),
.A2(n_53),
.B1(n_368),
.B2(n_371),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_33),
.Y(n_175)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_33),
.Y(n_411)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_36),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_37),
.Y(n_179)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_37),
.Y(n_332)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_44),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_44),
.Y(n_317)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21x1_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_63),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_63),
.B(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_63),
.B1(n_71),
.B2(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_54),
.A2(n_64),
.B(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_54),
.A2(n_81),
.B(n_238),
.Y(n_283)
);

OAI22x1_ASAP7_75t_SL g313 ( 
.A1(n_54),
.A2(n_63),
.B1(n_267),
.B2(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_54),
.A2(n_63),
.B1(n_369),
.B2(n_390),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_59),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_61),
.Y(n_350)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_279),
.C(n_288),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_239),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_67),
.A2(n_580),
.B(n_581),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_182),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g581 ( 
.A(n_68),
.B(n_182),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_167),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_78),
.B1(n_79),
.B2(n_166),
.Y(n_69)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_70),
.B(n_137),
.C(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_70),
.A2(n_166),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_70),
.B(n_167),
.C(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_74),
.Y(n_348)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_75),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_79),
.Y(n_281)
);

XNOR2x1_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.Y(n_79)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_80),
.Y(n_287)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_137),
.B2(n_165),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_92),
.B(n_165),
.C(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_103),
.B(n_130),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_94),
.B(n_119),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_94),
.Y(n_274)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

AOI21x1_ASAP7_75t_L g168 ( 
.A1(n_103),
.A2(n_169),
.B(n_180),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_103),
.A2(n_119),
.B1(n_169),
.B2(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_103),
.A2(n_119),
.B(n_285),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_103),
.A2(n_130),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_104),
.A2(n_131),
.B1(n_190),
.B2(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_104),
.A2(n_132),
.B(n_181),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_104),
.A2(n_131),
.B1(n_326),
.B2(n_394),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_L g407 ( 
.A1(n_104),
.A2(n_131),
.B1(n_394),
.B2(n_408),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_104),
.A2(n_131),
.B1(n_408),
.B2(n_536),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_119),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_111),
.B1(n_113),
.B2(n_116),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_111),
.Y(n_327)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

AO22x2_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_119)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_121),
.Y(n_460)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_122),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_123),
.Y(n_481)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_128),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_132),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_134),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_168),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_147),
.B(n_156),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_138),
.B(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_138),
.B(n_261),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_138),
.A2(n_147),
.B1(n_459),
.B2(n_461),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_138),
.A2(n_147),
.B1(n_461),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_157),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_139),
.A2(n_227),
.B1(n_234),
.B2(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_139),
.A2(n_234),
.B1(n_527),
.B2(n_528),
.Y(n_526)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_145),
.Y(n_139)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_140),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_140),
.Y(n_258)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_140),
.Y(n_302)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_140),
.Y(n_473)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_140),
.Y(n_511)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_141),
.Y(n_448)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_144),
.Y(n_305)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_144),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_147),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_147),
.A2(n_204),
.B(n_564),
.Y(n_563)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_151),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_155),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_157),
.A2(n_234),
.B(n_235),
.Y(n_388)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_176),
.Y(n_398)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_179),
.Y(n_542)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_205),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_183),
.A2(n_186),
.B1(n_187),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_183),
.Y(n_278)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g244 ( 
.A1(n_187),
.A2(n_188),
.B(n_196),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_198),
.B(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_203),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_205),
.A2(n_206),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_224),
.B(n_236),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_208),
.B1(n_236),
.B2(n_237),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_207),
.A2(n_208),
.B1(n_226),
.B2(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_214),
.B(n_221),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_212),
.Y(n_309)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_213),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_214),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_214),
.A2(n_471),
.B(n_477),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_214),
.A2(n_345),
.B1(n_502),
.B2(n_503),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_214),
.A2(n_490),
.B1(n_503),
.B2(n_517),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_216),
.Y(n_505)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_217),
.Y(n_476)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_218),
.Y(n_446)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_221),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_226),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_235),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_233),
.Y(n_468)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_275),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_240),
.B(n_275),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.C(n_245),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_241),
.Y(n_428)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_245),
.B(n_427),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_266),
.C(n_272),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g376 ( 
.A(n_246),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_259),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_247),
.B(n_259),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_248),
.Y(n_477)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_251),
.A2(n_352),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_266),
.B(n_273),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_268),
.A2(n_315),
.B1(n_316),
.B2(n_318),
.Y(n_314)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_269),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g578 ( 
.A1(n_279),
.A2(n_288),
.B(n_579),
.C(n_582),
.D(n_583),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_280),
.B(n_282),
.Y(n_582)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.CI(n_286),
.CON(n_282),
.SN(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_430),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_381),
.B(n_422),
.C(n_423),
.D(n_429),
.Y(n_291)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_292),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_372),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_293),
.B(n_372),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_320),
.C(n_322),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_294),
.A2(n_295),
.B1(n_320),
.B2(n_321),
.Y(n_383)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_312),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_296),
.B(n_313),
.C(n_319),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_310),
.Y(n_296)
);

XOR2x2_ASAP7_75t_L g399 ( 
.A(n_297),
.B(n_310),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B(n_306),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_298),
.A2(n_299),
.B1(n_352),
.B2(n_363),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_298),
.A2(n_489),
.B1(n_494),
.B2(n_495),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_298),
.A2(n_306),
.B(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_319),
.Y(n_312)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_315),
.A2(n_318),
.B1(n_395),
.B2(n_398),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_315),
.A2(n_318),
.B1(n_481),
.B2(n_482),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_315),
.A2(n_318),
.B1(n_455),
.B2(n_491),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_322),
.B(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_333),
.C(n_367),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_367),
.Y(n_386)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_330),
.Y(n_538)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_331),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_332),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_333),
.B(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_351),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_334),
.B(n_351),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_345),
.B(n_450),
.Y(n_449)
);

OAI21xp33_ASAP7_75t_SL g459 ( 
.A1(n_345),
.A2(n_449),
.B(n_460),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_345),
.B(n_545),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_358),
.Y(n_362)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_366),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_373),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_374),
.B(n_376),
.C(n_378),
.Y(n_425)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.C(n_400),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_384),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.C(n_399),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_399),
.Y(n_421)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.C(n_393),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_393),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_389),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx2_ASAP7_75t_SL g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_420),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_420),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.C(n_406),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_402),
.B(n_575),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_404),
.A2(n_405),
.B1(n_406),
.B2(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_406),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_412),
.C(n_414),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g566 ( 
.A(n_407),
.B(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_412),
.A2(n_413),
.B1(n_415),
.B2(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_415),
.Y(n_568)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

INVx6_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NOR3xp33_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_432),
.C(n_435),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_426),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_436),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_571),
.B(n_577),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_558),
.B(n_570),
.Y(n_437)
);

OAI21x1_ASAP7_75t_SL g438 ( 
.A1(n_439),
.A2(n_522),
.B(n_557),
.Y(n_438)
);

AOI21x1_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_486),
.B(n_521),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_469),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_441),
.B(n_469),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_457),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_442),
.A2(n_457),
.B1(n_458),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_442),
.Y(n_498)
);

OAI32xp33_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_444),
.A3(n_447),
.B1(n_449),
.B2(n_452),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_446),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_451),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_466),
.Y(n_547)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_478),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_470),
.B(n_479),
.C(n_485),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_471),
.Y(n_494)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_485),
.Y(n_478)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_480),
.Y(n_527)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_487),
.A2(n_499),
.B(n_520),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_497),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_497),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_515),
.B(n_519),
.Y(n_499)
);

NOR2x1_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_506),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_512),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_516),
.B(n_518),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_516),
.B(n_518),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_524),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_523),
.B(n_524),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_539),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_535),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_526),
.B(n_535),
.C(n_539),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_528),
.Y(n_564)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_532),
.Y(n_543)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_555),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_540),
.B(n_555),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_552),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_560),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_559),
.B(n_560),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_561),
.A2(n_565),
.B1(n_566),
.B2(n_569),
.Y(n_560)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_561),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_563),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_562),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_565),
.C(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_574),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_572),
.B(n_574),
.Y(n_577)
);


endmodule