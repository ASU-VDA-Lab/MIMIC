module fake_ibex_673_n_2548 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_483, n_141, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_479, n_225, n_360, n_272, n_23, n_468, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_482, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_460, n_476, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2548);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_141;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_479;
input n_225;
input n_360;
input n_272;
input n_23;
input n_468;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_460;
input n_476;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2548;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_2475;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_2311;
wire n_1937;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_787;
wire n_523;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_646;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_553;
wire n_554;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2112;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2509;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2470;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_1831;
wire n_864;
wire n_608;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2390;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_660;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_607;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2524;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_961;
wire n_634;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_2180;
wire n_1952;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_2528;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2251;
wire n_722;
wire n_2012;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2447;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2417;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_2518;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2487;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2513;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2303;
wire n_949;
wire n_704;
wire n_2357;
wire n_2104;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2435;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_2430;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_182),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_253),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_199),
.B(n_62),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g490 ( 
.A(n_360),
.B(n_2),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_12),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_332),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_198),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_33),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_72),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_95),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_129),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_11),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_145),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_31),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_374),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_195),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_65),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_87),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_131),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_440),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_14),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_264),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_339),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_454),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_444),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_57),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_478),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_74),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_283),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_126),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_332),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_310),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_79),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_240),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_301),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_215),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_272),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_458),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_57),
.Y(n_525)
);

INVxp33_ASAP7_75t_SL g526 ( 
.A(n_174),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_15),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_128),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_65),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_288),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_24),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_471),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_25),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_315),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_29),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_L g536 ( 
.A(n_251),
.B(n_363),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_248),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_466),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_461),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_164),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_264),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_475),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_224),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_305),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_417),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_220),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_412),
.Y(n_547)
);

BUFx5_ASAP7_75t_L g548 ( 
.A(n_42),
.Y(n_548)
);

BUFx5_ASAP7_75t_L g549 ( 
.A(n_5),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_131),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_73),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_437),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_371),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_162),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_346),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_252),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_56),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_321),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_149),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_31),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_290),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_291),
.Y(n_562)
);

BUFx5_ASAP7_75t_L g563 ( 
.A(n_108),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_252),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_480),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_317),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_418),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_467),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_229),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_L g570 ( 
.A(n_316),
.B(n_368),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_233),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_256),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_393),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_66),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_379),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_288),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_80),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_396),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_14),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_226),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_269),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_10),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_150),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_477),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_276),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_468),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_250),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_479),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_325),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_389),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_470),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_274),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_12),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_221),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_465),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_193),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_421),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_338),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_256),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_55),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_413),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_30),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_432),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_202),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_270),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_349),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_346),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_198),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_154),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_369),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_287),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_84),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_280),
.Y(n_613)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_314),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_425),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_433),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_254),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_228),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_36),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_392),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_143),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_119),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_7),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_339),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_98),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_91),
.Y(n_626)
);

BUFx2_ASAP7_75t_SL g627 ( 
.A(n_20),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_17),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_67),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_403),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_453),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_187),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_11),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_455),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_430),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_410),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_303),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_184),
.Y(n_638)
);

CKINVDCx16_ASAP7_75t_R g639 ( 
.A(n_46),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_446),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_103),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_92),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_195),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_298),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_258),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_72),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_55),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_409),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_400),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_327),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_366),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_331),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_172),
.Y(n_653)
);

CKINVDCx14_ASAP7_75t_R g654 ( 
.A(n_89),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_214),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_88),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_291),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_337),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_394),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_190),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_95),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_334),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_424),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_263),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_463),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_277),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_196),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_459),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_271),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_180),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_456),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_450),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_405),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_354),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_429),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_91),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_113),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_397),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_428),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_247),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_457),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_274),
.Y(n_682)
);

INVx1_ASAP7_75t_SL g683 ( 
.A(n_485),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_476),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_245),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_352),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_88),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_431),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_141),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_338),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_351),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_462),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_185),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_139),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_64),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_90),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_353),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_216),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_87),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_46),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_401),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_284),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_101),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_483),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_8),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_190),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_21),
.Y(n_707)
);

CKINVDCx14_ASAP7_75t_R g708 ( 
.A(n_203),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_181),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_434),
.B(n_230),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_246),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_324),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_64),
.Y(n_713)
);

CKINVDCx16_ASAP7_75t_R g714 ( 
.A(n_70),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_277),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_161),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_214),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_261),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_99),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_184),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_194),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_194),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_345),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_445),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_415),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_411),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_276),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_35),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_318),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_L g730 ( 
.A(n_316),
.B(n_92),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_5),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_451),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_426),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_223),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_448),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_144),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_148),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_473),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_452),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_19),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_135),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_129),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_344),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_317),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_464),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_51),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_261),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_406),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_315),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_271),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_32),
.Y(n_751)
);

NOR2xp67_ASAP7_75t_L g752 ( 
.A(n_245),
.B(n_402),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_328),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_179),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_257),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_51),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_239),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_322),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_191),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_319),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_211),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_246),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_484),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_208),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_362),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_438),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_414),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_469),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_270),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_132),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_243),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_460),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_321),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_358),
.Y(n_774)
);

CKINVDCx11_ASAP7_75t_R g775 ( 
.A(n_62),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_427),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_37),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_L g778 ( 
.A(n_279),
.B(n_340),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_192),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_204),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_336),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_137),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_482),
.B(n_69),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_420),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_29),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_443),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_416),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_42),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_481),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_117),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_300),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_213),
.Y(n_792)
);

NOR2xp67_ASAP7_75t_L g793 ( 
.A(n_367),
.B(n_83),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_90),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_231),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_40),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_24),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_419),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_408),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_449),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_262),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_84),
.Y(n_802)
);

CKINVDCx14_ASAP7_75t_R g803 ( 
.A(n_435),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_319),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_107),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_355),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_292),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_282),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_486),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_309),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_168),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_119),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_172),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_161),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_250),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_152),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_56),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_524),
.B(n_356),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_511),
.A2(n_359),
.B(n_357),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_548),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_532),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_548),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_548),
.Y(n_823)
);

BUFx12f_ASAP7_75t_L g824 ( 
.A(n_547),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_548),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_548),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_700),
.Y(n_827)
);

OAI21x1_ASAP7_75t_L g828 ( 
.A1(n_511),
.A2(n_364),
.B(n_361),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_700),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_548),
.Y(n_830)
);

AND2x6_ASAP7_75t_L g831 ( 
.A(n_631),
.B(n_365),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_548),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_549),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_549),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_522),
.B(n_0),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_487),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_487),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_549),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_654),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_547),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_654),
.Y(n_841)
);

OA21x2_ASAP7_75t_L g842 ( 
.A1(n_684),
.A2(n_372),
.B(n_370),
.Y(n_842)
);

OA21x2_ASAP7_75t_L g843 ( 
.A1(n_684),
.A2(n_375),
.B(n_373),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_532),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_549),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_506),
.B(n_1),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_547),
.B(n_3),
.Y(n_847)
);

BUFx12f_ASAP7_75t_L g848 ( 
.A(n_775),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_708),
.Y(n_849)
);

OA21x2_ASAP7_75t_L g850 ( 
.A1(n_726),
.A2(n_377),
.B(n_376),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_549),
.Y(n_851)
);

INVx5_ASAP7_75t_L g852 ( 
.A(n_532),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_549),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_687),
.B(n_4),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_563),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_505),
.B(n_4),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_631),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_708),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_563),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_515),
.B(n_6),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_519),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_701),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_726),
.A2(n_380),
.B(n_378),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_707),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_701),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_541),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_798),
.A2(n_382),
.B(n_381),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_733),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_701),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_515),
.B(n_9),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_563),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_541),
.B(n_10),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_558),
.B(n_13),
.Y(n_873)
);

NOR2x1_ASAP7_75t_L g874 ( 
.A(n_618),
.B(n_383),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_701),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_733),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_563),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_526),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_563),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_618),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_642),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_563),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_526),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_883)
);

BUFx12f_ASAP7_75t_L g884 ( 
.A(n_775),
.Y(n_884)
);

OA21x2_ASAP7_75t_L g885 ( 
.A1(n_798),
.A2(n_553),
.B(n_542),
.Y(n_885)
);

NOR2x1_ASAP7_75t_L g886 ( 
.A(n_642),
.B(n_384),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_563),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_565),
.A2(n_386),
.B(n_385),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_739),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_748),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_567),
.A2(n_388),
.B(n_387),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_803),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_803),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_513),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_794),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_794),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_748),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_748),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_756),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_498),
.B(n_19),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_498),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_505),
.B(n_20),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_509),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_568),
.A2(n_391),
.B(n_390),
.Y(n_904)
);

BUFx12f_ASAP7_75t_L g905 ( 
.A(n_707),
.Y(n_905)
);

OA21x2_ASAP7_75t_L g906 ( 
.A1(n_586),
.A2(n_398),
.B(n_395),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_509),
.Y(n_907)
);

BUFx8_ASAP7_75t_L g908 ( 
.A(n_783),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_518),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_660),
.B(n_21),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_581),
.A2(n_25),
.B1(n_22),
.B2(n_23),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_513),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_518),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_660),
.B(n_22),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_527),
.B(n_399),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_614),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_578),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_799),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_639),
.B(n_26),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_799),
.Y(n_920)
);

CKINVDCx6p67_ASAP7_75t_R g921 ( 
.A(n_848),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_841),
.Y(n_922)
);

AND3x2_ASAP7_75t_L g923 ( 
.A(n_919),
.B(n_757),
.C(n_667),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_840),
.B(n_512),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_905),
.B(n_627),
.Y(n_925)
);

NAND2xp33_ASAP7_75t_L g926 ( 
.A(n_831),
.B(n_748),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_820),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_831),
.B(n_892),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_820),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_831),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_L g931 ( 
.A(n_831),
.B(n_635),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_860),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_822),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_L g934 ( 
.A(n_856),
.B(n_731),
.C(n_666),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_841),
.B(n_714),
.Y(n_935)
);

INVx8_ASAP7_75t_L g936 ( 
.A(n_824),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_860),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_860),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_822),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_823),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_834),
.B(n_591),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_861),
.B(n_899),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_823),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_825),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_870),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_848),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_821),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_825),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_826),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_900),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_870),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_834),
.B(n_610),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_826),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_840),
.B(n_512),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_830),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_830),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_870),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_856),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_900),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_840),
.B(n_808),
.Y(n_960)
);

INVx5_ASAP7_75t_L g961 ( 
.A(n_831),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_880),
.B(n_530),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_832),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_872),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_864),
.B(n_615),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_832),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_880),
.B(n_707),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_836),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_902),
.B(n_761),
.C(n_816),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_833),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_900),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_833),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_857),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_827),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_838),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_L g976 ( 
.A(n_892),
.B(n_635),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_902),
.B(n_816),
.C(n_520),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_838),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_851),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_845),
.B(n_636),
.Y(n_980)
);

NAND3xp33_ASAP7_75t_L g981 ( 
.A(n_910),
.B(n_520),
.C(n_517),
.Y(n_981)
);

BUFx6f_ASAP7_75t_SL g982 ( 
.A(n_818),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_829),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_894),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_853),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_845),
.B(n_640),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_884),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_868),
.B(n_920),
.Y(n_988)
);

INVxp67_ASAP7_75t_SL g989 ( 
.A(n_910),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_866),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_914),
.A2(n_491),
.B1(n_494),
.B2(n_488),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_864),
.B(n_648),
.Y(n_992)
);

AO21x2_ASAP7_75t_L g993 ( 
.A1(n_819),
.A2(n_651),
.B(n_649),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_881),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_881),
.B(n_530),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_855),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_859),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_818),
.A2(n_914),
.B1(n_836),
.B2(n_849),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_L g999 ( 
.A(n_835),
.B(n_535),
.C(n_529),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_876),
.B(n_920),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_859),
.Y(n_1001)
);

INVx5_ASAP7_75t_L g1002 ( 
.A(n_881),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_895),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_894),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_871),
.B(n_663),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_882),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_896),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_887),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_905),
.B(n_711),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_824),
.B(n_711),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_887),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_885),
.Y(n_1012)
);

AND2x2_ASAP7_75t_SL g1013 ( 
.A(n_842),
.B(n_533),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_893),
.B(n_837),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_877),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_837),
.B(n_671),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_877),
.Y(n_1017)
);

AOI21x1_ASAP7_75t_L g1018 ( 
.A1(n_819),
.A2(n_673),
.B(n_672),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_879),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_879),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_907),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_909),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_889),
.B(n_674),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_821),
.Y(n_1024)
);

OAI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_839),
.A2(n_858),
.B1(n_884),
.B2(n_911),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_821),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_844),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_885),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_889),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_893),
.B(n_637),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_828),
.A2(n_692),
.B(n_679),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_918),
.B(n_704),
.Y(n_1032)
);

AO21x2_ASAP7_75t_L g1033 ( 
.A1(n_828),
.A2(n_735),
.B(n_732),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_885),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_918),
.Y(n_1035)
);

BUFx10_ASAP7_75t_L g1036 ( 
.A(n_849),
.Y(n_1036)
);

INVx6_ASAP7_75t_L g1037 ( 
.A(n_852),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_913),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_913),
.B(n_638),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_874),
.B(n_738),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_886),
.B(n_745),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_L g1042 ( 
.A(n_854),
.B(n_771),
.C(n_644),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_913),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_885),
.A2(n_496),
.B1(n_497),
.B2(n_495),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_901),
.B(n_644),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_903),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_903),
.B(n_771),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_873),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_852),
.B(n_763),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_908),
.B(n_773),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_908),
.B(n_765),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_SL g1052 ( 
.A(n_908),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_852),
.B(n_766),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_846),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_919),
.B(n_711),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_852),
.B(n_773),
.Y(n_1056)
);

INVxp33_ASAP7_75t_L g1057 ( 
.A(n_847),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_863),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_852),
.B(n_779),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_863),
.Y(n_1060)
);

NAND2xp33_ASAP7_75t_L g1061 ( 
.A(n_862),
.B(n_774),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_867),
.Y(n_1062)
);

BUFx10_ASAP7_75t_L g1063 ( 
.A(n_912),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_867),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_865),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_917),
.B(n_772),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_842),
.Y(n_1067)
);

INVxp33_ASAP7_75t_L g1068 ( 
.A(n_916),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_842),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_842),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_869),
.B(n_806),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_912),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_843),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_843),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_843),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1048),
.B(n_774),
.Y(n_1076)
);

NAND2x1_ASAP7_75t_L g1077 ( 
.A(n_964),
.B(n_843),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_982),
.A2(n_883),
.B1(n_878),
.B2(n_601),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_942),
.B(n_917),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_958),
.B(n_776),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_925),
.B(n_578),
.Y(n_1081)
);

NAND2xp33_ASAP7_75t_L g1082 ( 
.A(n_961),
.B(n_936),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_925),
.B(n_601),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_922),
.B(n_779),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_936),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_989),
.B(n_786),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1072),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_960),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_984),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_935),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_982),
.A2(n_1055),
.B1(n_998),
.B2(n_967),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_932),
.B(n_787),
.Y(n_1092)
);

INVx8_ASAP7_75t_L g1093 ( 
.A(n_936),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_924),
.B(n_954),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_L g1095 ( 
.A(n_977),
.B(n_791),
.C(n_780),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_968),
.B(n_780),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_936),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1054),
.B(n_538),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_937),
.B(n_938),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_1063),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_1009),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1030),
.B(n_539),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_930),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_1063),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_SL g1105 ( 
.A(n_1052),
.B(n_634),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1010),
.B(n_791),
.Y(n_1106)
);

INVxp67_ASAP7_75t_L g1107 ( 
.A(n_1063),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_930),
.B(n_501),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_925),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_990),
.Y(n_1110)
);

BUFx5_ASAP7_75t_L g1111 ( 
.A(n_1058),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1016),
.B(n_683),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_994),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_995),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_934),
.B(n_510),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_995),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_1052),
.Y(n_1117)
);

INVxp67_ASAP7_75t_SL g1118 ( 
.A(n_1012),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1038),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_995),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_SL g1121 ( 
.A(n_925),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1043),
.Y(n_1122)
);

NAND2xp33_ASAP7_75t_L g1123 ( 
.A(n_1044),
.B(n_545),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1014),
.B(n_552),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_921),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_921),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_SL g1127 ( 
.A1(n_984),
.A2(n_551),
.B1(n_554),
.B2(n_521),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_945),
.B(n_573),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_950),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_931),
.A2(n_915),
.B(n_850),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_969),
.B(n_575),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_951),
.B(n_850),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_957),
.B(n_850),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_962),
.B(n_492),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1043),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1057),
.B(n_965),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_992),
.B(n_584),
.Y(n_1137)
);

HB1xp67_ASAP7_75t_L g1138 ( 
.A(n_1052),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1051),
.B(n_588),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_999),
.B(n_590),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_962),
.B(n_595),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1043),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_982),
.A2(n_688),
.B1(n_697),
.B2(n_634),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1039),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_950),
.A2(n_500),
.B1(n_507),
.B2(n_499),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_946),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1057),
.B(n_981),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1042),
.B(n_597),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1068),
.A2(n_697),
.B1(n_767),
.B2(n_688),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_959),
.B(n_971),
.Y(n_1150)
);

AOI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_931),
.A2(n_514),
.B1(n_516),
.B2(n_508),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1050),
.B(n_603),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1036),
.B(n_962),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1045),
.Y(n_1154)
);

NOR3xp33_ASAP7_75t_L g1155 ( 
.A(n_1025),
.B(n_612),
.C(n_528),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_987),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1036),
.B(n_616),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1002),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1068),
.A2(n_525),
.B1(n_531),
.B2(n_523),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1012),
.B(n_1028),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1036),
.B(n_620),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1046),
.Y(n_1162)
);

AND2x6_ASAP7_75t_L g1163 ( 
.A(n_1067),
.B(n_533),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1021),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1022),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1047),
.B(n_630),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_991),
.A2(n_784),
.B1(n_789),
.B2(n_767),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_974),
.B(n_659),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1002),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_983),
.B(n_665),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1066),
.B(n_976),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_1040),
.B(n_489),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1056),
.B(n_668),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1002),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1034),
.A2(n_546),
.B1(n_559),
.B2(n_550),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_976),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_973),
.B(n_675),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1003),
.B(n_678),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1015),
.B(n_906),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_1059),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1019),
.B(n_906),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1007),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_973),
.B(n_681),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1000),
.B(n_724),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_987),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1029),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1017),
.B(n_725),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1035),
.Y(n_1188)
);

INVx4_ASAP7_75t_L g1189 ( 
.A(n_1037),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_923),
.B(n_493),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_928),
.A2(n_560),
.B1(n_572),
.B2(n_561),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1004),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_941),
.B(n_768),
.Y(n_1193)
);

INVx5_ASAP7_75t_L g1194 ( 
.A(n_1037),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1017),
.B(n_800),
.Y(n_1195)
);

INVx6_ASAP7_75t_L g1196 ( 
.A(n_1037),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1041),
.B(n_502),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1041),
.B(n_503),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_988),
.B(n_504),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_952),
.B(n_537),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1004),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1023),
.B(n_540),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1067),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_980),
.B(n_698),
.Y(n_1204)
);

OAI221xp5_ASAP7_75t_L g1205 ( 
.A1(n_1032),
.A2(n_676),
.B1(n_770),
.B2(n_661),
.C(n_657),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1020),
.B(n_888),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_927),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1020),
.B(n_888),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_928),
.A2(n_1062),
.B1(n_1064),
.B2(n_1060),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_926),
.B(n_562),
.C(n_556),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1018),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1032),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_L g1213 ( 
.A(n_1070),
.B(n_784),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_986),
.A2(n_809),
.B1(n_789),
.B2(n_566),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_986),
.B(n_698),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1013),
.B(n_891),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1005),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_929),
.B(n_891),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_933),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1005),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1031),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1073),
.B(n_564),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_939),
.B(n_698),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_940),
.B(n_904),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1061),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_940),
.B(n_534),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_943),
.B(n_534),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_943),
.B(n_543),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_944),
.B(n_543),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_993),
.B(n_569),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_948),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_949),
.B(n_698),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_993),
.B(n_809),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_953),
.B(n_544),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_993),
.A2(n_580),
.B1(n_583),
.B2(n_577),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1074),
.A2(n_551),
.B1(n_554),
.B2(n_521),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_955),
.B(n_571),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_956),
.B(n_576),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_956),
.B(n_582),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1033),
.A2(n_593),
.B1(n_599),
.B2(n_589),
.Y(n_1240)
);

OR2x2_ASAP7_75t_SL g1241 ( 
.A(n_926),
.B(n_587),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_963),
.B(n_544),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_963),
.B(n_555),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_966),
.B(n_555),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1033),
.B(n_807),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1071),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1049),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1073),
.B(n_585),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1069),
.A2(n_813),
.B1(n_592),
.B2(n_596),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1049),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_970),
.B(n_557),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_972),
.B(n_712),
.Y(n_1252)
);

INVxp33_ASAP7_75t_L g1253 ( 
.A(n_1053),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1075),
.A2(n_594),
.B1(n_600),
.B2(n_598),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1075),
.A2(n_626),
.B1(n_646),
.B2(n_587),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_975),
.B(n_604),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_978),
.Y(n_1257)
);

NAND2x1_ASAP7_75t_L g1258 ( 
.A(n_979),
.B(n_557),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_979),
.B(n_607),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_985),
.B(n_712),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_947),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_996),
.Y(n_1262)
);

BUFx5_ASAP7_75t_L g1263 ( 
.A(n_996),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_997),
.A2(n_617),
.B1(n_619),
.B2(n_611),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_997),
.A2(n_625),
.B1(n_645),
.B2(n_623),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1001),
.B(n_658),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1006),
.B(n_669),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1008),
.A2(n_536),
.B(n_490),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1011),
.B(n_792),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1024),
.B(n_574),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1024),
.A2(n_710),
.B(n_570),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1026),
.B(n_685),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1026),
.B(n_574),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_947),
.B(n_792),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1027),
.B(n_689),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1093),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1132),
.A2(n_1133),
.B(n_1118),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1085),
.B(n_693),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1097),
.B(n_730),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1088),
.B(n_626),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1117),
.B(n_778),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1080),
.B(n_694),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1093),
.B(n_699),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1080),
.B(n_702),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1090),
.A2(n_602),
.B(n_606),
.C(n_605),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1096),
.B(n_646),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1099),
.A2(n_677),
.B1(n_690),
.B2(n_662),
.Y(n_1287)
);

AOI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1213),
.A2(n_709),
.B1(n_715),
.B2(n_706),
.Y(n_1288)
);

CKINVDCx6p67_ASAP7_75t_R g1289 ( 
.A(n_1093),
.Y(n_1289)
);

AOI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1245),
.A2(n_609),
.B(n_608),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1086),
.B(n_718),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1086),
.B(n_1154),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1099),
.A2(n_677),
.B1(n_690),
.B2(n_662),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1155),
.A2(n_613),
.B(n_624),
.C(n_622),
.Y(n_1294)
);

INVx11_ASAP7_75t_L g1295 ( 
.A(n_1121),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1087),
.B(n_695),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1150),
.A2(n_716),
.B1(n_717),
.B2(n_695),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1262),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1126),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1101),
.B(n_716),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1079),
.B(n_717),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1144),
.B(n_721),
.Y(n_1302)
);

CKINVDCx14_ASAP7_75t_R g1303 ( 
.A(n_1125),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1205),
.A2(n_632),
.B(n_641),
.C(n_628),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1076),
.B(n_722),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1103),
.B(n_728),
.Y(n_1306)
);

OR2x6_ASAP7_75t_L g1307 ( 
.A(n_1167),
.B(n_579),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1089),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1084),
.B(n_720),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1189),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1105),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1256),
.B(n_729),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1233),
.A2(n_737),
.B1(n_753),
.B2(n_746),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1150),
.A2(n_1241),
.B1(n_1233),
.B2(n_1175),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1109),
.B(n_720),
.Y(n_1315)
);

NOR3xp33_ASAP7_75t_L g1316 ( 
.A(n_1167),
.B(n_1127),
.C(n_1255),
.Y(n_1316)
);

CKINVDCx10_ASAP7_75t_R g1317 ( 
.A(n_1121),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1094),
.A2(n_652),
.B(n_653),
.C(n_643),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1266),
.B(n_759),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1146),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1255),
.B(n_1149),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1129),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1209),
.A2(n_1181),
.B(n_1179),
.Y(n_1323)
);

CKINVDCx10_ASAP7_75t_R g1324 ( 
.A(n_1192),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1092),
.B(n_764),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1263),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1182),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1189),
.Y(n_1328)
);

AOI21xp33_ASAP7_75t_L g1329 ( 
.A1(n_1230),
.A2(n_1171),
.B(n_1222),
.Y(n_1329)
);

INVx3_ASAP7_75t_SL g1330 ( 
.A(n_1081),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1103),
.B(n_769),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1092),
.B(n_797),
.Y(n_1332)
);

BUFx12f_ASAP7_75t_L g1333 ( 
.A(n_1117),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1103),
.B(n_805),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1151),
.A2(n_777),
.B1(n_782),
.B2(n_760),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1128),
.A2(n_1078),
.B(n_1134),
.C(n_1153),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1106),
.B(n_760),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1248),
.A2(n_656),
.B(n_664),
.C(n_655),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1136),
.B(n_810),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1147),
.B(n_670),
.Y(n_1340)
);

NAND2xp33_ASAP7_75t_R g1341 ( 
.A(n_1081),
.B(n_27),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_SL g1342 ( 
.A(n_1083),
.B(n_777),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1206),
.A2(n_1208),
.B(n_1218),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1164),
.B(n_680),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1203),
.B(n_752),
.Y(n_1345)
);

O2A1O1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1128),
.A2(n_686),
.B(n_691),
.C(n_682),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1165),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1201),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1083),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1263),
.Y(n_1350)
);

AND2x2_ASAP7_75t_SL g1351 ( 
.A(n_1143),
.B(n_782),
.Y(n_1351)
);

CKINVDCx10_ASAP7_75t_R g1352 ( 
.A(n_1172),
.Y(n_1352)
);

AND2x2_ASAP7_75t_SL g1353 ( 
.A(n_1214),
.B(n_1082),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1263),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1156),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1145),
.B(n_1098),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1224),
.A2(n_793),
.B(n_703),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1091),
.B(n_801),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1180),
.B(n_696),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1100),
.B(n_801),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1102),
.B(n_705),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1235),
.A2(n_719),
.B(n_713),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1078),
.A2(n_727),
.B1(n_734),
.B2(n_723),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1162),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_L g1365 ( 
.A(n_1104),
.B(n_736),
.Y(n_1365)
);

AO22x1_ASAP7_75t_L g1366 ( 
.A1(n_1107),
.A2(n_741),
.B1(n_742),
.B2(n_740),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1211),
.A2(n_1065),
.B(n_744),
.Y(n_1367)
);

OAI321xp33_ASAP7_75t_L g1368 ( 
.A1(n_1271),
.A2(n_750),
.A3(n_747),
.B1(n_751),
.B2(n_749),
.C(n_743),
.Y(n_1368)
);

OAI21xp33_ASAP7_75t_L g1369 ( 
.A1(n_1159),
.A2(n_1254),
.B(n_1249),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1221),
.A2(n_1065),
.B(n_755),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1240),
.A2(n_1220),
.B(n_1217),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1176),
.A2(n_758),
.B1(n_762),
.B2(n_754),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1187),
.A2(n_1065),
.B(n_785),
.Y(n_1373)
);

AND2x4_ASAP7_75t_SL g1374 ( 
.A(n_1138),
.B(n_621),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1095),
.A2(n_788),
.B1(n_790),
.B2(n_781),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1114),
.A2(n_796),
.B(n_802),
.C(n_795),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1116),
.A2(n_811),
.B(n_812),
.C(n_804),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1112),
.A2(n_817),
.B1(n_815),
.B2(n_629),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1185),
.B(n_621),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1202),
.B(n_633),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1195),
.A2(n_650),
.B(n_647),
.Y(n_1381)
);

AO21x1_ASAP7_75t_L g1382 ( 
.A1(n_1268),
.A2(n_650),
.B(n_647),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_1196),
.Y(n_1383)
);

OAI321xp33_ASAP7_75t_L g1384 ( 
.A1(n_1191),
.A2(n_814),
.A3(n_897),
.B1(n_898),
.B2(n_890),
.C(n_875),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1139),
.B(n_28),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1120),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1115),
.B(n_30),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1199),
.A2(n_897),
.B(n_890),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1141),
.B(n_1124),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1172),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1190),
.B(n_32),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1196),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_R g1393 ( 
.A(n_1123),
.B(n_33),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1257),
.A2(n_407),
.B(n_404),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1200),
.B(n_34),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1110),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1113),
.A2(n_1170),
.B(n_1168),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1263),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1111),
.B(n_37),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1258),
.Y(n_1400)
);

OR2x6_ASAP7_75t_L g1401 ( 
.A(n_1236),
.B(n_38),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1197),
.B(n_39),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1186),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_1403)
);

NOR3xp33_ASAP7_75t_L g1404 ( 
.A(n_1140),
.B(n_41),
.C(n_43),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1212),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1131),
.B(n_43),
.C(n_44),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1264),
.A2(n_47),
.B1(n_44),
.B2(n_45),
.Y(n_1407)
);

NAND3xp33_ASAP7_75t_L g1408 ( 
.A(n_1152),
.B(n_45),
.C(n_47),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1166),
.B(n_48),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1246),
.A2(n_423),
.B(n_422),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1226),
.A2(n_1228),
.B1(n_1229),
.B2(n_1227),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1196),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1259),
.B(n_1267),
.Y(n_1413)
);

BUFx4f_ASAP7_75t_L g1414 ( 
.A(n_1163),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1111),
.Y(n_1415)
);

NAND3x1_ASAP7_75t_L g1416 ( 
.A(n_1265),
.B(n_49),
.C(n_50),
.Y(n_1416)
);

AO21x1_ASAP7_75t_L g1417 ( 
.A1(n_1270),
.A2(n_52),
.B(n_53),
.Y(n_1417)
);

O2A1O1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1226),
.A2(n_58),
.B(n_53),
.C(n_54),
.Y(n_1418)
);

BUFx12f_ASAP7_75t_L g1419 ( 
.A(n_1172),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1227),
.A2(n_1229),
.B(n_1234),
.C(n_1228),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1188),
.B(n_54),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1237),
.B(n_58),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1158),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1238),
.B(n_59),
.Y(n_1424)
);

INVx4_ASAP7_75t_L g1425 ( 
.A(n_1163),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1242),
.A2(n_1243),
.B1(n_1251),
.B2(n_1244),
.Y(n_1426)
);

OAI321xp33_ASAP7_75t_L g1427 ( 
.A1(n_1239),
.A2(n_59),
.A3(n_60),
.B1(n_61),
.B2(n_63),
.C(n_66),
.Y(n_1427)
);

NOR2x1_ASAP7_75t_L g1428 ( 
.A(n_1157),
.B(n_60),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1244),
.A2(n_68),
.B1(n_63),
.B2(n_67),
.Y(n_1429)
);

OAI22x1_ASAP7_75t_L g1430 ( 
.A1(n_1161),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1207),
.A2(n_439),
.B(n_436),
.Y(n_1431)
);

AO21x1_ASAP7_75t_L g1432 ( 
.A1(n_1270),
.A2(n_1273),
.B(n_1251),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1198),
.B(n_71),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_SL g1434 ( 
.A1(n_1225),
.A2(n_442),
.B(n_447),
.C(n_441),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1272),
.B(n_74),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1275),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1163),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1177),
.B(n_78),
.Y(n_1438)
);

BUFx8_ASAP7_75t_L g1439 ( 
.A(n_1163),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1163),
.A2(n_1148),
.B1(n_1178),
.B2(n_1137),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1210),
.B(n_78),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1194),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1219),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1194),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1253),
.B(n_81),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1119),
.A2(n_85),
.B(n_82),
.C(n_83),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1231),
.Y(n_1447)
);

INVx3_ASAP7_75t_SL g1448 ( 
.A(n_1204),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1194),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1122),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1169),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1174),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1183),
.A2(n_1193),
.B1(n_1250),
.B2(n_1247),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1135),
.B(n_86),
.Y(n_1454)
);

OAI22x1_ASAP7_75t_L g1455 ( 
.A1(n_1142),
.A2(n_96),
.B1(n_93),
.B2(n_94),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1273),
.A2(n_474),
.B(n_472),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1184),
.B(n_93),
.Y(n_1457)
);

O2A1O1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1215),
.A2(n_97),
.B(n_94),
.C(n_96),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1261),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1173),
.B(n_97),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1108),
.B(n_98),
.Y(n_1461)
);

O2A1O1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1223),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1232),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1252),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1260),
.B(n_102),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1269),
.A2(n_106),
.B(n_104),
.C(n_105),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1261),
.B(n_105),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1274),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1094),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1097),
.B(n_110),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1216),
.A2(n_112),
.B(n_113),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1080),
.B(n_112),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1088),
.B(n_114),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1080),
.B(n_114),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1262),
.Y(n_1475)
);

OAI21xp33_ASAP7_75t_L g1476 ( 
.A1(n_1090),
.A2(n_115),
.B(n_116),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1203),
.Y(n_1477)
);

AOI21xp33_ASAP7_75t_L g1478 ( 
.A1(n_1245),
.A2(n_115),
.B(n_116),
.Y(n_1478)
);

AND2x2_ASAP7_75t_SL g1479 ( 
.A(n_1081),
.B(n_117),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_SL g1480 ( 
.A(n_1085),
.B(n_118),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1099),
.A2(n_121),
.B1(n_118),
.B2(n_120),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1090),
.B(n_121),
.Y(n_1482)
);

A2O1A1Ixp33_ASAP7_75t_L g1483 ( 
.A1(n_1094),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1099),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1088),
.B(n_125),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_SL g1486 ( 
.A(n_1085),
.B(n_126),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1080),
.B(n_127),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1099),
.A2(n_132),
.B1(n_128),
.B2(n_130),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1080),
.B(n_130),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1093),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1160),
.A2(n_133),
.B(n_134),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1292),
.B(n_134),
.Y(n_1492)
);

NAND2x1_ASAP7_75t_L g1493 ( 
.A(n_1276),
.B(n_135),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1369),
.B(n_1336),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1276),
.B(n_136),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1287),
.A2(n_136),
.B(n_137),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1356),
.B(n_1327),
.Y(n_1497)
);

INVx1_ASAP7_75t_SL g1498 ( 
.A(n_1320),
.Y(n_1498)
);

AO31x2_ASAP7_75t_L g1499 ( 
.A1(n_1432),
.A2(n_140),
.A3(n_138),
.B(n_139),
.Y(n_1499)
);

AO31x2_ASAP7_75t_L g1500 ( 
.A1(n_1323),
.A2(n_142),
.A3(n_138),
.B(n_140),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1347),
.B(n_142),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1364),
.B(n_1290),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1289),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_SL g1504 ( 
.A1(n_1425),
.A2(n_146),
.B(n_147),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1290),
.B(n_1436),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_SL g1506 ( 
.A1(n_1425),
.A2(n_1314),
.B(n_1471),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1421),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_SL g1508 ( 
.A1(n_1314),
.A2(n_148),
.B(n_149),
.Y(n_1508)
);

OAI21xp33_ASAP7_75t_L g1509 ( 
.A1(n_1342),
.A2(n_150),
.B(n_151),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1343),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1329),
.A2(n_153),
.B(n_155),
.C(n_156),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1307),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1318),
.B(n_157),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_SL g1514 ( 
.A(n_1307),
.B(n_158),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1307),
.B(n_159),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1396),
.B(n_159),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1490),
.B(n_160),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1490),
.B(n_160),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1296),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1447),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1411),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1357),
.A2(n_166),
.B(n_167),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1333),
.B(n_352),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1313),
.B(n_169),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1386),
.Y(n_1525)
);

INVx6_ASAP7_75t_SL g1526 ( 
.A(n_1470),
.Y(n_1526)
);

NOR2x1_ASAP7_75t_SL g1527 ( 
.A(n_1457),
.B(n_1411),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1287),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1408),
.B(n_170),
.C(n_171),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1329),
.A2(n_170),
.B(n_171),
.C(n_173),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1344),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1426),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_1532)
);

NOR2x1_ASAP7_75t_L g1533 ( 
.A(n_1299),
.B(n_175),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1470),
.Y(n_1534)
);

NAND2x1_ASAP7_75t_L g1535 ( 
.A(n_1449),
.B(n_178),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1355),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1348),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1479),
.B(n_1316),
.Y(n_1538)
);

A2O1A1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1471),
.A2(n_183),
.B(n_185),
.C(n_186),
.Y(n_1539)
);

INVx4_ASAP7_75t_L g1540 ( 
.A(n_1295),
.Y(n_1540)
);

AO31x2_ASAP7_75t_L g1541 ( 
.A1(n_1417),
.A2(n_188),
.A3(n_189),
.B(n_191),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1361),
.B(n_192),
.Y(n_1542)
);

BUFx4f_ASAP7_75t_SL g1543 ( 
.A(n_1308),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1426),
.A2(n_193),
.B(n_196),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1414),
.B(n_197),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1413),
.A2(n_197),
.B(n_200),
.Y(n_1546)
);

AO21x2_ASAP7_75t_L g1547 ( 
.A1(n_1357),
.A2(n_201),
.B(n_202),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1380),
.B(n_203),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1280),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1293),
.B(n_205),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1367),
.A2(n_206),
.B(n_207),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1301),
.B(n_207),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1370),
.A2(n_208),
.B(n_209),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1340),
.B(n_1338),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1482),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1372),
.B(n_209),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1309),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1322),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1286),
.B(n_210),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1359),
.B(n_212),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1394),
.A2(n_213),
.B(n_215),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1401),
.B(n_351),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1449),
.Y(n_1563)
);

AO31x2_ASAP7_75t_L g1564 ( 
.A1(n_1469),
.A2(n_216),
.A3(n_217),
.B(n_218),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1435),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1324),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1442),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1293),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1389),
.B(n_219),
.Y(n_1569)
);

A2O1A1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1478),
.A2(n_219),
.B(n_220),
.C(n_222),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1330),
.Y(n_1571)
);

NOR2x1_ASAP7_75t_L g1572 ( 
.A(n_1401),
.B(n_225),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1401),
.B(n_226),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1472),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1474),
.Y(n_1575)
);

NAND2xp33_ASAP7_75t_SL g1576 ( 
.A(n_1393),
.B(n_227),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1487),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1442),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1297),
.A2(n_1337),
.B1(n_1335),
.B2(n_1360),
.Y(n_1579)
);

NAND2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1414),
.B(n_230),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1297),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1374),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1373),
.A2(n_232),
.B(n_233),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1321),
.B(n_234),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1346),
.B(n_234),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_SL g1586 ( 
.A(n_1457),
.B(n_235),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1387),
.B(n_236),
.C(n_237),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1282),
.B(n_238),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1335),
.B(n_238),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1317),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1284),
.B(n_239),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1303),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1440),
.B(n_241),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1349),
.B(n_242),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1291),
.B(n_244),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1489),
.Y(n_1596)
);

AOI221xp5_ASAP7_75t_L g1597 ( 
.A1(n_1285),
.A2(n_249),
.B1(n_253),
.B2(n_254),
.C(n_255),
.Y(n_1597)
);

OA22x2_ASAP7_75t_L g1598 ( 
.A1(n_1363),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1376),
.B(n_259),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1439),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1377),
.B(n_260),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_SL g1602 ( 
.A(n_1341),
.B(n_263),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1378),
.B(n_265),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1325),
.B(n_265),
.Y(n_1604)
);

CKINVDCx16_ASAP7_75t_R g1605 ( 
.A(n_1390),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1332),
.B(n_1473),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1388),
.A2(n_266),
.B(n_267),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1485),
.B(n_266),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1353),
.B(n_267),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1339),
.B(n_268),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1352),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1304),
.B(n_272),
.Y(n_1612)
);

NAND2x1p5_ASAP7_75t_L g1613 ( 
.A(n_1298),
.B(n_273),
.Y(n_1613)
);

INVx4_ASAP7_75t_L g1614 ( 
.A(n_1298),
.Y(n_1614)
);

AOI211x1_ASAP7_75t_L g1615 ( 
.A1(n_1478),
.A2(n_275),
.B(n_278),
.C(n_279),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1459),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_1439),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1415),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1326),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1366),
.B(n_281),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1454),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1443),
.B(n_285),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1371),
.A2(n_286),
.B(n_287),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1450),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1300),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1351),
.B(n_1311),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1455),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1419),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1305),
.B(n_289),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1430),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1358),
.B(n_290),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1456),
.A2(n_293),
.B(n_294),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1288),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1409),
.A2(n_295),
.B(n_296),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1418),
.A2(n_297),
.B(n_298),
.C(n_299),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1362),
.B(n_1312),
.Y(n_1636)
);

O2A1O1Ixp5_ASAP7_75t_L g1637 ( 
.A1(n_1467),
.A2(n_297),
.B(n_299),
.C(n_300),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1319),
.B(n_302),
.Y(n_1638)
);

A2O1A1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1483),
.A2(n_304),
.B(n_306),
.C(n_307),
.Y(n_1639)
);

AO31x2_ASAP7_75t_L g1640 ( 
.A1(n_1481),
.A2(n_306),
.A3(n_308),
.B(n_309),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1457),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1381),
.A2(n_308),
.B(n_310),
.Y(n_1642)
);

AO22x2_ASAP7_75t_L g1643 ( 
.A1(n_1481),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_1643)
);

NOR2xp67_ASAP7_75t_L g1644 ( 
.A(n_1315),
.B(n_311),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1437),
.A2(n_314),
.B1(n_318),
.B2(n_320),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1402),
.B(n_322),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1422),
.A2(n_323),
.B(n_324),
.Y(n_1647)
);

AO31x2_ASAP7_75t_L g1648 ( 
.A1(n_1484),
.A2(n_323),
.A3(n_325),
.B(n_326),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1433),
.B(n_326),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1350),
.Y(n_1650)
);

NOR2xp67_ASAP7_75t_L g1651 ( 
.A(n_1368),
.B(n_327),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1424),
.A2(n_328),
.B(n_329),
.Y(n_1652)
);

AND3x2_ASAP7_75t_L g1653 ( 
.A(n_1404),
.B(n_329),
.C(n_330),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1484),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1488),
.A2(n_335),
.B(n_336),
.C(n_337),
.Y(n_1655)
);

AOI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1365),
.A2(n_341),
.B(n_342),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1294),
.B(n_342),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1379),
.A2(n_1391),
.B1(n_1445),
.B2(n_1385),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1375),
.B(n_343),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1405),
.B(n_343),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1354),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1488),
.A2(n_1453),
.B1(n_1429),
.B2(n_1475),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1302),
.B(n_1395),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1398),
.Y(n_1664)
);

AOI221x1_ASAP7_75t_L g1665 ( 
.A1(n_1476),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.C(n_350),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_SL g1666 ( 
.A(n_1283),
.B(n_1429),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1461),
.B(n_1438),
.Y(n_1667)
);

AND3x2_ASAP7_75t_L g1668 ( 
.A(n_1281),
.B(n_1279),
.C(n_1416),
.Y(n_1668)
);

BUFx12f_ASAP7_75t_L g1669 ( 
.A(n_1281),
.Y(n_1669)
);

AO31x2_ASAP7_75t_L g1670 ( 
.A1(n_1446),
.A2(n_1403),
.A3(n_1491),
.B(n_1410),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1407),
.B(n_1278),
.Y(n_1671)
);

INVx2_ASAP7_75t_SL g1672 ( 
.A(n_1279),
.Y(n_1672)
);

NOR2xp67_ASAP7_75t_L g1673 ( 
.A(n_1406),
.B(n_1460),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1480),
.B(n_1486),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1465),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1428),
.B(n_1306),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1468),
.A2(n_1464),
.B(n_1458),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1331),
.B(n_1334),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1462),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1444),
.B(n_1383),
.Y(n_1680)
);

NAND2xp33_ASAP7_75t_L g1681 ( 
.A(n_1448),
.B(n_1310),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1383),
.B(n_1392),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1441),
.A2(n_1452),
.B1(n_1451),
.B2(n_1423),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1466),
.Y(n_1684)
);

AND3x4_ASAP7_75t_L g1685 ( 
.A(n_1400),
.B(n_1427),
.C(n_1468),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1392),
.B(n_1412),
.Y(n_1686)
);

AO31x2_ASAP7_75t_L g1687 ( 
.A1(n_1434),
.A2(n_1384),
.A3(n_1444),
.B(n_1310),
.Y(n_1687)
);

O2A1O1Ixp5_ASAP7_75t_SL g1688 ( 
.A1(n_1412),
.A2(n_1271),
.B(n_1345),
.C(n_1357),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1328),
.Y(n_1689)
);

INVx6_ASAP7_75t_L g1690 ( 
.A(n_1328),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1463),
.B(n_1307),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1292),
.B(n_958),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1327),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1299),
.B(n_1126),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1292),
.B(n_958),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1276),
.B(n_1490),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1304),
.A2(n_1338),
.B1(n_1294),
.B2(n_1369),
.C(n_1285),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1292),
.B(n_958),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1292),
.B(n_958),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1307),
.B(n_1479),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1292),
.B(n_958),
.Y(n_1705)
);

NOR2x1_ASAP7_75t_L g1706 ( 
.A(n_1299),
.B(n_1126),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1289),
.Y(n_1707)
);

NAND2xp33_ASAP7_75t_SL g1708 ( 
.A(n_1425),
.B(n_1393),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1292),
.B(n_958),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1431),
.Y(n_1710)
);

AO31x2_ASAP7_75t_L g1711 ( 
.A1(n_1432),
.A2(n_1323),
.A3(n_1382),
.B(n_1417),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_SL g1712 ( 
.A(n_1316),
.B(n_1393),
.C(n_912),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1292),
.B(n_958),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1289),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1276),
.B(n_1490),
.Y(n_1715)
);

INVx3_ASAP7_75t_SL g1716 ( 
.A(n_1289),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1292),
.B(n_958),
.Y(n_1717)
);

NAND2x1p5_ASAP7_75t_L g1718 ( 
.A(n_1276),
.B(n_1490),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1292),
.B(n_958),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1327),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1277),
.A2(n_1323),
.B(n_1216),
.Y(n_1722)
);

NAND2x1p5_ASAP7_75t_L g1723 ( 
.A(n_1276),
.B(n_1490),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1307),
.B(n_1479),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1307),
.B(n_1479),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1292),
.B(n_958),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1292),
.B(n_958),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1327),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1292),
.B(n_958),
.Y(n_1731)
);

OAI21x1_ASAP7_75t_SL g1732 ( 
.A1(n_1425),
.A2(n_1314),
.B(n_1471),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1292),
.B(n_958),
.Y(n_1733)
);

INVx5_ASAP7_75t_L g1734 ( 
.A(n_1276),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1292),
.B(n_958),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1292),
.B(n_958),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1277),
.A2(n_1323),
.B(n_1216),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1292),
.B(n_958),
.Y(n_1738)
);

AOI211x1_ASAP7_75t_L g1739 ( 
.A1(n_1369),
.A2(n_1290),
.B(n_1314),
.C(n_1471),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1289),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1327),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1292),
.B(n_958),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1289),
.Y(n_1743)
);

A2O1A1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1329),
.A2(n_1420),
.B(n_1397),
.C(n_1290),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1327),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1320),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1292),
.B(n_958),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1327),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1749)
);

OA21x2_ASAP7_75t_L g1750 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1431),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_SL g1751 ( 
.A(n_1289),
.B(n_1093),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1292),
.B(n_958),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1277),
.A2(n_1323),
.B(n_1216),
.Y(n_1754)
);

AO31x2_ASAP7_75t_L g1755 ( 
.A1(n_1432),
.A2(n_1323),
.A3(n_1382),
.B(n_1417),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1327),
.Y(n_1756)
);

BUFx3_ASAP7_75t_L g1757 ( 
.A(n_1289),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1327),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1327),
.Y(n_1759)
);

BUFx6f_ASAP7_75t_L g1760 ( 
.A(n_1477),
.Y(n_1760)
);

NOR4xp25_ASAP7_75t_L g1761 ( 
.A(n_1416),
.B(n_1314),
.C(n_1427),
.D(n_1481),
.Y(n_1761)
);

O2A1O1Ixp5_ASAP7_75t_L g1762 ( 
.A1(n_1382),
.A2(n_1329),
.B(n_1357),
.C(n_1399),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1320),
.Y(n_1763)
);

AO31x2_ASAP7_75t_L g1764 ( 
.A1(n_1432),
.A2(n_1323),
.A3(n_1382),
.B(n_1417),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1289),
.Y(n_1765)
);

NOR2xp67_ASAP7_75t_L g1766 ( 
.A(n_1333),
.B(n_1125),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1292),
.B(n_958),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1276),
.B(n_1490),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1292),
.B(n_958),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1292),
.B(n_958),
.Y(n_1770)
);

OAI21x1_ASAP7_75t_SL g1771 ( 
.A1(n_1425),
.A2(n_1314),
.B(n_1471),
.Y(n_1771)
);

AO31x2_ASAP7_75t_L g1772 ( 
.A1(n_1432),
.A2(n_1323),
.A3(n_1382),
.B(n_1417),
.Y(n_1772)
);

OA22x2_ASAP7_75t_L g1773 ( 
.A1(n_1307),
.A2(n_1401),
.B1(n_1167),
.B2(n_1149),
.Y(n_1773)
);

OA21x2_ASAP7_75t_L g1774 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1431),
.Y(n_1774)
);

BUFx3_ASAP7_75t_L g1775 ( 
.A(n_1289),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1313),
.B(n_1091),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1323),
.A2(n_1130),
.B(n_1077),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1327),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1562),
.A2(n_1523),
.B1(n_1566),
.B2(n_1579),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1693),
.Y(n_1780)
);

INVx1_ASAP7_75t_SL g1781 ( 
.A(n_1716),
.Y(n_1781)
);

CKINVDCx20_ASAP7_75t_R g1782 ( 
.A(n_1716),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1757),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1773),
.A2(n_1538),
.B1(n_1626),
.B2(n_1562),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1721),
.Y(n_1785)
);

NAND2x1p5_ASAP7_75t_L g1786 ( 
.A(n_1757),
.B(n_1775),
.Y(n_1786)
);

NAND2x1p5_ASAP7_75t_L g1787 ( 
.A(n_1775),
.B(n_1734),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1568),
.B(n_1528),
.Y(n_1788)
);

OA21x2_ASAP7_75t_L g1789 ( 
.A1(n_1704),
.A2(n_1727),
.B(n_1719),
.Y(n_1789)
);

AOI21xp33_ASAP7_75t_L g1790 ( 
.A1(n_1494),
.A2(n_1569),
.B(n_1658),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1730),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1741),
.Y(n_1792)
);

A2O1A1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1655),
.A2(n_1744),
.B(n_1544),
.C(n_1539),
.Y(n_1793)
);

AO21x2_ASAP7_75t_L g1794 ( 
.A1(n_1719),
.A2(n_1728),
.B(n_1727),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1517),
.Y(n_1795)
);

OA21x2_ASAP7_75t_L g1796 ( 
.A1(n_1749),
.A2(n_1777),
.B(n_1753),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1773),
.A2(n_1562),
.B1(n_1581),
.B2(n_1528),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1702),
.B(n_1537),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1745),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1748),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1503),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1718),
.Y(n_1802)
);

OR2x4_ASAP7_75t_L g1803 ( 
.A(n_1712),
.B(n_1589),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_SL g1804 ( 
.A1(n_1701),
.A2(n_1724),
.B1(n_1725),
.B2(n_1586),
.Y(n_1804)
);

AO21x2_ASAP7_75t_L g1805 ( 
.A1(n_1753),
.A2(n_1777),
.B(n_1732),
.Y(n_1805)
);

BUFx2_ASAP7_75t_L g1806 ( 
.A(n_1526),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1756),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1744),
.A2(n_1762),
.B(n_1569),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1758),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1762),
.A2(n_1688),
.B(n_1636),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1536),
.Y(n_1811)
);

NAND2x1p5_ASAP7_75t_L g1812 ( 
.A(n_1734),
.B(n_1517),
.Y(n_1812)
);

AO22x2_ASAP7_75t_L g1813 ( 
.A1(n_1739),
.A2(n_1771),
.B1(n_1506),
.B2(n_1685),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1759),
.Y(n_1814)
);

INVxp67_ASAP7_75t_SL g1815 ( 
.A(n_1512),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1718),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1707),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1778),
.Y(n_1818)
);

AO21x2_ASAP7_75t_L g1819 ( 
.A1(n_1722),
.A2(n_1754),
.B(n_1737),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1531),
.B(n_1692),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1712),
.A2(n_1602),
.B1(n_1776),
.B2(n_1576),
.Y(n_1821)
);

INVx8_ASAP7_75t_L g1822 ( 
.A(n_1523),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1624),
.Y(n_1823)
);

AND2x6_ASAP7_75t_SL g1824 ( 
.A(n_1523),
.B(n_1590),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1695),
.B(n_1699),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1552),
.B(n_1559),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1525),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1520),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1707),
.Y(n_1829)
);

OAI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1710),
.A2(n_1774),
.B(n_1750),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1592),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1558),
.B(n_1527),
.Y(n_1832)
);

OAI21x1_ASAP7_75t_L g1833 ( 
.A1(n_1710),
.A2(n_1774),
.B(n_1750),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1550),
.B(n_1700),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1606),
.A2(n_1663),
.B(n_1662),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1705),
.B(n_1709),
.Y(n_1836)
);

AOI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1625),
.A2(n_1776),
.B1(n_1697),
.B2(n_1761),
.C(n_1505),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1713),
.B(n_1717),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1625),
.B(n_1631),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1502),
.A2(n_1554),
.B(n_1677),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1714),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_SL g1842 ( 
.A1(n_1666),
.A2(n_1514),
.B(n_1508),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1760),
.Y(n_1843)
);

AOI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1524),
.A2(n_1565),
.B1(n_1555),
.B2(n_1507),
.C(n_1496),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1534),
.A2(n_1526),
.B1(n_1512),
.B2(n_1584),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1643),
.A2(n_1641),
.B1(n_1515),
.B2(n_1598),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1534),
.B(n_1720),
.Y(n_1847)
);

NAND3x1_ASAP7_75t_L g1848 ( 
.A(n_1572),
.B(n_1573),
.C(n_1627),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1760),
.Y(n_1849)
);

BUFx2_ASAP7_75t_SL g1850 ( 
.A(n_1766),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1760),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1685),
.A2(n_1622),
.B1(n_1497),
.B2(n_1580),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1501),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1726),
.B(n_1729),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1516),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1731),
.B(n_1733),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1735),
.B(n_1736),
.Y(n_1857)
);

BUFx2_ASAP7_75t_L g1858 ( 
.A(n_1571),
.Y(n_1858)
);

CKINVDCx16_ASAP7_75t_R g1859 ( 
.A(n_1751),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1602),
.A2(n_1576),
.B1(n_1598),
.B2(n_1524),
.Y(n_1860)
);

NOR2xp33_ASAP7_75t_L g1861 ( 
.A(n_1738),
.B(n_1742),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1747),
.B(n_1752),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1767),
.B(n_1769),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1613),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1622),
.A2(n_1580),
.B1(n_1492),
.B2(n_1518),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1770),
.B(n_1675),
.Y(n_1866)
);

BUFx3_ASAP7_75t_L g1867 ( 
.A(n_1714),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1582),
.B(n_1740),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1615),
.B(n_1635),
.C(n_1539),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1740),
.B(n_1743),
.Y(n_1870)
);

AO22x2_ASAP7_75t_L g1871 ( 
.A1(n_1630),
.A2(n_1665),
.B1(n_1654),
.B2(n_1504),
.Y(n_1871)
);

OAI222xp33_ASAP7_75t_L g1872 ( 
.A1(n_1557),
.A2(n_1495),
.B1(n_1655),
.B2(n_1519),
.C1(n_1549),
.C2(n_1532),
.Y(n_1872)
);

INVx8_ASAP7_75t_L g1873 ( 
.A(n_1734),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1543),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1743),
.B(n_1765),
.Y(n_1875)
);

OR2x6_ASAP7_75t_L g1876 ( 
.A(n_1540),
.B(n_1600),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1495),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1533),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1594),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1513),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1521),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1617),
.B(n_1765),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1640),
.Y(n_1883)
);

BUFx2_ASAP7_75t_L g1884 ( 
.A(n_1543),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1574),
.B(n_1575),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1618),
.Y(n_1886)
);

NAND2x1_ASAP7_75t_L g1887 ( 
.A(n_1567),
.B(n_1578),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1577),
.B(n_1596),
.Y(n_1888)
);

BUFx4f_ASAP7_75t_SL g1889 ( 
.A(n_1498),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1691),
.B(n_1594),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1650),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1696),
.B(n_1715),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1611),
.B(n_1605),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1723),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1651),
.Y(n_1895)
);

INVx2_ASAP7_75t_SL g1896 ( 
.A(n_1540),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1621),
.B(n_1671),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1667),
.B(n_1560),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1669),
.Y(n_1899)
);

CKINVDCx20_ASAP7_75t_R g1900 ( 
.A(n_1746),
.Y(n_1900)
);

A2O1A1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1639),
.A2(n_1511),
.B(n_1530),
.C(n_1623),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1664),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_1694),
.Y(n_1903)
);

INVx4_ASAP7_75t_SL g1904 ( 
.A(n_1640),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1648),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1706),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1609),
.A2(n_1708),
.B1(n_1556),
.B2(n_1644),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1672),
.B(n_1603),
.Y(n_1908)
);

OAI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1588),
.A2(n_1591),
.B(n_1595),
.Y(n_1909)
);

BUFx12f_ASAP7_75t_L g1910 ( 
.A(n_1628),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1612),
.A2(n_1585),
.B1(n_1657),
.B2(n_1601),
.Y(n_1911)
);

OR2x6_ASAP7_75t_L g1912 ( 
.A(n_1632),
.B(n_1561),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1708),
.Y(n_1913)
);

BUFx12f_ASAP7_75t_L g1914 ( 
.A(n_1680),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1660),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1620),
.B(n_1668),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1711),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1599),
.A2(n_1597),
.B1(n_1509),
.B2(n_1668),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_SL g1919 ( 
.A(n_1763),
.B(n_1614),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1638),
.B(n_1629),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1711),
.Y(n_1921)
);

OAI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1604),
.A2(n_1684),
.B(n_1679),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1711),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1542),
.B(n_1610),
.Y(n_1924)
);

BUFx2_ASAP7_75t_L g1925 ( 
.A(n_1614),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1674),
.A2(n_1646),
.B(n_1649),
.Y(n_1926)
);

OR2x6_ASAP7_75t_L g1927 ( 
.A(n_1493),
.B(n_1696),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1548),
.A2(n_1608),
.B1(n_1683),
.B2(n_1570),
.Y(n_1928)
);

A2O1A1Ixp33_ASAP7_75t_L g1929 ( 
.A1(n_1639),
.A2(n_1511),
.B(n_1530),
.C(n_1570),
.Y(n_1929)
);

OAI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1673),
.A2(n_1553),
.B(n_1551),
.Y(n_1930)
);

BUFx2_ASAP7_75t_SL g1931 ( 
.A(n_1715),
.Y(n_1931)
);

OAI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1647),
.A2(n_1652),
.B1(n_1645),
.B2(n_1546),
.Y(n_1932)
);

BUFx3_ASAP7_75t_L g1933 ( 
.A(n_1768),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1768),
.B(n_1656),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1659),
.B(n_1678),
.Y(n_1935)
);

OAI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1551),
.A2(n_1553),
.B(n_1642),
.Y(n_1936)
);

AOI22xp33_ASAP7_75t_L g1937 ( 
.A1(n_1633),
.A2(n_1546),
.B1(n_1634),
.B2(n_1587),
.Y(n_1937)
);

AOI21xp33_ASAP7_75t_L g1938 ( 
.A1(n_1676),
.A2(n_1681),
.B(n_1545),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1680),
.B(n_1563),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_SL g1940 ( 
.A(n_1653),
.B(n_1529),
.Y(n_1940)
);

A2O1A1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1583),
.A2(n_1607),
.B(n_1637),
.C(n_1535),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1682),
.A2(n_1686),
.B(n_1689),
.Y(n_1942)
);

INVx1_ASAP7_75t_SL g1943 ( 
.A(n_1690),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1522),
.A2(n_1547),
.B1(n_1653),
.B2(n_1681),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1772),
.B(n_1764),
.Y(n_1945)
);

CKINVDCx6p67_ASAP7_75t_R g1946 ( 
.A(n_1616),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_SL g1947 ( 
.A1(n_1690),
.A2(n_1564),
.B1(n_1541),
.B2(n_1661),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1687),
.A2(n_1772),
.B(n_1764),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1690),
.Y(n_1949)
);

AO21x2_ASAP7_75t_L g1950 ( 
.A1(n_1755),
.A2(n_1772),
.B(n_1764),
.Y(n_1950)
);

OAI21x1_ASAP7_75t_L g1951 ( 
.A1(n_1687),
.A2(n_1772),
.B(n_1755),
.Y(n_1951)
);

O2A1O1Ixp33_ASAP7_75t_SL g1952 ( 
.A1(n_1755),
.A2(n_1670),
.B(n_1499),
.C(n_1564),
.Y(n_1952)
);

OAI21x1_ASAP7_75t_L g1953 ( 
.A1(n_1687),
.A2(n_1755),
.B(n_1670),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1619),
.A2(n_1661),
.B1(n_1616),
.B2(n_1564),
.Y(n_1954)
);

OAI21x1_ASAP7_75t_L g1955 ( 
.A1(n_1670),
.A2(n_1500),
.B(n_1499),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1499),
.B(n_1500),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1661),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1773),
.A2(n_1316),
.B1(n_1307),
.B2(n_1538),
.Y(n_1958)
);

AO21x2_ASAP7_75t_L g1959 ( 
.A1(n_1698),
.A2(n_1704),
.B(n_1703),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1716),
.Y(n_1960)
);

BUFx3_ASAP7_75t_L g1961 ( 
.A(n_1716),
.Y(n_1961)
);

BUFx12f_ASAP7_75t_L g1962 ( 
.A(n_1566),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1693),
.Y(n_1963)
);

INVx1_ASAP7_75t_SL g1964 ( 
.A(n_1716),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1693),
.Y(n_1965)
);

OAI211xp5_ASAP7_75t_SL g1966 ( 
.A1(n_1579),
.A2(n_1363),
.B(n_1625),
.C(n_1573),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1568),
.B(n_1528),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1544),
.B(n_1761),
.Y(n_1968)
);

BUFx2_ASAP7_75t_L g1969 ( 
.A(n_1526),
.Y(n_1969)
);

AOI22xp33_ASAP7_75t_L g1970 ( 
.A1(n_1773),
.A2(n_1316),
.B1(n_1307),
.B2(n_1538),
.Y(n_1970)
);

CKINVDCx11_ASAP7_75t_R g1971 ( 
.A(n_1716),
.Y(n_1971)
);

OAI22xp5_ASAP7_75t_L g1972 ( 
.A1(n_1579),
.A2(n_1307),
.B1(n_1534),
.B2(n_1702),
.Y(n_1972)
);

INVx6_ASAP7_75t_L g1973 ( 
.A(n_1734),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1716),
.Y(n_1974)
);

AO21x1_ASAP7_75t_L g1975 ( 
.A1(n_1576),
.A2(n_1544),
.B(n_1593),
.Y(n_1975)
);

AO31x2_ASAP7_75t_L g1976 ( 
.A1(n_1510),
.A2(n_1703),
.A3(n_1704),
.B(n_1698),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1568),
.B(n_1528),
.Y(n_1977)
);

AOI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1773),
.A2(n_1316),
.B1(n_1307),
.B2(n_1538),
.Y(n_1978)
);

INVx4_ASAP7_75t_L g1979 ( 
.A(n_1873),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1966),
.B(n_1861),
.Y(n_1980)
);

BUFx3_ASAP7_75t_L g1981 ( 
.A(n_1873),
.Y(n_1981)
);

INVx1_ASAP7_75t_SL g1982 ( 
.A(n_1782),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1823),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1828),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1780),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1785),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1791),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1792),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1856),
.B(n_1861),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1799),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1800),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1807),
.Y(n_1992)
);

OR2x6_ASAP7_75t_L g1993 ( 
.A(n_1812),
.B(n_1873),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1809),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1812),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1862),
.B(n_1836),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1814),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1818),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1811),
.Y(n_1999)
);

CKINVDCx8_ASAP7_75t_R g2000 ( 
.A(n_1824),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1961),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1798),
.B(n_1797),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1835),
.B(n_1797),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1779),
.A2(n_1958),
.B1(n_1978),
.B2(n_1970),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1973),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1958),
.B(n_1970),
.Y(n_2006)
);

HB1xp67_ASAP7_75t_L g2007 ( 
.A(n_1902),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1902),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1827),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1858),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1963),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1973),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1886),
.B(n_1891),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1965),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1795),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1973),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1862),
.B(n_1854),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1885),
.Y(n_2018)
);

BUFx12f_ASAP7_75t_L g2019 ( 
.A(n_1971),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1961),
.Y(n_2020)
);

OR2x6_ASAP7_75t_L g2021 ( 
.A(n_1913),
.B(n_1822),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1795),
.Y(n_2022)
);

CKINVDCx6p67_ASAP7_75t_R g2023 ( 
.A(n_1971),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1888),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1820),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1863),
.B(n_1834),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1840),
.B(n_1788),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1866),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1897),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1878),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1884),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1822),
.B(n_1870),
.Y(n_2032)
);

AO21x2_ASAP7_75t_L g2033 ( 
.A1(n_1810),
.A2(n_1808),
.B(n_1956),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1784),
.B(n_1837),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1782),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1825),
.B(n_1838),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1815),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1815),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1848),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1846),
.B(n_1880),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1848),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1976),
.Y(n_2042)
);

OAI21x1_ASAP7_75t_SL g2043 ( 
.A1(n_1975),
.A2(n_1842),
.B(n_1865),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1857),
.Y(n_2044)
);

AND2x4_ASAP7_75t_L g2045 ( 
.A(n_1832),
.B(n_1864),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1839),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1846),
.B(n_1890),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_1832),
.B(n_1877),
.Y(n_2048)
);

HB1xp67_ASAP7_75t_L g2049 ( 
.A(n_1957),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1946),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1813),
.B(n_1860),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1976),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1787),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_1974),
.Y(n_2054)
);

AOI22xp33_ASAP7_75t_L g2055 ( 
.A1(n_1844),
.A2(n_1821),
.B1(n_1972),
.B2(n_1790),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1977),
.B(n_1967),
.Y(n_2056)
);

BUFx2_ASAP7_75t_L g2057 ( 
.A(n_1787),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1976),
.Y(n_2058)
);

NOR2xp67_ASAP7_75t_L g2059 ( 
.A(n_1960),
.B(n_1896),
.Y(n_2059)
);

AND2x6_ASAP7_75t_L g2060 ( 
.A(n_1843),
.B(n_1849),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1847),
.B(n_1826),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_SL g2062 ( 
.A1(n_1822),
.A2(n_1859),
.B1(n_1852),
.B2(n_1845),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_SL g2063 ( 
.A(n_1927),
.B(n_1931),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1847),
.B(n_1821),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1789),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1813),
.B(n_1860),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_1957),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1908),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1882),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1879),
.B(n_1881),
.Y(n_2070)
);

INVx1_ASAP7_75t_SL g2071 ( 
.A(n_1974),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1883),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_1803),
.B(n_1879),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1934),
.B(n_1853),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1905),
.Y(n_2075)
);

OR2x6_ASAP7_75t_L g2076 ( 
.A(n_1912),
.B(n_1850),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1875),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1925),
.Y(n_2078)
);

OR2x2_ASAP7_75t_L g2079 ( 
.A(n_1868),
.B(n_1892),
.Y(n_2079)
);

INVx1_ASAP7_75t_SL g2080 ( 
.A(n_1781),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1803),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1796),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_1914),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1915),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1796),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1796),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1855),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1906),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_1920),
.A2(n_1911),
.B1(n_1932),
.B2(n_1918),
.Y(n_2089)
);

OR2x6_ASAP7_75t_L g2090 ( 
.A(n_1912),
.B(n_1927),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1898),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1935),
.Y(n_2092)
);

AO21x2_ASAP7_75t_L g2093 ( 
.A1(n_1793),
.A2(n_1968),
.B(n_1833),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1960),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_1914),
.Y(n_2095)
);

BUFx4f_ASAP7_75t_SL g2096 ( 
.A(n_1962),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1904),
.Y(n_2097)
);

INVx4_ASAP7_75t_L g2098 ( 
.A(n_1802),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1895),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_L g2100 ( 
.A(n_1872),
.B(n_1920),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1817),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1817),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1829),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1829),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1910),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_1786),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1841),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1922),
.B(n_1911),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1841),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1867),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1867),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1950),
.B(n_1947),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_1786),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_1802),
.B(n_1816),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1794),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1804),
.B(n_1916),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1949),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_1816),
.B(n_1894),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2051),
.B(n_1955),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2051),
.B(n_1955),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1996),
.B(n_1893),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2072),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2007),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2066),
.B(n_1950),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2066),
.B(n_1947),
.Y(n_2125)
);

INVx2_ASAP7_75t_SL g2126 ( 
.A(n_1993),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2075),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_2090),
.B(n_1805),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1983),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1984),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2087),
.Y(n_2131)
);

OR2x2_ASAP7_75t_SL g2132 ( 
.A(n_2039),
.B(n_1869),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2008),
.Y(n_2133)
);

AND2x4_ASAP7_75t_SL g2134 ( 
.A(n_1979),
.B(n_1876),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2060),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_2077),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2027),
.B(n_1917),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_1999),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2003),
.B(n_1921),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_2100),
.A2(n_1918),
.B1(n_1804),
.B2(n_1912),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1985),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2108),
.B(n_1923),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2108),
.B(n_1923),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1986),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1987),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1988),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1990),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2036),
.B(n_1929),
.Y(n_2148)
);

INVxp67_ASAP7_75t_L g2149 ( 
.A(n_2010),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1991),
.Y(n_2150)
);

INVx2_ASAP7_75t_SL g2151 ( 
.A(n_1993),
.Y(n_2151)
);

INVx2_ASAP7_75t_SL g2152 ( 
.A(n_1993),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1992),
.Y(n_2153)
);

INVxp67_ASAP7_75t_SL g2154 ( 
.A(n_2013),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2056),
.B(n_1945),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2036),
.B(n_1929),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2056),
.B(n_1819),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1994),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2025),
.B(n_1932),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1997),
.Y(n_2160)
);

CKINVDCx8_ASAP7_75t_R g2161 ( 
.A(n_1993),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2047),
.B(n_1954),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_2090),
.B(n_1805),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_2049),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2047),
.B(n_1954),
.Y(n_2165)
);

HB1xp67_ASAP7_75t_L g2166 ( 
.A(n_2067),
.Y(n_2166)
);

AOI22xp33_ASAP7_75t_SL g2167 ( 
.A1(n_2100),
.A2(n_2063),
.B1(n_2034),
.B2(n_2006),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1998),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_2015),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_2022),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2006),
.B(n_1953),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_1981),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2009),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2112),
.B(n_1948),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2112),
.B(n_1951),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2002),
.B(n_1794),
.Y(n_2176)
);

INVx5_ASAP7_75t_L g2177 ( 
.A(n_1979),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_2078),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2011),
.Y(n_2179)
);

OR2x2_ASAP7_75t_L g2180 ( 
.A(n_2002),
.B(n_1959),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2014),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2084),
.Y(n_2182)
);

NAND2xp33_ASAP7_75t_R g2183 ( 
.A(n_2105),
.B(n_1876),
.Y(n_2183)
);

BUFx3_ASAP7_75t_L g2184 ( 
.A(n_1981),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2018),
.B(n_1907),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2024),
.B(n_1903),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2093),
.B(n_2040),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2026),
.B(n_1989),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2028),
.B(n_2017),
.Y(n_2189)
);

HB1xp67_ASAP7_75t_L g2190 ( 
.A(n_2037),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2038),
.B(n_1830),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2070),
.B(n_1830),
.Y(n_2192)
);

HB1xp67_ASAP7_75t_L g2193 ( 
.A(n_2001),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2061),
.B(n_1833),
.Y(n_2194)
);

BUFx2_ASAP7_75t_L g2195 ( 
.A(n_2060),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2029),
.B(n_1939),
.Y(n_2196)
);

INVx1_ASAP7_75t_SL g2197 ( 
.A(n_2001),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2069),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2068),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2046),
.Y(n_2200)
);

HB1xp67_ASAP7_75t_L g2201 ( 
.A(n_2053),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2065),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_2057),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2044),
.B(n_2091),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2092),
.B(n_1939),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2074),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1980),
.B(n_1939),
.Y(n_2207)
);

BUFx3_ASAP7_75t_L g2208 ( 
.A(n_1979),
.Y(n_2208)
);

NOR2xp67_ASAP7_75t_SL g2209 ( 
.A(n_2000),
.B(n_1851),
.Y(n_2209)
);

BUFx3_ASAP7_75t_L g2210 ( 
.A(n_2050),
.Y(n_2210)
);

OR2x6_ASAP7_75t_L g2211 ( 
.A(n_2021),
.B(n_1871),
.Y(n_2211)
);

INVx1_ASAP7_75t_SL g2212 ( 
.A(n_2094),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2171),
.B(n_2033),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2122),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2206),
.B(n_2034),
.Y(n_2215)
);

BUFx2_ASAP7_75t_L g2216 ( 
.A(n_2154),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2122),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2171),
.B(n_2033),
.Y(n_2218)
);

NAND2x1p5_ASAP7_75t_L g2219 ( 
.A(n_2177),
.B(n_1995),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2119),
.B(n_2042),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2131),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2119),
.B(n_2042),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2200),
.B(n_2089),
.Y(n_2223)
);

INVx4_ASAP7_75t_L g2224 ( 
.A(n_2177),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2123),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2182),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2129),
.Y(n_2227)
);

INVxp67_ASAP7_75t_L g2228 ( 
.A(n_2193),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_2135),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2128),
.B(n_2097),
.Y(n_2230)
);

HB1xp67_ASAP7_75t_L g2231 ( 
.A(n_2133),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2199),
.B(n_2089),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2130),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2127),
.Y(n_2234)
);

OR2x2_ASAP7_75t_L g2235 ( 
.A(n_2194),
.B(n_2081),
.Y(n_2235)
);

INVx3_ASAP7_75t_L g2236 ( 
.A(n_2135),
.Y(n_2236)
);

HB1xp67_ASAP7_75t_L g2237 ( 
.A(n_2169),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2202),
.Y(n_2238)
);

BUFx2_ASAP7_75t_L g2239 ( 
.A(n_2195),
.Y(n_2239)
);

BUFx3_ASAP7_75t_L g2240 ( 
.A(n_2172),
.Y(n_2240)
);

HB1xp67_ASAP7_75t_L g2241 ( 
.A(n_2170),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2120),
.B(n_2052),
.Y(n_2242)
);

BUFx2_ASAP7_75t_L g2243 ( 
.A(n_2195),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2120),
.B(n_2052),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_2136),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2141),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2124),
.B(n_2058),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2144),
.Y(n_2248)
);

OR2x2_ASAP7_75t_L g2249 ( 
.A(n_2157),
.B(n_2155),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2145),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2146),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2147),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_2174),
.B(n_2115),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2150),
.Y(n_2254)
);

INVx2_ASAP7_75t_SL g2255 ( 
.A(n_2177),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2153),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2174),
.B(n_2082),
.Y(n_2257)
);

NOR2xp67_ASAP7_75t_L g2258 ( 
.A(n_2177),
.B(n_2019),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2198),
.B(n_2148),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2156),
.B(n_2073),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2158),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2160),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2175),
.B(n_2085),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2168),
.B(n_2073),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2175),
.B(n_2086),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2173),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2179),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2181),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2191),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2178),
.Y(n_2270)
);

HB1xp67_ASAP7_75t_L g2271 ( 
.A(n_2138),
.Y(n_2271)
);

INVx2_ASAP7_75t_SL g2272 ( 
.A(n_2177),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2189),
.B(n_2055),
.Y(n_2273)
);

BUFx12f_ASAP7_75t_L g2274 ( 
.A(n_2208),
.Y(n_2274)
);

NAND2x1_ASAP7_75t_SL g2275 ( 
.A(n_2135),
.B(n_2041),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2137),
.B(n_2139),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2191),
.Y(n_2277)
);

INVx1_ASAP7_75t_SL g2278 ( 
.A(n_2197),
.Y(n_2278)
);

INVx1_ASAP7_75t_SL g2279 ( 
.A(n_2172),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2214),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_2249),
.B(n_2176),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2260),
.B(n_2159),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2214),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2217),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2217),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2234),
.Y(n_2286)
);

INVxp67_ASAP7_75t_L g2287 ( 
.A(n_2225),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2276),
.B(n_2190),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2257),
.B(n_2263),
.Y(n_2289)
);

NAND2x1_ASAP7_75t_SL g2290 ( 
.A(n_2258),
.B(n_2059),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2257),
.B(n_2187),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2276),
.B(n_2187),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_L g2293 ( 
.A(n_2273),
.B(n_2207),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2230),
.B(n_2128),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2249),
.B(n_2180),
.Y(n_2295)
);

NOR2x1p5_ASAP7_75t_L g2296 ( 
.A(n_2274),
.B(n_2023),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_2245),
.B(n_2231),
.Y(n_2297)
);

INVxp33_ASAP7_75t_L g2298 ( 
.A(n_2224),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2216),
.B(n_2192),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2265),
.B(n_2213),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_2240),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2213),
.B(n_2125),
.Y(n_2302)
);

OR2x2_ASAP7_75t_L g2303 ( 
.A(n_2216),
.B(n_2192),
.Y(n_2303)
);

INVx2_ASAP7_75t_SL g2304 ( 
.A(n_2240),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2238),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2237),
.B(n_2142),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2241),
.B(n_2142),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2218),
.B(n_2125),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2259),
.B(n_2143),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2218),
.B(n_2180),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2220),
.B(n_2162),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2270),
.B(n_2271),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2220),
.B(n_2162),
.Y(n_2313)
);

AND2x4_ASAP7_75t_L g2314 ( 
.A(n_2230),
.B(n_2163),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2238),
.Y(n_2315)
);

INVxp67_ASAP7_75t_L g2316 ( 
.A(n_2279),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2215),
.B(n_2264),
.Y(n_2317)
);

NOR2x1_ASAP7_75t_SL g2318 ( 
.A(n_2274),
.B(n_2076),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2232),
.B(n_2223),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2222),
.B(n_2165),
.Y(n_2320)
);

BUFx3_ASAP7_75t_L g2321 ( 
.A(n_2224),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2293),
.B(n_2228),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2300),
.B(n_2253),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2288),
.Y(n_2324)
);

OR2x2_ASAP7_75t_L g2325 ( 
.A(n_2310),
.B(n_2269),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2305),
.Y(n_2326)
);

AOI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2293),
.A2(n_2149),
.B1(n_2121),
.B2(n_1980),
.C(n_2164),
.Y(n_2327)
);

INVxp67_ASAP7_75t_SL g2328 ( 
.A(n_2299),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2280),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2300),
.B(n_2253),
.Y(n_2330)
);

NOR2x1p5_ASAP7_75t_L g2331 ( 
.A(n_2321),
.B(n_2224),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2282),
.A2(n_2167),
.B1(n_2140),
.B2(n_2004),
.Y(n_2332)
);

INVx2_ASAP7_75t_SL g2333 ( 
.A(n_2321),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2303),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2289),
.B(n_2222),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2283),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2289),
.B(n_2242),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2305),
.Y(n_2338)
);

OR2x2_ASAP7_75t_L g2339 ( 
.A(n_2310),
.B(n_2292),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2302),
.B(n_2235),
.Y(n_2340)
);

NAND4xp75_ASAP7_75t_L g2341 ( 
.A(n_2318),
.B(n_2272),
.C(n_2255),
.D(n_2126),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2315),
.Y(n_2342)
);

INVxp67_ASAP7_75t_L g2343 ( 
.A(n_2301),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_2294),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2284),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2291),
.B(n_2242),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2291),
.B(n_2244),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2312),
.Y(n_2348)
);

NAND4xp25_ASAP7_75t_L g2349 ( 
.A(n_2297),
.B(n_2004),
.C(n_2055),
.D(n_2062),
.Y(n_2349)
);

NAND2x1p5_ASAP7_75t_L g2350 ( 
.A(n_2296),
.B(n_2255),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2311),
.B(n_2244),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2302),
.B(n_2235),
.Y(n_2352)
);

OR2x2_ASAP7_75t_L g2353 ( 
.A(n_2281),
.B(n_2269),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2308),
.B(n_2221),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2287),
.B(n_2000),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2311),
.B(n_2247),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2315),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2285),
.Y(n_2358)
);

OR2x2_ASAP7_75t_L g2359 ( 
.A(n_2281),
.B(n_2277),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_2295),
.B(n_2277),
.Y(n_2360)
);

INVxp67_ASAP7_75t_SL g2361 ( 
.A(n_2298),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2286),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2334),
.B(n_2308),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_2323),
.B(n_2320),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2329),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2326),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2326),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2338),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2323),
.B(n_2320),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2338),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_2348),
.B(n_2316),
.Y(n_2371)
);

OAI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2350),
.A2(n_2298),
.B1(n_2161),
.B2(n_2301),
.Y(n_2372)
);

OAI221xp5_ASAP7_75t_L g2373 ( 
.A1(n_2332),
.A2(n_2319),
.B1(n_2317),
.B2(n_2307),
.C(n_2306),
.Y(n_2373)
);

AOI321xp33_ASAP7_75t_L g2374 ( 
.A1(n_2327),
.A2(n_2116),
.A3(n_2309),
.B1(n_2165),
.B2(n_2314),
.C(n_2294),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2329),
.Y(n_2375)
);

OR2x2_ASAP7_75t_L g2376 ( 
.A(n_2339),
.B(n_2295),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2336),
.Y(n_2377)
);

AOI211xp5_ASAP7_75t_SL g2378 ( 
.A1(n_2355),
.A2(n_2096),
.B(n_2290),
.C(n_2236),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2342),
.Y(n_2379)
);

INVxp67_ASAP7_75t_SL g2380 ( 
.A(n_2361),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2356),
.B(n_2313),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2342),
.Y(n_2382)
);

O2A1O1Ixp5_ASAP7_75t_L g2383 ( 
.A1(n_2328),
.A2(n_2294),
.B(n_2314),
.C(n_2230),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2333),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2357),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2357),
.Y(n_2386)
);

OAI322xp33_ASAP7_75t_L g2387 ( 
.A1(n_2339),
.A2(n_2278),
.A3(n_2188),
.B1(n_2304),
.B2(n_2248),
.C1(n_2267),
.C2(n_2233),
.Y(n_2387)
);

OAI22xp33_ASAP7_75t_SL g2388 ( 
.A1(n_2350),
.A2(n_2304),
.B1(n_2161),
.B2(n_2272),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2325),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_2322),
.B(n_2019),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2325),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2353),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2336),
.Y(n_2393)
);

OAI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2350),
.A2(n_2314),
.B1(n_2243),
.B2(n_2239),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2353),
.Y(n_2395)
);

NAND2x1_ASAP7_75t_SL g2396 ( 
.A(n_2344),
.B(n_2229),
.Y(n_2396)
);

OAI21xp33_ASAP7_75t_L g2397 ( 
.A1(n_2354),
.A2(n_2352),
.B(n_2340),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2345),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2345),
.Y(n_2399)
);

OAI211xp5_ASAP7_75t_L g2400 ( 
.A1(n_2349),
.A2(n_2071),
.B(n_1982),
.C(n_2054),
.Y(n_2400)
);

AND3x1_ASAP7_75t_L g2401 ( 
.A(n_2344),
.B(n_2023),
.C(n_1919),
.Y(n_2401)
);

OAI21xp5_ASAP7_75t_SL g2402 ( 
.A1(n_2378),
.A2(n_2134),
.B(n_2333),
.Y(n_2402)
);

OAI22xp5_ASAP7_75t_L g2403 ( 
.A1(n_2401),
.A2(n_2341),
.B1(n_2344),
.B2(n_2331),
.Y(n_2403)
);

NAND4xp25_ASAP7_75t_L g2404 ( 
.A(n_2374),
.B(n_2183),
.C(n_2054),
.D(n_2035),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2376),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2376),
.Y(n_2406)
);

OAI332xp33_ASAP7_75t_L g2407 ( 
.A1(n_2373),
.A2(n_1964),
.A3(n_2324),
.B1(n_2080),
.B2(n_2212),
.B3(n_2064),
.C1(n_1874),
.C2(n_2185),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2393),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2393),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2398),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2398),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2399),
.Y(n_2412)
);

INVx1_ASAP7_75t_SL g2413 ( 
.A(n_2384),
.Y(n_2413)
);

OAI211xp5_ASAP7_75t_SL g2414 ( 
.A1(n_2400),
.A2(n_2343),
.B(n_2186),
.C(n_2166),
.Y(n_2414)
);

OAI31xp33_ASAP7_75t_L g2415 ( 
.A1(n_2388),
.A2(n_2134),
.A3(n_2208),
.B(n_2239),
.Y(n_2415)
);

AOI21xp5_ASAP7_75t_L g2416 ( 
.A1(n_2383),
.A2(n_2076),
.B(n_2243),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2399),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2364),
.B(n_2330),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2392),
.B(n_2359),
.Y(n_2419)
);

INVx1_ASAP7_75t_SL g2420 ( 
.A(n_2390),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2366),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2365),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2397),
.B(n_2356),
.Y(n_2423)
);

OAI322xp33_ASAP7_75t_L g2424 ( 
.A1(n_2380),
.A2(n_2360),
.A3(n_2359),
.B1(n_2362),
.B2(n_2358),
.C1(n_2246),
.C2(n_2226),
.Y(n_2424)
);

OAI211xp5_ASAP7_75t_SL g2425 ( 
.A1(n_2371),
.A2(n_2088),
.B(n_2204),
.C(n_1944),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_2372),
.B(n_2096),
.Y(n_2426)
);

AOI21xp5_ASAP7_75t_L g2427 ( 
.A1(n_2387),
.A2(n_2394),
.B(n_2363),
.Y(n_2427)
);

OAI211xp5_ASAP7_75t_L g2428 ( 
.A1(n_2426),
.A2(n_2035),
.B(n_2396),
.C(n_1900),
.Y(n_2428)
);

OAI22xp5_ASAP7_75t_L g2429 ( 
.A1(n_2427),
.A2(n_2341),
.B1(n_2381),
.B2(n_2369),
.Y(n_2429)
);

AOI21xp33_ASAP7_75t_L g2430 ( 
.A1(n_2426),
.A2(n_2020),
.B(n_1783),
.Y(n_2430)
);

AOI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_2414),
.A2(n_2416),
.B(n_2403),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2421),
.Y(n_2432)
);

AOI22xp5_ASAP7_75t_L g2433 ( 
.A1(n_2414),
.A2(n_2391),
.B1(n_2395),
.B2(n_2392),
.Y(n_2433)
);

AOI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2402),
.A2(n_2076),
.B(n_2375),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2405),
.Y(n_2435)
);

NAND3xp33_ASAP7_75t_L g2436 ( 
.A(n_2415),
.B(n_2377),
.C(n_1944),
.Y(n_2436)
);

AOI221xp5_ASAP7_75t_L g2437 ( 
.A1(n_2424),
.A2(n_2391),
.B1(n_2227),
.B2(n_2252),
.C(n_2251),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2406),
.B(n_2423),
.Y(n_2438)
);

AOI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2413),
.A2(n_2076),
.B(n_2370),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2422),
.Y(n_2440)
);

OAI22x1_ASAP7_75t_SL g2441 ( 
.A1(n_2420),
.A2(n_1900),
.B1(n_2105),
.B2(n_1831),
.Y(n_2441)
);

OAI221xp5_ASAP7_75t_L g2442 ( 
.A1(n_2404),
.A2(n_2425),
.B1(n_2396),
.B2(n_2410),
.C(n_2409),
.Y(n_2442)
);

OAI222xp33_ASAP7_75t_L g2443 ( 
.A1(n_2419),
.A2(n_2389),
.B1(n_2395),
.B2(n_2364),
.C1(n_2369),
.C2(n_2211),
.Y(n_2443)
);

AOI221xp5_ASAP7_75t_L g2444 ( 
.A1(n_2407),
.A2(n_2250),
.B1(n_2261),
.B2(n_2256),
.C(n_2254),
.Y(n_2444)
);

OAI222xp33_ASAP7_75t_L g2445 ( 
.A1(n_2418),
.A2(n_2389),
.B1(n_2211),
.B2(n_2360),
.C1(n_2337),
.C2(n_2335),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2408),
.B(n_2351),
.Y(n_2446)
);

O2A1O1Ixp33_ASAP7_75t_L g2447 ( 
.A1(n_2425),
.A2(n_2095),
.B(n_2083),
.C(n_2043),
.Y(n_2447)
);

AOI311xp33_ASAP7_75t_L g2448 ( 
.A1(n_2411),
.A2(n_2382),
.A3(n_2385),
.B(n_2379),
.C(n_2370),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_SL g2449 ( 
.A(n_2421),
.B(n_1962),
.Y(n_2449)
);

OAI21xp5_ASAP7_75t_L g2450 ( 
.A1(n_2412),
.A2(n_2417),
.B(n_2219),
.Y(n_2450)
);

O2A1O1Ixp33_ASAP7_75t_L g2451 ( 
.A1(n_2426),
.A2(n_2020),
.B(n_2203),
.C(n_2201),
.Y(n_2451)
);

AOI211xp5_ASAP7_75t_L g2452 ( 
.A1(n_2426),
.A2(n_2209),
.B(n_2184),
.C(n_1899),
.Y(n_2452)
);

OAI211xp5_ASAP7_75t_L g2453 ( 
.A1(n_2426),
.A2(n_2094),
.B(n_2031),
.C(n_2275),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2405),
.B(n_2351),
.Y(n_2454)
);

OAI221xp5_ASAP7_75t_L g2455 ( 
.A1(n_2415),
.A2(n_2385),
.B1(n_2382),
.B2(n_2379),
.C(n_1940),
.Y(n_2455)
);

INVx2_ASAP7_75t_SL g2456 ( 
.A(n_2441),
.Y(n_2456)
);

HB1xp67_ASAP7_75t_L g2457 ( 
.A(n_2435),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2440),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2438),
.B(n_2366),
.Y(n_2459)
);

NAND5xp2_ASAP7_75t_L g2460 ( 
.A(n_2431),
.B(n_2219),
.C(n_1937),
.D(n_1930),
.E(n_1901),
.Y(n_2460)
);

NAND5xp2_ASAP7_75t_L g2461 ( 
.A(n_2452),
.B(n_2219),
.C(n_1937),
.D(n_1889),
.E(n_1969),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_SL g2462 ( 
.A(n_2451),
.B(n_1889),
.Y(n_2462)
);

NOR3xp33_ASAP7_75t_L g2463 ( 
.A(n_2429),
.B(n_1801),
.C(n_1831),
.Y(n_2463)
);

NOR3xp33_ASAP7_75t_L g2464 ( 
.A(n_2428),
.B(n_1806),
.C(n_1928),
.Y(n_2464)
);

OAI21xp33_ASAP7_75t_L g2465 ( 
.A1(n_2442),
.A2(n_2368),
.B(n_2367),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2432),
.Y(n_2466)
);

NAND3xp33_ASAP7_75t_SL g2467 ( 
.A(n_2437),
.B(n_2113),
.C(n_2106),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2453),
.B(n_2367),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_SL g2469 ( 
.A(n_2437),
.B(n_2184),
.Y(n_2469)
);

NOR3xp33_ASAP7_75t_L g2470 ( 
.A(n_2455),
.B(n_1938),
.C(n_1909),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2446),
.Y(n_2471)
);

HB1xp67_ASAP7_75t_L g2472 ( 
.A(n_2433),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2444),
.B(n_2335),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2454),
.Y(n_2474)
);

INVx1_ASAP7_75t_SL g2475 ( 
.A(n_2449),
.Y(n_2475)
);

HB1xp67_ASAP7_75t_L g2476 ( 
.A(n_2457),
.Y(n_2476)
);

AND5x1_ASAP7_75t_L g2477 ( 
.A(n_2463),
.B(n_2439),
.C(n_2434),
.D(n_2447),
.E(n_2444),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_2456),
.B(n_2443),
.Y(n_2478)
);

NOR2x1_ASAP7_75t_L g2479 ( 
.A(n_2467),
.B(n_1876),
.Y(n_2479)
);

NOR3xp33_ASAP7_75t_L g2480 ( 
.A(n_2460),
.B(n_2445),
.C(n_2430),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2458),
.Y(n_2481)
);

NOR2x1_ASAP7_75t_L g2482 ( 
.A(n_2469),
.B(n_2436),
.Y(n_2482)
);

OAI211xp5_ASAP7_75t_SL g2483 ( 
.A1(n_2456),
.A2(n_2472),
.B(n_2475),
.C(n_2465),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2466),
.Y(n_2484)
);

NOR3xp33_ASAP7_75t_L g2485 ( 
.A(n_2461),
.B(n_2450),
.C(n_2050),
.Y(n_2485)
);

AND5x1_ASAP7_75t_L g2486 ( 
.A(n_2462),
.B(n_2448),
.C(n_1952),
.D(n_1910),
.E(n_1941),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2474),
.Y(n_2487)
);

NOR2x1_ASAP7_75t_L g2488 ( 
.A(n_2469),
.B(n_2050),
.Y(n_2488)
);

NAND3xp33_ASAP7_75t_SL g2489 ( 
.A(n_2464),
.B(n_2468),
.C(n_2473),
.Y(n_2489)
);

AOI211xp5_ASAP7_75t_L g2490 ( 
.A1(n_2470),
.A2(n_2209),
.B(n_2210),
.C(n_2151),
.Y(n_2490)
);

NOR3xp33_ASAP7_75t_SL g2491 ( 
.A(n_2468),
.B(n_2030),
.C(n_1936),
.Y(n_2491)
);

AND3x1_ASAP7_75t_L g2492 ( 
.A(n_2466),
.B(n_2151),
.C(n_2126),
.Y(n_2492)
);

NAND3xp33_ASAP7_75t_L g2493 ( 
.A(n_2471),
.B(n_2102),
.C(n_2101),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2476),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2484),
.Y(n_2495)
);

OAI322xp33_ASAP7_75t_L g2496 ( 
.A1(n_2478),
.A2(n_2487),
.A3(n_2481),
.B1(n_2483),
.B2(n_2477),
.C1(n_2489),
.C2(n_2471),
.Y(n_2496)
);

NOR3xp33_ASAP7_75t_L g2497 ( 
.A(n_2489),
.B(n_2459),
.C(n_1924),
.Y(n_2497)
);

OR2x2_ASAP7_75t_L g2498 ( 
.A(n_2493),
.B(n_2337),
.Y(n_2498)
);

OR2x2_ASAP7_75t_L g2499 ( 
.A(n_2480),
.B(n_2346),
.Y(n_2499)
);

NOR3x1_ASAP7_75t_L g2500 ( 
.A(n_2479),
.B(n_2152),
.C(n_2032),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2482),
.B(n_2330),
.Y(n_2501)
);

NOR3xp33_ASAP7_75t_L g2502 ( 
.A(n_2488),
.B(n_1926),
.C(n_1943),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2491),
.Y(n_2503)
);

NOR2x1_ASAP7_75t_L g2504 ( 
.A(n_2486),
.B(n_2021),
.Y(n_2504)
);

NOR3x2_ASAP7_75t_L g2505 ( 
.A(n_2485),
.B(n_2079),
.C(n_2021),
.Y(n_2505)
);

NAND4xp75_ASAP7_75t_L g2506 ( 
.A(n_2492),
.B(n_2152),
.C(n_2005),
.D(n_2016),
.Y(n_2506)
);

OR3x2_ASAP7_75t_L g2507 ( 
.A(n_2503),
.B(n_2490),
.C(n_2104),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2494),
.Y(n_2508)
);

AND2x4_ASAP7_75t_L g2509 ( 
.A(n_2494),
.B(n_2346),
.Y(n_2509)
);

OR2x2_ASAP7_75t_L g2510 ( 
.A(n_2499),
.B(n_2347),
.Y(n_2510)
);

NOR3xp33_ASAP7_75t_L g2511 ( 
.A(n_2496),
.B(n_2012),
.C(n_2005),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2495),
.B(n_2497),
.Y(n_2512)
);

AOI22xp5_ASAP7_75t_L g2513 ( 
.A1(n_2504),
.A2(n_2021),
.B1(n_2211),
.B2(n_2210),
.Y(n_2513)
);

NAND3xp33_ASAP7_75t_L g2514 ( 
.A(n_2502),
.B(n_2107),
.C(n_2103),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2501),
.B(n_2347),
.Y(n_2515)
);

INVx1_ASAP7_75t_SL g2516 ( 
.A(n_2505),
.Y(n_2516)
);

NOR2x1_ASAP7_75t_L g2517 ( 
.A(n_2506),
.B(n_1927),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2508),
.Y(n_2518)
);

OAI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2507),
.A2(n_2498),
.B1(n_2500),
.B2(n_2132),
.Y(n_2519)
);

NAND3x1_ASAP7_75t_L g2520 ( 
.A(n_2512),
.B(n_2511),
.C(n_2517),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2509),
.Y(n_2521)
);

OAI211xp5_ASAP7_75t_SL g2522 ( 
.A1(n_2516),
.A2(n_2117),
.B(n_2110),
.C(n_2111),
.Y(n_2522)
);

AOI21xp33_ASAP7_75t_L g2523 ( 
.A1(n_2510),
.A2(n_2109),
.B(n_2016),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2515),
.B(n_2368),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2514),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2513),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2516),
.B(n_2262),
.Y(n_2527)
);

AOI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2516),
.A2(n_2211),
.B1(n_2045),
.B2(n_2048),
.Y(n_2528)
);

OAI21x1_ASAP7_75t_L g2529 ( 
.A1(n_2520),
.A2(n_2012),
.B(n_2275),
.Y(n_2529)
);

AOI21xp5_ASAP7_75t_L g2530 ( 
.A1(n_2518),
.A2(n_1887),
.B(n_1942),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2521),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2527),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2525),
.B(n_2266),
.Y(n_2533)
);

AO21x1_ASAP7_75t_L g2534 ( 
.A1(n_2526),
.A2(n_2098),
.B(n_2268),
.Y(n_2534)
);

A2O1A1Ixp33_ASAP7_75t_L g2535 ( 
.A1(n_2531),
.A2(n_2522),
.B(n_2528),
.C(n_2519),
.Y(n_2535)
);

OAI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_2532),
.A2(n_2524),
.B1(n_2523),
.B2(n_2132),
.Y(n_2536)
);

OR2x6_ASAP7_75t_L g2537 ( 
.A(n_2534),
.B(n_1933),
.Y(n_2537)
);

AO21x2_ASAP7_75t_L g2538 ( 
.A1(n_2533),
.A2(n_2205),
.B(n_2196),
.Y(n_2538)
);

OA22x2_ASAP7_75t_L g2539 ( 
.A1(n_2529),
.A2(n_2386),
.B1(n_2012),
.B2(n_2098),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2530),
.B(n_2386),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_L g2541 ( 
.A(n_2535),
.B(n_2098),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2536),
.Y(n_2542)
);

AOI21xp33_ASAP7_75t_L g2543 ( 
.A1(n_2537),
.A2(n_2539),
.B(n_2540),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2542),
.B(n_2541),
.Y(n_2544)
);

AOI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2543),
.A2(n_2538),
.B1(n_2118),
.B2(n_2114),
.Y(n_2545)
);

OR2x6_ASAP7_75t_L g2546 ( 
.A(n_2544),
.B(n_2545),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2546),
.B(n_2229),
.Y(n_2547)
);

AOI22xp33_ASAP7_75t_L g2548 ( 
.A1(n_2547),
.A2(n_2236),
.B1(n_2229),
.B2(n_2099),
.Y(n_2548)
);


endmodule