module fake_jpeg_139_n_449 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_449);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_449;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_47),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g141 ( 
.A(n_52),
.Y(n_141)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_55),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_58),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_59),
.B(n_62),
.Y(n_125)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_23),
.B(n_8),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_64),
.B(n_66),
.Y(n_128)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_72),
.Y(n_132)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_8),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_34),
.B(n_8),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_38),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_79),
.B(n_88),
.Y(n_120)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_39),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_33),
.B(n_7),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_18),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_38),
.CON(n_103),
.SN(n_103)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_103),
.B(n_100),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_112),
.B(n_24),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_40),
.B(n_29),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_26),
.Y(n_153)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_53),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_36),
.B1(n_20),
.B2(n_28),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_86),
.A2(n_65),
.B1(n_54),
.B2(n_63),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_85),
.B1(n_70),
.B2(n_71),
.Y(n_159)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_44),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_41),
.Y(n_144)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_149),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_78),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_163),
.Y(n_202)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g208 ( 
.A(n_148),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_90),
.Y(n_149)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_154),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_76),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_45),
.B1(n_61),
.B2(n_56),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_155),
.A2(n_161),
.B1(n_173),
.B2(n_111),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_159),
.A2(n_160),
.B1(n_175),
.B2(n_177),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_124),
.A2(n_76),
.B1(n_29),
.B2(n_32),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_73),
.B1(n_58),
.B2(n_18),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_77),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_186),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_32),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_164),
.B(n_176),
.Y(n_195)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

BUFx2_ASAP7_75t_R g168 ( 
.A(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_178),
.Y(n_211)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

BUFx8_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_97),
.A2(n_36),
.B1(n_28),
.B2(n_77),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_114),
.B(n_80),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_180),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_109),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_131),
.B(n_28),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_183),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_163),
.B(n_170),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_140),
.B(n_83),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_96),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_95),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_126),
.B(n_9),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_97),
.B(n_69),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_172),
.C(n_147),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_205),
.C(n_217),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_136),
.B(n_103),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_204),
.B(n_212),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_122),
.B(n_116),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_99),
.C(n_134),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_138),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_159),
.A2(n_130),
.B(n_133),
.C(n_142),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_213),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_96),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_159),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_204),
.B1(n_214),
.B2(n_202),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_223),
.B1(n_224),
.B2(n_218),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_184),
.B1(n_159),
.B2(n_173),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_150),
.B1(n_107),
.B2(n_200),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_SL g261 ( 
.A1(n_222),
.A2(n_233),
.B(n_174),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_166),
.B1(n_178),
.B2(n_169),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_146),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

AND2x6_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_213),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

INVx13_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_231),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_235),
.Y(n_244)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_209),
.A2(n_152),
.B1(n_171),
.B2(n_158),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_240),
.Y(n_251)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_162),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_205),
.C(n_199),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_216),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_239),
.Y(n_250)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_148),
.Y(n_240)
);

NAND2x1p5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_162),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_197),
.B(n_190),
.Y(n_260)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_242),
.A2(n_190),
.B1(n_197),
.B2(n_146),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_201),
.B1(n_194),
.B2(n_215),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_243),
.A2(n_249),
.B1(n_257),
.B2(n_261),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_247),
.A2(n_253),
.B1(n_262),
.B2(n_239),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_248),
.A2(n_260),
.B(n_264),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_224),
.A2(n_201),
.B1(n_215),
.B2(n_203),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_219),
.A2(n_203),
.B1(n_216),
.B2(n_207),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_226),
.B1(n_241),
.B2(n_236),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_195),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_256),
.C(n_259),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_238),
.A2(n_213),
.B1(n_195),
.B2(n_199),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_199),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_200),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_236),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_177),
.B(n_168),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_188),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_241),
.C(n_232),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_240),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_268),
.B(n_269),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_220),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_276),
.C(n_279),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_272),
.B(n_273),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_226),
.B(n_248),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_274),
.A2(n_243),
.B(n_260),
.Y(n_296)
);

INVx13_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_254),
.B1(n_246),
.B2(n_258),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_250),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_223),
.Y(n_278)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_233),
.C(n_188),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_251),
.B(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_283),
.B(n_285),
.Y(n_303)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_244),
.Y(n_284)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_189),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_286),
.Y(n_310)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_189),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_289),
.B(n_266),
.Y(n_307)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_290),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_289),
.C(n_268),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_300),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_271),
.A2(n_247),
.B(n_233),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_299),
.B(n_296),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_274),
.A2(n_271),
.B(n_282),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_278),
.B1(n_277),
.B2(n_279),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_305),
.A2(n_246),
.B1(n_230),
.B2(n_275),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_233),
.B(n_256),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_267),
.C(n_272),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_254),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_269),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_242),
.Y(n_312)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_312),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_235),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_315),
.B(n_141),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_267),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_321),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_L g346 ( 
.A1(n_319),
.A2(n_299),
.B(n_309),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_297),
.A2(n_301),
.B1(n_298),
.B2(n_291),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_320),
.A2(n_327),
.B1(n_302),
.B2(n_314),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_270),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_326),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_285),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_324),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_283),
.Y(n_325)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_325),
.Y(n_354)
);

BUFx12f_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_287),
.B1(n_286),
.B2(n_290),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_330),
.B1(n_293),
.B2(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_294),
.Y(n_329)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_305),
.A2(n_275),
.B1(n_229),
.B2(n_191),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_333),
.C(n_334),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_129),
.C(n_101),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_117),
.C(n_165),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_292),
.B(n_165),
.C(n_93),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_339),
.C(n_310),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_311),
.B(n_208),
.Y(n_337)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_302),
.B(n_309),
.C(n_298),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_355),
.B1(n_361),
.B2(n_326),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_329),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_348),
.Y(n_372)
);

XNOR2x1_ASAP7_75t_SL g345 ( 
.A(n_316),
.B(n_294),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_350),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_346),
.A2(n_323),
.B(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_336),
.A2(n_303),
.B1(n_312),
.B2(n_295),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_330),
.A2(n_303),
.B1(n_295),
.B2(n_229),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_356),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_206),
.C(n_231),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_360),
.C(n_362),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_331),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_353),
.B(n_323),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_320),
.A2(n_206),
.B1(n_150),
.B2(n_157),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_318),
.A2(n_206),
.B1(n_208),
.B2(n_231),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_358),
.B(n_335),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_315),
.B(n_208),
.C(n_107),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_137),
.B1(n_138),
.B2(n_151),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_333),
.B(n_339),
.C(n_332),
.Y(n_362)
);

BUFx12_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_367),
.Y(n_383)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_354),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_374),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_371),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_370),
.A2(n_361),
.B1(n_343),
.B2(n_352),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_338),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_334),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_373),
.B(n_375),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_344),
.B(n_326),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_357),
.A2(n_326),
.B1(n_156),
.B2(n_151),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_376),
.A2(n_378),
.B1(n_380),
.B2(n_363),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_186),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_381),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_346),
.A2(n_359),
.B1(n_347),
.B2(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_14),
.Y(n_395)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_385),
.A2(n_388),
.B1(n_396),
.B2(n_379),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_380),
.A2(n_343),
.B1(n_353),
.B2(n_341),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_387),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_341),
.C(n_137),
.Y(n_387)
);

AOI211xp5_ASAP7_75t_L g388 ( 
.A1(n_366),
.A2(n_365),
.B(n_364),
.C(n_372),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_377),
.B(n_156),
.C(n_123),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_390),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_378),
.A2(n_121),
.B1(n_115),
.B2(n_119),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_92),
.C(n_60),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_391),
.B(n_13),
.Y(n_410)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_395),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_364),
.A2(n_7),
.B1(n_12),
.B2(n_3),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_365),
.A2(n_9),
.B(n_12),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_6),
.B(n_11),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_398),
.B(n_368),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_402),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_371),
.Y(n_402)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_403),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_388),
.A2(n_376),
.B1(n_374),
.B2(n_4),
.Y(n_404)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_393),
.A2(n_9),
.B(n_12),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_408),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_392),
.B(n_394),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_406),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_11),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_397),
.A2(n_13),
.B(n_4),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_10),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_396),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_412),
.B(n_392),
.Y(n_413)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_413),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_422),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_387),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_407),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_399),
.A2(n_391),
.B(n_389),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_416),
.A2(n_403),
.B(n_404),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_4),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_401),
.B(n_5),
.C(n_10),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_424),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_427),
.B(n_429),
.Y(n_434)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_426),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_417),
.B(n_408),
.Y(n_427)
);

BUFx24_ASAP7_75t_SL g429 ( 
.A(n_419),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_420),
.A2(n_5),
.B(n_10),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_430),
.A2(n_418),
.B(n_421),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_5),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_431),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_435),
.B(n_11),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_433),
.A2(n_420),
.B1(n_416),
.B2(n_10),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_437),
.B(n_428),
.C(n_432),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_426),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_439),
.A2(n_0),
.B1(n_1),
.B2(n_436),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_440),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_441),
.A2(n_442),
.B(n_443),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_11),
.C(n_0),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_434),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_444),
.C(n_0),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_447),
.A2(n_0),
.B(n_1),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_0),
.Y(n_449)
);


endmodule