module fake_jpeg_20435_n_237 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_237);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_17),
.B1(n_11),
.B2(n_23),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_36),
.B1(n_26),
.B2(n_12),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_54),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_32),
.Y(n_60)
);

BUFx2_ASAP7_75t_SL g46 ( 
.A(n_39),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_32),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_31),
.B1(n_17),
.B2(n_11),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_52),
.B1(n_55),
.B2(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_26),
.B1(n_27),
.B2(n_25),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_26),
.C(n_15),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_11),
.B1(n_28),
.B2(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_60),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_40),
.C(n_35),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_63),
.C(n_68),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_40),
.C(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_26),
.C(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_11),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_77),
.Y(n_104)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_43),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_88),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_52),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_84),
.B(n_87),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_46),
.B(n_36),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_91),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_83),
.B1(n_42),
.B2(n_64),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_90),
.B(n_100),
.C(n_53),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_56),
.B(n_57),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_42),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_71),
.B1(n_60),
.B2(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_30),
.B1(n_39),
.B2(n_27),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_98),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_63),
.B(n_68),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_85),
.B1(n_87),
.B2(n_81),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_79),
.B1(n_74),
.B2(n_88),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_30),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_53),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_116),
.B1(n_91),
.B2(n_37),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_111),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_113),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_96),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_34),
.B(n_30),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_62),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_128),
.C(n_127),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_62),
.B1(n_58),
.B2(n_49),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_16),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_119),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_123),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_12),
.B1(n_37),
.B2(n_25),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_91),
.B1(n_39),
.B2(n_44),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_13),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_30),
.B1(n_24),
.B2(n_22),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_44),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_16),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_16),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_89),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_100),
.C(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_124),
.C(n_119),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_131),
.A2(n_139),
.B(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_21),
.B1(n_12),
.B2(n_18),
.Y(n_134)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_19),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_23),
.B1(n_15),
.B2(n_21),
.Y(n_138)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_129),
.B(n_21),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_15),
.B1(n_23),
.B2(n_22),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_152),
.B1(n_121),
.B2(n_119),
.Y(n_155)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_10),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_148),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_108),
.B1(n_120),
.B2(n_126),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_24),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_34),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_151),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_159),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_22),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_135),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_170),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_22),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_147),
.B(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_20),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_154),
.C(n_170),
.Y(n_171)
);

BUFx4f_ASAP7_75t_SL g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_20),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_183),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_136),
.C(n_150),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_167),
.C(n_14),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_181),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_132),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_149),
.B1(n_145),
.B2(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_164),
.B1(n_150),
.B2(n_144),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_159),
.B(n_165),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_131),
.B(n_151),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_20),
.B(n_13),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_174),
.B1(n_179),
.B2(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_133),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_191),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_168),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_184),
.A2(n_163),
.B1(n_167),
.B2(n_152),
.C(n_9),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_193),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_197),
.Y(n_204)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_14),
.A3(n_20),
.B1(n_13),
.B2(n_19),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_178),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_200),
.B(n_203),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_175),
.B1(n_196),
.B2(n_194),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_201),
.A2(n_195),
.B1(n_2),
.B2(n_3),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_207),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_178),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_8),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_182),
.B1(n_179),
.B2(n_10),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_214),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_1),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_213),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_13),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_13),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_19),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_8),
.B(n_2),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_201),
.B(n_8),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_222),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_210),
.B(n_13),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_212),
.C(n_214),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_19),
.C(n_5),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_213),
.A3(n_215),
.B1(n_13),
.B2(n_19),
.C1(n_6),
.C2(n_7),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_227),
.B(n_4),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_225),
.A2(n_220),
.B(n_222),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_230),
.B(n_228),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_232),
.C(n_226),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_233),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_19),
.B1(n_6),
.B2(n_7),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_19),
.C(n_4),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_4),
.Y(n_237)
);


endmodule