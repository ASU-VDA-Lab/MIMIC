module real_jpeg_5464_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_10;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_11;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_65;
wire n_33;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_1),
.A2(n_39),
.B1(n_83),
.B2(n_86),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_1),
.A2(n_39),
.B1(n_96),
.B2(n_100),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_2),
.B(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_2),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_2),
.A2(n_71),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_2),
.A2(n_118),
.B(n_119),
.C(n_125),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_2),
.B(n_139),
.C(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_2),
.A2(n_71),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_2),
.B(n_65),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_2),
.B(n_16),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_5),
.Y(n_129)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_5),
.Y(n_162)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_5),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_25),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_8),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_133),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_131),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_88),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_12),
.B(n_88),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_51),
.C(n_61),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_13),
.A2(n_14),
.B1(n_51),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_33),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_24),
.Y(n_15)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_16),
.B(n_34),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_16)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_21),
.Y(n_167)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_42),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_27),
.B(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_27),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_29),
.Y(n_147)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_42),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_54),
.B1(n_57),
.B2(n_59),
.Y(n_53)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_42),
.B(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_51),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_52),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_54),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_75),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_77),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_67),
.B(n_77),
.Y(n_176)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_71),
.A2(n_120),
.B(n_123),
.Y(n_119)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_76),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_77),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_82),
.B(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_116),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_152),
.B(n_184),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_149),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_137),
.B1(n_142),
.B2(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_168),
.B(n_183),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_177),
.B(n_182),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_181),
.Y(n_182)
);


endmodule