module fake_jpeg_19252_n_263 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_263);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_11),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_34),
.B1(n_24),
.B2(n_32),
.Y(n_42)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_24),
.B1(n_26),
.B2(n_18),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_24),
.B1(n_32),
.B2(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_56),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_48),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_24),
.B1(n_18),
.B2(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_49),
.Y(n_68)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_SL g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_54),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_26),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_30),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_12),
.B(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_18),
.B1(n_38),
.B2(n_21),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_29),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_47),
.B1(n_17),
.B2(n_23),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_70),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_75),
.Y(n_81)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_84),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_42),
.B1(n_48),
.B2(n_45),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_93),
.B1(n_74),
.B2(n_73),
.Y(n_113)
);

OAI21x1_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_57),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_88),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_67),
.B(n_31),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_58),
.C(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_94),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_53),
.Y(n_95)
);

AO21x2_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_77),
.B(n_71),
.Y(n_97)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_76),
.B1(n_66),
.B2(n_67),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_109),
.B1(n_114),
.B2(n_93),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g103 ( 
.A(n_94),
.Y(n_103)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_106),
.Y(n_127)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_85),
.B(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_64),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_67),
.B1(n_74),
.B2(n_73),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_110),
.B(n_112),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_113),
.A2(n_96),
.B1(n_90),
.B2(n_111),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_73),
.B1(n_75),
.B2(n_47),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_22),
.B(n_16),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_91),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_29),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_108),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_134),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_126),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_125),
.B1(n_131),
.B2(n_133),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_159)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_88),
.C(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_81),
.C(n_55),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_137),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_21),
.B1(n_65),
.B2(n_69),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_113),
.B1(n_97),
.B2(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_139),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_31),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_19),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_69),
.C(n_29),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_28),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_97),
.B(n_53),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_19),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_19),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_106),
.B(n_97),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_165),
.B1(n_123),
.B2(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_103),
.B1(n_116),
.B2(n_69),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_153),
.B1(n_156),
.B2(n_12),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_9),
.B(n_1),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_152),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_16),
.B(n_23),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_21),
.B1(n_13),
.B2(n_15),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_161),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_17),
.B1(n_13),
.B2(n_15),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_159),
.A2(n_160),
.B1(n_13),
.B2(n_11),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_29),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_140),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_122),
.B(n_132),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_167),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_117),
.A2(n_6),
.B(n_2),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_131),
.B1(n_129),
.B2(n_126),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_178),
.C(n_182),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_165),
.B(n_158),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_137),
.B1(n_17),
.B2(n_15),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_175),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_13),
.B1(n_16),
.B2(n_11),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_156),
.B1(n_151),
.B2(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_16),
.B1(n_12),
.B2(n_30),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_183),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_148),
.B(n_20),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_29),
.C(n_30),
.Y(n_182)
);

AO21x2_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_27),
.B(n_28),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_29),
.C(n_27),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_154),
.C(n_163),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_189),
.B(n_144),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_204),
.B1(n_159),
.B2(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_186),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_166),
.B(n_180),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_178),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_170),
.C(n_187),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_29),
.C(n_20),
.Y(n_216)
);

OAI221xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_167),
.B1(n_152),
.B2(n_149),
.C(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_173),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_209),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_208),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_155),
.Y(n_209)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_211),
.A2(n_212),
.B1(n_197),
.B2(n_194),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_183),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_183),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_20),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_192),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g220 ( 
.A(n_214),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_220),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_226),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_188),
.C(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_217),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_196),
.C(n_193),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_207),
.A2(n_195),
.B(n_200),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_193),
.B(n_191),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_197),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_231),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_194),
.C(n_199),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_235),
.Y(n_244)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_234),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_191),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_225),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_237),
.C(n_218),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_6),
.C(n_2),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_6),
.B1(n_2),
.B2(n_3),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_4),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_245),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_228),
.B(n_3),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_242),
.A2(n_5),
.B(n_7),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_7),
.B1(n_4),
.B2(n_5),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

AOI321xp33_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_7),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_10),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_5),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_239),
.C(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_8),
.C(n_9),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_249),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_239),
.B(n_250),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_257),
.B1(n_255),
.B2(n_8),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_8),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_9),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_10),
.B(n_0),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_10),
.C(n_0),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_0),
.Y(n_263)
);


endmodule