module real_aes_2881_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
INVx1_ASAP7_75t_L g23 ( .A(n_0), .Y(n_23) );
NAND3xp33_ASAP7_75t_SL g10 ( .A(n_1), .B(n_11), .C(n_12), .Y(n_10) );
INVx3_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
INVx1_ASAP7_75t_L g25 ( .A(n_3), .Y(n_25) );
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
AND2x2_ASAP7_75t_L g26 ( .A(n_4), .B(n_18), .Y(n_26) );
INVx1_ASAP7_75t_L g18 ( .A(n_5), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g6 ( .A(n_7), .B(n_19), .Y(n_6) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_8), .Y(n_7) );
NAND2xp5_ASAP7_75t_SL g8 ( .A(n_9), .B(n_15), .Y(n_8) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
INVx2_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g15 ( .A(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_21), .B(n_26), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_22), .B(n_24), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
INVx2_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
endmodule