module fake_jpeg_4464_n_60 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_60);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_25;
wire n_56;
wire n_31;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;

INVx4_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_7),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_14),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_39),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_3),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

OAI32xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_41),
.A3(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_47)
);

AND2x4_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_4),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_23),
.A2(n_6),
.B1(n_11),
.B2(n_27),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_20),
.A2(n_22),
.B1(n_28),
.B2(n_24),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_21),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

AND2x6_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_41),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_41),
.B2(n_49),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_49),
.B1(n_42),
.B2(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_37),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_45),
.C(n_42),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_33),
.C(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

AOI322xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_54),
.A3(n_30),
.B1(n_22),
.B2(n_44),
.C1(n_39),
.C2(n_46),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_32),
.B1(n_31),
.B2(n_40),
.Y(n_60)
);


endmodule