module fake_ariane_416_n_777 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_777);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_777;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_74),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_45),
.Y(n_162)
);

BUFx4f_ASAP7_75t_SL g163 ( 
.A(n_3),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_68),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_21),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_86),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_75),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_60),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_43),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_25),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_14),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_22),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_36),
.B(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_55),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_8),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_8),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_99),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_23),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_63),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_70),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_65),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_11),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_57),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_2),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_84),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_2),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_9),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_146),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_30),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_52),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_59),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_127),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_40),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_61),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_117),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_123),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

AOI22x1_ASAP7_75t_SL g216 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_161),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_163),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_160),
.A2(n_0),
.B(n_1),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_4),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_174),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_164),
.A2(n_5),
.B(n_6),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_7),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_165),
.B(n_18),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_162),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_162),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g241 ( 
.A(n_167),
.B(n_19),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g243 ( 
.A1(n_168),
.A2(n_83),
.B(n_153),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_170),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_169),
.B(n_10),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_185),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_205),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

CKINVDCx6p67_ASAP7_75t_R g256 ( 
.A(n_175),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_240),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_175),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_193),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_182),
.Y(n_264)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_245),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_214),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_191),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_192),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_221),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_229),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_194),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_220),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_230),
.B(n_196),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_231),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_231),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_231),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_225),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_227),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_244),
.A2(n_213),
.B(n_202),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_247),
.Y(n_294)
);

BUFx6f_ASAP7_75t_SL g295 ( 
.A(n_253),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_206),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_218),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_228),
.Y(n_300)
);

AO21x2_ASAP7_75t_L g301 ( 
.A1(n_243),
.A2(n_207),
.B(n_210),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_246),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_249),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_224),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_269),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_249),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_298),
.B(n_234),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_264),
.A2(n_235),
.B1(n_232),
.B2(n_236),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_260),
.B(n_249),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_237),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_248),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_237),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_280),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_300),
.B(n_235),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_248),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_272),
.B(n_224),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_265),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_252),
.Y(n_327)
);

AND2x4_ASAP7_75t_SL g328 ( 
.A(n_265),
.B(n_222),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_239),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_262),
.B(n_225),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_L g334 ( 
.A(n_299),
.B(n_239),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_262),
.B(n_282),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_225),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_273),
.B(n_226),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_285),
.B(n_226),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_L g340 ( 
.A(n_287),
.B(n_241),
.C(n_182),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_288),
.B(n_222),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_289),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_292),
.B(n_296),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_303),
.B(n_163),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_281),
.B(n_247),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_297),
.B(n_205),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_251),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_305),
.B(n_247),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_217),
.Y(n_354)
);

BUFx6f_ASAP7_75t_SL g355 ( 
.A(n_284),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_259),
.B(n_166),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_301),
.A2(n_233),
.B1(n_223),
.B2(n_238),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_304),
.B(n_247),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_259),
.B(n_171),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_257),
.B(n_267),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_295),
.B(n_217),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_259),
.B(n_172),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_257),
.B(n_267),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_268),
.Y(n_365)
);

OR2x6_ASAP7_75t_L g366 ( 
.A(n_295),
.B(n_216),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_259),
.B(n_173),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_294),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_268),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_271),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_301),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_310),
.B(n_176),
.Y(n_372)
);

AO21x1_ASAP7_75t_L g373 ( 
.A1(n_340),
.A2(n_243),
.B(n_293),
.Y(n_373)
);

OAI321xp33_ASAP7_75t_L g374 ( 
.A1(n_317),
.A2(n_279),
.A3(n_277),
.B1(n_274),
.B2(n_271),
.C(n_294),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_327),
.B(n_259),
.Y(n_375)
);

O2A1O1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_307),
.A2(n_233),
.B(n_223),
.C(n_301),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_323),
.A2(n_319),
.B1(n_309),
.B2(n_338),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_314),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_371),
.A2(n_233),
.B(n_223),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_312),
.A2(n_313),
.B(n_314),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_313),
.B(n_177),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_189),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_330),
.B(n_12),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_315),
.B(n_195),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_357),
.A2(n_238),
.B(n_274),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_308),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_318),
.A2(n_279),
.B(n_277),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_321),
.B(n_197),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_316),
.A2(n_198),
.B1(n_208),
.B2(n_211),
.Y(n_392)
);

O2A1O1Ixp5_ASAP7_75t_L g393 ( 
.A1(n_339),
.A2(n_238),
.B(n_212),
.C(n_14),
.Y(n_393)
);

OAI21xp33_ASAP7_75t_L g394 ( 
.A1(n_325),
.A2(n_294),
.B(n_275),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_336),
.A2(n_217),
.B(n_275),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_344),
.A2(n_217),
.B(n_275),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_319),
.A2(n_275),
.B(n_294),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_238),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_306),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_352),
.A2(n_275),
.B(n_294),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_321),
.A2(n_87),
.B(n_152),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_324),
.B(n_12),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_324),
.B(n_13),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_306),
.Y(n_404)
);

AND2x2_ASAP7_75t_SL g405 ( 
.A(n_328),
.B(n_13),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_322),
.B(n_15),
.Y(n_407)
);

NOR3xp33_ASAP7_75t_L g408 ( 
.A(n_326),
.B(n_15),
.C(n_16),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_20),
.Y(n_409)
);

OAI321xp33_ASAP7_75t_L g410 ( 
.A1(n_341),
.A2(n_16),
.A3(n_17),
.B1(n_157),
.B2(n_26),
.C(n_27),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g411 ( 
.A(n_311),
.B(n_334),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_350),
.A2(n_90),
.B(n_24),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_325),
.B(n_17),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_350),
.A2(n_28),
.B(n_29),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_320),
.A2(n_31),
.B(n_32),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_354),
.A2(n_33),
.B(n_34),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_333),
.A2(n_360),
.B(n_356),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_357),
.A2(n_35),
.B(n_37),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_362),
.B(n_38),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_329),
.B(n_39),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_362),
.B(n_41),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g423 ( 
.A1(n_361),
.A2(n_42),
.B(n_44),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_360),
.A2(n_363),
.B(n_367),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_343),
.B(n_151),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_340),
.B(n_46),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_345),
.B(n_47),
.Y(n_427)
);

AOI21x1_ASAP7_75t_L g428 ( 
.A1(n_364),
.A2(n_48),
.B(n_49),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_346),
.B(n_50),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_355),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_347),
.B(n_149),
.Y(n_431)
);

O2A1O1Ixp5_ASAP7_75t_L g432 ( 
.A1(n_351),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_342),
.B(n_145),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_359),
.A2(n_56),
.B(n_58),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_349),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_368),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_358),
.B(n_370),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_365),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_355),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_358),
.A2(n_62),
.B(n_66),
.C(n_67),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_142),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_380),
.A2(n_353),
.B(n_366),
.Y(n_442)
);

AOI21x1_ASAP7_75t_L g443 ( 
.A1(n_398),
.A2(n_353),
.B(n_366),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_399),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_381),
.A2(n_419),
.B(n_417),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

AO31x2_ASAP7_75t_L g447 ( 
.A1(n_373),
.A2(n_69),
.A3(n_71),
.B(n_72),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_366),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_419),
.A2(n_73),
.B(n_76),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_388),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_377),
.A2(n_77),
.B(n_78),
.C(n_79),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_80),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_81),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_398),
.A2(n_82),
.B(n_88),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_402),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_372),
.B(n_93),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_391),
.A2(n_403),
.B(n_424),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_384),
.B(n_94),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_437),
.A2(n_95),
.B(n_96),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_385),
.B(n_97),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_405),
.B(n_98),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_379),
.A2(n_100),
.B(n_101),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_378),
.B(n_102),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_104),
.Y(n_465)
);

AOI21xp33_ASAP7_75t_L g466 ( 
.A1(n_426),
.A2(n_105),
.B(n_107),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_378),
.B(n_108),
.Y(n_467)
);

BUFx8_ASAP7_75t_L g468 ( 
.A(n_411),
.Y(n_468)
);

NOR2x1_ASAP7_75t_SL g469 ( 
.A(n_399),
.B(n_109),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_439),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_110),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_379),
.A2(n_112),
.B(n_113),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

AO21x1_ASAP7_75t_L g474 ( 
.A1(n_421),
.A2(n_431),
.B(n_420),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_409),
.B(n_114),
.Y(n_475)
);

AOI21x1_ASAP7_75t_L g476 ( 
.A1(n_397),
.A2(n_115),
.B(n_116),
.Y(n_476)
);

AOI21x1_ASAP7_75t_L g477 ( 
.A1(n_390),
.A2(n_120),
.B(n_121),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_389),
.A2(n_404),
.B(n_421),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_392),
.B(n_122),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_392),
.B(n_124),
.Y(n_480)
);

AOI21x1_ASAP7_75t_L g481 ( 
.A1(n_400),
.A2(n_425),
.B(n_433),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_387),
.A2(n_126),
.B(n_128),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_375),
.B(n_131),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_406),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_418),
.B(n_132),
.Y(n_485)
);

BUFx2_ASAP7_75t_SL g486 ( 
.A(n_427),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_387),
.A2(n_134),
.B(n_135),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_376),
.A2(n_136),
.B(n_137),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_438),
.B(n_141),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_438),
.B(n_138),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_401),
.A2(n_140),
.B(n_395),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_394),
.A2(n_407),
.B(n_396),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_408),
.B(n_407),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_429),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_441),
.B(n_414),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_423),
.A2(n_428),
.B(n_415),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_412),
.B(n_440),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_374),
.B(n_410),
.Y(n_498)
);

AOI21x1_ASAP7_75t_L g499 ( 
.A1(n_445),
.A2(n_434),
.B(n_416),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_450),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_446),
.Y(n_501)
);

OAI21x1_ASAP7_75t_SL g502 ( 
.A1(n_488),
.A2(n_432),
.B(n_393),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_462),
.B(n_493),
.Y(n_503)
);

OAI21x1_ASAP7_75t_SL g504 ( 
.A1(n_488),
.A2(n_442),
.B(n_480),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_444),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_496),
.A2(n_481),
.B(n_478),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_473),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_448),
.B(n_470),
.Y(n_509)
);

OAI21x1_ASAP7_75t_SL g510 ( 
.A1(n_479),
.A2(n_443),
.B(n_469),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_484),
.Y(n_511)
);

INVx6_ASAP7_75t_L g512 ( 
.A(n_444),
.Y(n_512)
);

AOI21x1_ASAP7_75t_L g513 ( 
.A1(n_492),
.A2(n_458),
.B(n_474),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_452),
.B(n_454),
.Y(n_514)
);

AOI22x1_ASAP7_75t_L g515 ( 
.A1(n_453),
.A2(n_497),
.B1(n_455),
.B2(n_460),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_471),
.Y(n_516)
);

CKINVDCx6p67_ASAP7_75t_R g517 ( 
.A(n_471),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_482),
.A2(n_487),
.B(n_472),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_452),
.B(n_444),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_468),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_473),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_485),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_473),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_477),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_475),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_495),
.A2(n_457),
.B(n_449),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_465),
.B(n_475),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_463),
.A2(n_491),
.B(n_467),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_459),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_489),
.A2(n_490),
.B(n_483),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_486),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_494),
.A2(n_464),
.B(n_456),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_451),
.A2(n_466),
.B(n_461),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_456),
.A2(n_447),
.B(n_466),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_447),
.Y(n_536)
);

AO21x2_ASAP7_75t_L g537 ( 
.A1(n_447),
.A2(n_492),
.B(n_488),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_488),
.B(n_298),
.C(n_264),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_496),
.A2(n_481),
.B(n_445),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_462),
.B(n_450),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_498),
.A2(n_256),
.B1(n_317),
.B2(n_341),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_450),
.B(n_471),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_453),
.B(n_461),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_450),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_496),
.A2(n_481),
.B(n_445),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_516),
.A2(n_503),
.B1(n_541),
.B2(n_540),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_542),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_501),
.Y(n_548)
);

NAND2x1_ASAP7_75t_L g549 ( 
.A(n_504),
.B(n_510),
.Y(n_549)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

CKINVDCx11_ASAP7_75t_R g551 ( 
.A(n_520),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_503),
.A2(n_538),
.B1(n_517),
.B2(n_540),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_517),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_518),
.A2(n_545),
.B(n_539),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_542),
.B(n_528),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_544),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_513),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_519),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_508),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_518),
.A2(n_545),
.B(n_539),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_508),
.Y(n_563)
);

INVxp33_ASAP7_75t_L g564 ( 
.A(n_509),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_507),
.A2(n_529),
.B(n_499),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_521),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_526),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g569 ( 
.A1(n_536),
.A2(n_535),
.B(n_524),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_522),
.A2(n_511),
.B1(n_528),
.B2(n_542),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_521),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_506),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_526),
.B(n_519),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_519),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_529),
.A2(n_527),
.B(n_531),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_523),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_530),
.B(n_512),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_532),
.A2(n_515),
.B1(n_535),
.B2(n_534),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_543),
.A2(n_532),
.B1(n_514),
.B2(n_537),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_514),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_512),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_533),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_505),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_566),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_548),
.B(n_512),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_578),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_578),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_559),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_581),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_581),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_572),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_555),
.B(n_537),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_549),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_547),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_555),
.B(n_512),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_553),
.B(n_506),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_557),
.B(n_543),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_557),
.B(n_533),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_569),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_556),
.B(n_520),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_553),
.Y(n_602)
);

NOR2x1_ASAP7_75t_L g603 ( 
.A(n_568),
.B(n_534),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_569),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_560),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_558),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_569),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_546),
.A2(n_534),
.B1(n_502),
.B2(n_531),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_558),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_583),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_553),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_556),
.B(n_574),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_574),
.Y(n_613)
);

AOI222xp33_ASAP7_75t_L g614 ( 
.A1(n_570),
.A2(n_551),
.B1(n_573),
.B2(n_550),
.C1(n_580),
.C2(n_575),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_583),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_560),
.B(n_567),
.Y(n_616)
);

NAND2x1p5_ASAP7_75t_L g617 ( 
.A(n_568),
.B(n_552),
.Y(n_617)
);

AOI221xp5_ASAP7_75t_L g618 ( 
.A1(n_552),
.A2(n_579),
.B1(n_567),
.B2(n_571),
.C(n_563),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_559),
.B(n_575),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_559),
.B(n_575),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_562),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_577),
.Y(n_622)
);

AOI211xp5_ASAP7_75t_L g623 ( 
.A1(n_568),
.A2(n_582),
.B(n_575),
.C(n_576),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_575),
.B(n_568),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_592),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_590),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_593),
.B(n_562),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_593),
.B(n_562),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_591),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_602),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_599),
.B(n_561),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_610),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_599),
.B(n_561),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_592),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_610),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_612),
.B(n_582),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_624),
.B(n_582),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_612),
.B(n_547),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_587),
.B(n_554),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_594),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_588),
.B(n_554),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_602),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_615),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_615),
.Y(n_644)
);

NOR2xp67_ASAP7_75t_L g645 ( 
.A(n_584),
.B(n_573),
.Y(n_645)
);

OAI221xp5_ASAP7_75t_SL g646 ( 
.A1(n_618),
.A2(n_547),
.B1(n_549),
.B2(n_576),
.C(n_565),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_609),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_606),
.B(n_565),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_598),
.B(n_613),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_601),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_609),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_598),
.Y(n_652)
);

BUFx4f_ASAP7_75t_L g653 ( 
.A(n_617),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_613),
.B(n_606),
.Y(n_654)
);

NOR2x1_ASAP7_75t_SL g655 ( 
.A(n_602),
.B(n_611),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_608),
.A2(n_617),
.B1(n_586),
.B2(n_611),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_585),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_585),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_596),
.B(n_616),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_629),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_626),
.B(n_596),
.Y(n_661)
);

AND2x4_ASAP7_75t_SL g662 ( 
.A(n_642),
.B(n_624),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_625),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_627),
.B(n_628),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_652),
.B(n_605),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_632),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_655),
.B(n_630),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_654),
.B(n_607),
.Y(n_668)
);

NAND2x1p5_ASAP7_75t_L g669 ( 
.A(n_653),
.B(n_611),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_627),
.B(n_621),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_628),
.B(n_621),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_649),
.B(n_616),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_655),
.B(n_594),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_631),
.B(n_603),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_630),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_631),
.B(n_603),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_649),
.B(n_617),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_646),
.B(n_597),
.C(n_623),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_633),
.B(n_623),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_625),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_634),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_633),
.B(n_600),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_632),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_654),
.B(n_600),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_639),
.B(n_604),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_660),
.B(n_650),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_664),
.B(n_659),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_666),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_678),
.B(n_642),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_679),
.A2(n_614),
.B1(n_597),
.B2(n_656),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_664),
.B(n_639),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_662),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_672),
.B(n_644),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_683),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_661),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_665),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_679),
.B(n_641),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_668),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_682),
.B(n_641),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_663),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_668),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_695),
.B(n_682),
.Y(n_702)
);

AOI21x1_ASAP7_75t_L g703 ( 
.A1(n_689),
.A2(n_645),
.B(n_673),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_688),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_690),
.A2(n_614),
.B1(n_676),
.B2(n_674),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_696),
.B(n_674),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_694),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_689),
.A2(n_676),
.B1(n_677),
.B2(n_653),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_692),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_693),
.B(n_685),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_697),
.B(n_685),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_709),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_704),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_SL g714 ( 
.A1(n_705),
.A2(n_701),
.B1(n_698),
.B2(n_687),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_707),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_708),
.A2(n_667),
.B(n_673),
.Y(n_716)
);

AOI222xp33_ASAP7_75t_L g717 ( 
.A1(n_706),
.A2(n_686),
.B1(n_699),
.B2(n_671),
.C1(n_670),
.C2(n_647),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_714),
.A2(n_717),
.B1(n_716),
.B2(n_712),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_713),
.B(n_709),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_715),
.Y(n_720)
);

OAI21xp33_ASAP7_75t_SL g721 ( 
.A1(n_712),
.A2(n_711),
.B(n_691),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_713),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_712),
.A2(n_703),
.B1(n_710),
.B2(n_702),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_719),
.B(n_642),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_722),
.B(n_686),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_720),
.B(n_699),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_723),
.Y(n_727)
);

NOR4xp75_ASAP7_75t_L g728 ( 
.A(n_725),
.B(n_721),
.C(n_718),
.D(n_675),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_726),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_729),
.Y(n_730)
);

NOR3xp33_ASAP7_75t_L g731 ( 
.A(n_728),
.B(n_727),
.C(n_636),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_728),
.B(n_667),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_730),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_732),
.B(n_724),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_731),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_730),
.Y(n_736)
);

NOR2x1_ASAP7_75t_L g737 ( 
.A(n_730),
.B(n_667),
.Y(n_737)
);

XOR2x1_ASAP7_75t_L g738 ( 
.A(n_730),
.B(n_669),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_736),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_733),
.B(n_675),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_735),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_738),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_737),
.Y(n_743)
);

XOR2xp5_ASAP7_75t_L g744 ( 
.A(n_734),
.B(n_637),
.Y(n_744)
);

XOR2xp5_ASAP7_75t_L g745 ( 
.A(n_744),
.B(n_637),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_743),
.A2(n_673),
.B1(n_669),
.B2(n_635),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_SL g747 ( 
.A1(n_743),
.A2(n_662),
.B1(n_653),
.B2(n_637),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_741),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_739),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_740),
.Y(n_750)
);

OAI331xp33_ASAP7_75t_L g751 ( 
.A1(n_748),
.A2(n_742),
.A3(n_644),
.B1(n_643),
.B2(n_635),
.B3(n_638),
.C1(n_619),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_749),
.Y(n_752)
);

AOI21xp33_ASAP7_75t_L g753 ( 
.A1(n_750),
.A2(n_700),
.B(n_657),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_745),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_746),
.Y(n_755)
);

OAI22x1_ASAP7_75t_L g756 ( 
.A1(n_747),
.A2(n_640),
.B1(n_594),
.B2(n_589),
.Y(n_756)
);

AOI21x1_ASAP7_75t_L g757 ( 
.A1(n_748),
.A2(n_643),
.B(n_671),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_749),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_749),
.A2(n_648),
.B(n_640),
.Y(n_759)
);

AOI311xp33_ASAP7_75t_L g760 ( 
.A1(n_752),
.A2(n_658),
.A3(n_657),
.B(n_648),
.C(n_594),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_754),
.A2(n_700),
.B1(n_658),
.B2(n_651),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_758),
.Y(n_762)
);

AOI21xp33_ASAP7_75t_L g763 ( 
.A1(n_755),
.A2(n_651),
.B(n_647),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_759),
.Y(n_764)
);

AOI21xp33_ASAP7_75t_L g765 ( 
.A1(n_756),
.A2(n_684),
.B(n_622),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_757),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_751),
.A2(n_640),
.B(n_595),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_SL g768 ( 
.A1(n_762),
.A2(n_753),
.B(n_670),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_764),
.B(n_766),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_763),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_761),
.Y(n_771)
);

AO21x2_ASAP7_75t_L g772 ( 
.A1(n_767),
.A2(n_620),
.B(n_684),
.Y(n_772)
);

AO21x2_ASAP7_75t_L g773 ( 
.A1(n_769),
.A2(n_765),
.B(n_760),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_L g774 ( 
.A(n_770),
.B(n_589),
.Y(n_774)
);

INVx3_ASAP7_75t_L g775 ( 
.A(n_773),
.Y(n_775)
);

AOI221xp5_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_771),
.B1(n_774),
.B2(n_768),
.C(n_772),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_776),
.A2(n_622),
.B1(n_681),
.B2(n_680),
.Y(n_777)
);


endmodule