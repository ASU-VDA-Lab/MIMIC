module fake_netlist_6_4316_n_464 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_464);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_464;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_235;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_156;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_397;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_460;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_456;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_321;
wire n_331;
wire n_227;
wire n_406;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_164;
wire n_292;
wire n_307;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_319;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_459;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_17),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_58),
.B(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_107),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_44),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_43),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_55),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_7),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_40),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_62),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_25),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_10),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_86),
.Y(n_182)
);

INVxp33_ASAP7_75t_SL g183 ( 
.A(n_87),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_95),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_56),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_47),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_134),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_49),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_70),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_38),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_50),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_27),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_12),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_63),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_41),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_33),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_151),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_53),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_59),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_75),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_74),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_72),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_84),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_4),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_42),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_135),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_23),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_0),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_16),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_69),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_113),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_64),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_21),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_34),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_81),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_20),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_98),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_48),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_54),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_118),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_28),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_90),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_14),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_139),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_82),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_121),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_24),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_140),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_37),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_68),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_89),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_67),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_35),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_102),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_138),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_99),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_19),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_120),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_93),
.Y(n_254)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_3),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_155),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_29),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_126),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_127),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_79),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_9),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_83),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_124),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g264 ( 
.A(n_52),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_71),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_18),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_123),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_92),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_88),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_85),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_105),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_66),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_60),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_122),
.B(n_2),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_13),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_61),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_152),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_142),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_156),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_229),
.B(n_5),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_157),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_159),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_169),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_161),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_176),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_R g286 ( 
.A(n_174),
.B(n_6),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_187),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_162),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_168),
.B(n_8),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_164),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_165),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_188),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_193),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_177),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_189),
.Y(n_295)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_255),
.C(n_238),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_166),
.B(n_15),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_194),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_167),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_R g300 ( 
.A(n_182),
.B(n_22),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_202),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_205),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_222),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_171),
.Y(n_304)
);

AND3x2_ASAP7_75t_L g305 ( 
.A(n_179),
.B(n_26),
.C(n_31),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_223),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_173),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_178),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_224),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_232),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_180),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_240),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_243),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_251),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_192),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_263),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_266),
.Y(n_318)
);

NAND2xp33_ASAP7_75t_R g319 ( 
.A(n_183),
.B(n_32),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_195),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_220),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_181),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_198),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_212),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_184),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_R g326 ( 
.A(n_226),
.B(n_265),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_R g327 ( 
.A(n_268),
.B(n_36),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_237),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_185),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_R g330 ( 
.A(n_190),
.B(n_39),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_191),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_196),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_197),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_170),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_283),
.Y(n_336)
);

OAI221xp5_ASAP7_75t_L g337 ( 
.A1(n_296),
.A2(n_262),
.B1(n_172),
.B2(n_257),
.C(n_216),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_326),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_287),
.B(n_292),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_289),
.B(n_264),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_331),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_332),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_298),
.B(n_215),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_320),
.A2(n_250),
.B1(n_252),
.B2(n_276),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_209),
.Y(n_350)
);

AO22x2_ASAP7_75t_L g351 ( 
.A1(n_288),
.A2(n_210),
.B1(n_277),
.B2(n_275),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_290),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_233),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_175),
.Y(n_355)
);

OR2x2_ASAP7_75t_SL g356 ( 
.A(n_295),
.B(n_199),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

BUFx6f_ASAP7_75t_SL g358 ( 
.A(n_313),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_309),
.B(n_186),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

BUFx8_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_312),
.B(n_269),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_314),
.B(n_273),
.Y(n_366)
);

NAND2x1p5_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_160),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_315),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_158),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_163),
.Y(n_370)
);

BUFx8_ASAP7_75t_L g371 ( 
.A(n_329),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_342),
.B(n_321),
.Y(n_372)
);

NAND2x1p5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_200),
.Y(n_373)
);

BUFx12f_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_SL g375 ( 
.A1(n_337),
.A2(n_304),
.B(n_297),
.C(n_241),
.Y(n_375)
);

O2A1O1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_347),
.A2(n_299),
.B(n_304),
.C(n_242),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_356),
.A2(n_328),
.B1(n_324),
.B2(n_323),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_338),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_350),
.A2(n_259),
.B(n_239),
.Y(n_379)
);

NAND3xp33_ASAP7_75t_SL g380 ( 
.A(n_340),
.B(n_300),
.C(n_286),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_346),
.B(n_313),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_341),
.A2(n_335),
.B1(n_348),
.B2(n_359),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_327),
.Y(n_384)
);

INVx3_ASAP7_75t_SL g385 ( 
.A(n_369),
.Y(n_385)
);

O2A1O1Ixp33_ASAP7_75t_SL g386 ( 
.A1(n_354),
.A2(n_213),
.B(n_219),
.C(n_218),
.Y(n_386)
);

O2A1O1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_349),
.A2(n_211),
.B(n_214),
.C(n_278),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_364),
.A2(n_366),
.B(n_370),
.Y(n_388)
);

O2A1O1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_362),
.A2(n_207),
.B(n_208),
.C(n_272),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_358),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_294),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_357),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_343),
.B(n_204),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_367),
.A2(n_316),
.B1(n_246),
.B2(n_206),
.Y(n_394)
);

AOI22x1_ASAP7_75t_L g395 ( 
.A1(n_351),
.A2(n_201),
.B1(n_203),
.B2(n_271),
.Y(n_395)
);

BUFx12f_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_352),
.Y(n_397)
);

AO21x2_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_330),
.B(n_253),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_379),
.A2(n_365),
.B(n_360),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_393),
.A2(n_353),
.B(n_217),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_374),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_383),
.A2(n_247),
.B(n_225),
.Y(n_403)
);

AOI221x1_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_248),
.B1(n_227),
.B2(n_228),
.C(n_230),
.Y(n_404)
);

OAI21x1_ASAP7_75t_L g405 ( 
.A1(n_395),
.A2(n_254),
.B(n_231),
.Y(n_405)
);

OA21x2_ASAP7_75t_L g406 ( 
.A1(n_397),
.A2(n_344),
.B(n_334),
.Y(n_406)
);

AO21x2_ASAP7_75t_L g407 ( 
.A1(n_372),
.A2(n_249),
.B(n_234),
.Y(n_407)
);

AO21x2_ASAP7_75t_L g408 ( 
.A1(n_375),
.A2(n_256),
.B(n_235),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

BUFx12f_ASAP7_75t_L g411 ( 
.A(n_396),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_392),
.B(n_260),
.Y(n_412)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

AO21x2_ASAP7_75t_L g414 ( 
.A1(n_381),
.A2(n_258),
.B(n_236),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_261),
.B1(n_244),
.B2(n_245),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_377),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_402),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_408),
.A2(n_415),
.B1(n_399),
.B2(n_406),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_410),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_416),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_407),
.B(n_414),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_401),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_412),
.Y(n_424)
);

NAND2x1_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_267),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_373),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_411),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_376),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_413),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_390),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_429),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

BUFx5_ASAP7_75t_L g433 ( 
.A(n_430),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_426),
.A2(n_371),
.B1(n_221),
.B2(n_319),
.Y(n_434)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_420),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_424),
.A2(n_386),
.B(n_387),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_428),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_417),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_432),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_423),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_423),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_438),
.A2(n_434),
.B1(n_428),
.B2(n_437),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_435),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_440),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_439),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_444),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_446),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_422),
.Y(n_449)
);

NAND4xp25_ASAP7_75t_L g450 ( 
.A(n_447),
.B(n_389),
.C(n_427),
.D(n_419),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_445),
.Y(n_451)
);

OAI21xp33_ASAP7_75t_SL g452 ( 
.A1(n_450),
.A2(n_305),
.B(n_46),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_448),
.B(n_45),
.Y(n_453)
);

AOI221x1_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_451),
.B1(n_449),
.B2(n_425),
.C(n_80),
.Y(n_454)
);

AND4x2_ASAP7_75t_L g455 ( 
.A(n_452),
.B(n_51),
.C(n_57),
.D(n_78),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_454),
.B(n_91),
.Y(n_456)
);

AOI211xp5_ASAP7_75t_L g457 ( 
.A1(n_455),
.A2(n_94),
.B(n_96),
.C(n_97),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_456),
.Y(n_458)
);

INVx5_ASAP7_75t_L g459 ( 
.A(n_457),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_458),
.B(n_100),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_460),
.Y(n_461)
);

OAI221xp5_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_459),
.B1(n_103),
.B2(n_104),
.C(n_106),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_462),
.A2(n_150),
.B1(n_111),
.B2(n_112),
.Y(n_463)
);

AOI221xp5_ASAP7_75t_L g464 ( 
.A1(n_463),
.A2(n_101),
.B1(n_117),
.B2(n_119),
.C(n_125),
.Y(n_464)
);


endmodule