module fake_jpeg_28613_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_79),
.B(n_69),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_82),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_91),
.B(n_94),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_72),
.Y(n_96)
);

AND2x4_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_58),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_50),
.B1(n_67),
.B2(n_66),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_53),
.B(n_89),
.C(n_85),
.Y(n_121)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_107),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_52),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_58),
.B1(n_70),
.B2(n_61),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_112),
.B1(n_99),
.B2(n_111),
.Y(n_125)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_53),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_112),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_54),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_70),
.B1(n_68),
.B2(n_56),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_92),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_121),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_8),
.Y(n_137)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_24),
.A3(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_7),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_3),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_4),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_48),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_5),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_138),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_8),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_9),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_19),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_151),
.B(n_32),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_41),
.Y(n_146)
);

XNOR2x2_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_149),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_115),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_148),
.B(n_119),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_22),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_121),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_30),
.C(n_31),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_153),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_119),
.B1(n_127),
.B2(n_38),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_146),
.C(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_155),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_166),
.B1(n_161),
.B2(n_143),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_144),
.B(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_163),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_154),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_158),
.B(n_162),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_40),
.B(n_153),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_136),
.Y(n_173)
);


endmodule