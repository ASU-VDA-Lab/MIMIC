module fake_jpeg_23019_n_40 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_40);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_16),
.Y(n_22)
);

OR2x2_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_0),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_26),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_30),
.B1(n_9),
.B2(n_10),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_32),
.B1(n_13),
.B2(n_14),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_34),
.B(n_35),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_27),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

BUFx24_ASAP7_75t_SL g40 ( 
.A(n_39),
.Y(n_40)
);


endmodule