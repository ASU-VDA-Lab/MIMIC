module fake_netlist_1_1187_n_24 (n_1, n_2, n_4, n_3, n_5, n_0, n_24);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
INVx2_ASAP7_75t_SL g6 ( .A(n_2), .Y(n_6) );
INVx2_ASAP7_75t_SL g7 ( .A(n_0), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_3), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_2), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
A2O1A1Ixp33_ASAP7_75t_L g11 ( .A1(n_6), .A2(n_1), .B(n_3), .C(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_6), .B(n_1), .Y(n_13) );
OAI21x1_ASAP7_75t_L g14 ( .A1(n_9), .A2(n_4), .B(n_5), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_13), .B(n_7), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
NOR2x1_ASAP7_75t_L g17 ( .A(n_15), .B(n_13), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_15), .B(n_14), .Y(n_18) );
AOI221xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_11), .B1(n_12), .B2(n_8), .C(n_10), .Y(n_19) );
AOI22xp5_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_16), .B1(n_7), .B2(n_8), .Y(n_20) );
NAND4xp75_ASAP7_75t_L g21 ( .A(n_19), .B(n_10), .C(n_12), .D(n_16), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_20), .B(n_14), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_5), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
endmodule