module real_jpeg_14622_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_312, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_312;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_50),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_2),
.A2(n_50),
.B1(n_58),
.B2(n_62),
.Y(n_258)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_4),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_4),
.A2(n_58),
.B1(n_62),
.B2(n_165),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_165),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_165),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_7),
.A2(n_58),
.B1(n_62),
.B2(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_8),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_8),
.A2(n_37),
.B1(n_58),
.B2(n_62),
.Y(n_224)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_10),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_10),
.A2(n_29),
.B1(n_58),
.B2(n_62),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_10),
.A2(n_29),
.B1(n_45),
.B2(n_46),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_11),
.B(n_33),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_12),
.A2(n_53),
.B1(n_58),
.B2(n_62),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_13),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_13),
.A2(n_58),
.B1(n_62),
.B2(n_96),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_96),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_14),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_58),
.B1(n_62),
.B2(n_136),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_136),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_136),
.Y(n_244)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_16),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_16),
.B(n_58),
.C(n_61),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_16),
.B(n_44),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_16),
.A2(n_127),
.B(n_169),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_16),
.A2(n_32),
.B(n_43),
.C(n_196),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_153),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_16),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_16),
.B(n_25),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_110),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_20),
.B(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_70),
.C(n_78),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_70),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_38),
.B2(n_69),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_22),
.A2(n_23),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_23),
.B(n_39),
.C(n_55),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_24),
.A2(n_31),
.B(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_26),
.A2(n_30),
.B(n_153),
.C(n_240),
.Y(n_239)
);

AOI32xp33_ASAP7_75t_L g253 ( 
.A1(n_26),
.A2(n_32),
.A3(n_34),
.B1(n_241),
.B2(n_254),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_30),
.A2(n_135),
.B(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_30),
.A2(n_31),
.B1(n_135),
.B2(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_31),
.B(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_31),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_31),
.A2(n_92),
.B(n_268),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_54),
.B1(n_55),
.B2(n_68),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_48),
.B2(n_51),
.Y(n_39)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_40),
.B(n_203),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

AO22x1_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_42),
.A2(n_45),
.B(n_153),
.Y(n_196)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_44),
.B(n_203),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_64)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_46),
.B(n_157),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_52),
.A2(n_72),
.B1(n_74),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_55),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B(n_65),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_63),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_56),
.A2(n_63),
.B1(n_89),
.B2(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_56),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_56),
.A2(n_63),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_56),
.A2(n_63),
.B1(n_131),
.B2(n_247),
.Y(n_273)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_57),
.A2(n_164),
.B(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_57),
.B(n_153),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_57),
.A2(n_166),
.B(n_246),
.Y(n_245)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_62),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_63),
.B(n_155),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_71),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_72),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_72),
.A2(n_74),
.B1(n_216),
.B2(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_72),
.A2(n_202),
.B(n_244),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_74),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_74),
.A2(n_133),
.B(n_217),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_76),
.A2(n_152),
.B(n_154),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_76),
.A2(n_154),
.B(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B(n_91),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_80),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_82),
.B1(n_91),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_83),
.A2(n_84),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_83),
.B(n_170),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_83),
.A2(n_84),
.B1(n_126),
.B2(n_258),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_84),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_84),
.B(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_139),
.B(n_310),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_112),
.B(n_114),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_121),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_120),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_121),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.C(n_134),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_122),
.A2(n_123),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_124),
.A2(n_129),
.B1(n_130),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_124),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_127),
.A2(n_128),
.B1(n_198),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_127),
.A2(n_128),
.B1(n_224),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_128),
.A2(n_175),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_153),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_128),
.A2(n_183),
.B(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_132),
.B(n_134),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_138),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_304),
.B(n_309),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_292),
.B(n_303),
.Y(n_142)
);

OAI321xp33_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_260),
.A3(n_285),
.B1(n_290),
.B2(n_291),
.C(n_312),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_233),
.B(n_259),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_210),
.B(n_232),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_191),
.B(n_209),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_171),
.B(n_190),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_158),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_149),
.B(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_156),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_151),
.B1(n_156),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_167),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_163),
.C(n_167),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_168),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_179),
.B(n_189),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_177),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_184),
.B(n_188),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_193),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_204),
.C(n_208),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_197),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_199)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_225),
.B2(n_226),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_228),
.C(n_230),
.Y(n_234)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_219),
.C(n_223),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_234),
.B(n_235),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_249),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_236),
.B(n_250),
.C(n_251),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_242),
.B2(n_248),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_243),
.C(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_256),
.Y(n_270)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_275),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_271),
.C(n_274),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_263),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_270),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_269),
.C(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_274),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_284),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_279),
.C(n_284),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.C(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_302),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_302),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_297),
.C(n_298),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);


endmodule