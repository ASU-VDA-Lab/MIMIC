module real_jpeg_1024_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_4),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_60),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_60),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_5),
.A2(n_39),
.B1(n_40),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_68),
.Y(n_120)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_11),
.A2(n_22),
.B1(n_23),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_12),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_12),
.A2(n_39),
.B(n_44),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_12),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_12),
.B(n_25),
.C(n_28),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_12),
.B(n_51),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_12),
.B(n_103),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_91),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_89),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_81),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_17),
.B(n_81),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_56),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_31),
.B(n_34),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_20),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_20),
.A2(n_86),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_20),
.A2(n_102),
.B1(n_103),
.B2(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_46),
.Y(n_45)
);

OA22x2_ASAP7_75t_SL g64 ( 
.A1(n_22),
.A2(n_23),
.B1(n_41),
.B2(n_46),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI32xp33_ASAP7_75t_L g38 ( 
.A1(n_23),
.A2(n_39),
.A3(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_23),
.B(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_25),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_27),
.A2(n_32),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_28),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_28),
.B(n_115),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_47),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_38),
.B(n_47),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_46),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_40),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_52),
.B(n_53),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_48),
.A2(n_50),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_49),
.B(n_54),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_49),
.A2(n_51),
.B1(n_100),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_49),
.A2(n_51),
.B1(n_117),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_50),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_69),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_62),
.B1(n_64),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.C(n_87),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_87),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_130),
.B(n_135),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_111),
.B(n_129),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_104),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_104),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_101),
.C(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_123),
.B(n_128),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_118),
.B(n_122),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_121),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_127),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_133),
.Y(n_135)
);


endmodule