module fake_jpeg_2993_n_399 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_399);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_399;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_44),
.Y(n_127)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_46),
.Y(n_129)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_27),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g131 ( 
.A(n_48),
.Y(n_131)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_8),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_54),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_64),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_23),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_68),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_15),
.A2(n_9),
.B(n_13),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_80),
.Y(n_114)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_9),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_26),
.B(n_9),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_82),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_29),
.B(n_14),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_33),
.Y(n_95)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_86),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_85),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_22),
.B1(n_28),
.B2(n_39),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_88),
.A2(n_90),
.B1(n_94),
.B2(n_99),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_15),
.B1(n_27),
.B2(n_35),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_26),
.B1(n_28),
.B2(n_39),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_95),
.B(n_12),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_107),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_29),
.B1(n_31),
.B2(n_38),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_44),
.B(n_43),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_105),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_31),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_38),
.C(n_41),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_74),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_17),
.B1(n_41),
.B2(n_37),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_112),
.B1(n_74),
.B2(n_18),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_49),
.A2(n_18),
.B1(n_43),
.B2(n_36),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_18),
.B1(n_48),
.B2(n_79),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_45),
.A2(n_34),
.B1(n_30),
.B2(n_24),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_54),
.B(n_30),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_24),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_63),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_59),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_137),
.B(n_145),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_138),
.B(n_181),
.Y(n_225)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_139),
.Y(n_211)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_140),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_141),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_143),
.Y(n_192)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_146),
.A2(n_149),
.B1(n_151),
.B2(n_154),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_21),
.B(n_82),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_161),
.Y(n_190)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_21),
.B1(n_71),
.B2(n_46),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_107),
.A2(n_84),
.B1(n_82),
.B2(n_73),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_170),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_80),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_153),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_102),
.A2(n_73),
.B1(n_20),
.B2(n_65),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

MAJx3_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_62),
.C(n_2),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_159),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_168),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_59),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_160),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_11),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_3),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_119),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_125),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_171),
.A2(n_91),
.B1(n_106),
.B2(n_87),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_0),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_99),
.Y(n_205)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_96),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_180),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_177),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_183),
.Y(n_207)
);

INVx6_ASAP7_75t_SL g179 ( 
.A(n_116),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_179),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_118),
.Y(n_181)
);

AO22x2_ASAP7_75t_SL g182 ( 
.A1(n_98),
.A2(n_100),
.B1(n_124),
.B2(n_121),
.Y(n_182)
);

AO22x2_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_102),
.B1(n_121),
.B2(n_124),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_93),
.B(n_12),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_106),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_110),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_217),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_128),
.B(n_122),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_194),
.A2(n_201),
.B(n_168),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_157),
.A2(n_129),
.B(n_87),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_157),
.A2(n_129),
.B1(n_89),
.B2(n_91),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_159),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_116),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_150),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_145),
.B(n_100),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_98),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_148),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_142),
.B(n_92),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_172),
.C(n_159),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_234),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_143),
.C(n_180),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_215),
.C(n_192),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_231),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_237),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_167),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_236),
.Y(n_277)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_153),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_189),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_242),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_153),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_245),
.Y(n_282)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_139),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_190),
.B(n_173),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_179),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_198),
.A2(n_165),
.B1(n_182),
.B2(n_177),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_206),
.B1(n_194),
.B2(n_200),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_198),
.A2(n_182),
.B1(n_130),
.B2(n_155),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_249),
.A2(n_252),
.B1(n_203),
.B2(n_210),
.Y(n_286)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_198),
.A2(n_130),
.B1(n_144),
.B2(n_140),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_160),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_253),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_217),
.B(n_141),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_254),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_4),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_257),
.B(n_209),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_196),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_213),
.B(n_136),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_259),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_136),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_260),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_222),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_199),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_262),
.A2(n_266),
.B1(n_289),
.B2(n_249),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_215),
.B1(n_187),
.B2(n_204),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_274),
.C(n_275),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_239),
.A2(n_215),
.B(n_192),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_268),
.A2(n_228),
.B(n_245),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_219),
.C(n_199),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_204),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_234),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_281),
.B(n_247),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_227),
.B(n_216),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_285),
.C(n_231),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_226),
.B(n_216),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_246),
.B1(n_236),
.B2(n_230),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_228),
.A2(n_216),
.B1(n_185),
.B2(n_224),
.Y(n_289)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_298),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_248),
.B1(n_246),
.B2(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_251),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_299),
.A2(n_307),
.B(n_303),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_300),
.B(n_314),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_303),
.Y(n_319)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_251),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_287),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_304),
.B(n_305),
.Y(n_337)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_306),
.Y(n_334)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_313),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_SL g330 ( 
.A(n_309),
.B(n_312),
.C(n_279),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_263),
.A2(n_246),
.B1(n_228),
.B2(n_255),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_311),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_283),
.B(n_232),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_281),
.B(n_279),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_234),
.C(n_257),
.Y(n_314)
);

BUFx12_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_258),
.Y(n_338)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_269),
.B(n_284),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_268),
.C(n_267),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_331),
.C(n_332),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_316),
.A2(n_277),
.B1(n_282),
.B2(n_262),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_326),
.A2(n_271),
.B1(n_185),
.B2(n_241),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_300),
.B(n_265),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_327),
.B(n_335),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_301),
.A2(n_277),
.B1(n_289),
.B2(n_285),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_328),
.A2(n_329),
.B1(n_296),
.B2(n_254),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_338),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_274),
.C(n_275),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_294),
.B(n_276),
.C(n_266),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_333),
.A2(n_299),
.B(n_297),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_314),
.B(n_252),
.Y(n_335)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_337),
.B(n_313),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_342),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_334),
.B(n_302),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_343),
.A2(n_350),
.B(n_354),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_317),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_348),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_330),
.B(n_240),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_346),
.B(n_323),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_296),
.C(n_235),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_349),
.C(n_320),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_327),
.C(n_320),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_333),
.A2(n_296),
.B(n_255),
.Y(n_350)
);

A2O1A1O1Ixp25_ASAP7_75t_L g351 ( 
.A1(n_318),
.A2(n_250),
.B(n_243),
.C(n_308),
.D(n_291),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_351),
.A2(n_322),
.B(n_338),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_352),
.A2(n_325),
.B1(n_347),
.B2(n_323),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_322),
.A2(n_209),
.B(n_315),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_355),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_356),
.A2(n_354),
.B(n_351),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_203),
.C(n_186),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_335),
.C(n_328),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_359),
.B(n_364),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_350),
.A2(n_326),
.B1(n_318),
.B2(n_319),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_363),
.A2(n_368),
.B1(n_352),
.B2(n_353),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_325),
.C(n_321),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_353),
.B(n_329),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_365),
.Y(n_373)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_366),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_364),
.A2(n_344),
.B(n_343),
.Y(n_369)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_369),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_362),
.B(n_340),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_370),
.B(n_376),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_372),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_374),
.A2(n_357),
.B(n_367),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_361),
.B(n_349),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_357),
.A2(n_315),
.B(n_211),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_377),
.B(n_378),
.C(n_358),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_379),
.A2(n_383),
.B(n_373),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_380),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_359),
.C(n_360),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_382),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_224),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_372),
.B(n_365),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_388),
.A2(n_390),
.B1(n_391),
.B2(n_220),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_386),
.A2(n_373),
.B(n_363),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_186),
.B(n_197),
.Y(n_391)
);

AOI322xp5_ASAP7_75t_L g392 ( 
.A1(n_387),
.A2(n_383),
.A3(n_385),
.B1(n_197),
.B2(n_220),
.C1(n_164),
.C2(n_62),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_392),
.A2(n_393),
.B1(n_394),
.B2(n_220),
.Y(n_395)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_389),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_395),
.B(n_396),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_393),
.A2(n_13),
.B(n_5),
.Y(n_396)
);

BUFx24_ASAP7_75t_SL g398 ( 
.A(n_397),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_398),
.B(n_13),
.Y(n_399)
);


endmodule