module real_jpeg_3877_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_1),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_1),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_1),
.B(n_70),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_1),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_1),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_1),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_1),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_2),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_2),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_2),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_2),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_2),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_2),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_2),
.B(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_3),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_3),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_3),
.B(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_3),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_3),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_3),
.B(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_4),
.Y(n_171)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_4),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_5),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_5),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_5),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_5),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_5),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_5),
.B(n_368),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_5),
.B(n_409),
.Y(n_408)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_7),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_7),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_7),
.B(n_14),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_10),
.B(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_10),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_10),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_10),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_10),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_10),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_10),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_10),
.B(n_411),
.Y(n_410)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_11),
.Y(n_111)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_11),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_12),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_12),
.B(n_152),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_12),
.B(n_65),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_12),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_12),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_12),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_12),
.B(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_13),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_13),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_14),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_14),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_14),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_14),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_15),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_15),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_15),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_15),
.B(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_463),
.Y(n_16)
);

OAI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_218),
.B(n_460),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_182),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_SL g460 ( 
.A1(n_19),
.A2(n_461),
.B(n_462),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_138),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_20),
.B(n_138),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_99),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_21),
.B(n_100),
.C(n_115),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_68),
.C(n_80),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_22),
.B(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_48),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_23),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_33),
.B2(n_37),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_26),
.B(n_32),
.C(n_37),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_28),
.A2(n_32),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_28),
.B(n_205),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_28),
.A2(n_32),
.B1(n_204),
.B2(n_205),
.Y(n_427)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_29),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_30),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_39),
.C(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_33),
.A2(n_37),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_33),
.B(n_270),
.C(n_272),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_33),
.A2(n_37),
.B1(n_272),
.B2(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_35),
.Y(n_391)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_35),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_37),
.B(n_103),
.C(n_109),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_38),
.B(n_48),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_39),
.A2(n_119),
.B1(n_120),
.B2(n_127),
.Y(n_118)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_39),
.A2(n_44),
.B1(n_127),
.B2(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_43),
.Y(n_153)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_44),
.Y(n_149)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_47),
.Y(n_211)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_47),
.Y(n_365)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_47),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_55),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_55),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_56),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_61),
.C(n_64),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_56),
.B(n_196),
.Y(n_226)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_60),
.Y(n_271)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_60),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_62),
.B(n_195),
.C(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_63),
.A2(n_64),
.B1(n_472),
.B2(n_473),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_68),
.A2(n_80),
.B1(n_81),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_75),
.C(n_78),
.Y(n_117)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_72),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_72),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_74),
.B(n_84),
.C(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_74),
.A2(n_78),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_75),
.Y(n_79)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_91),
.C(n_95),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_82),
.A2(n_83),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.C(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_84),
.A2(n_89),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_84),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_84),
.A2(n_162),
.B1(n_168),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_84),
.A2(n_162),
.B1(n_381),
.B2(n_386),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_84),
.B(n_386),
.Y(n_428)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_86),
.Y(n_379)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_86),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_87),
.A2(n_161),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_87),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_87),
.B(n_242),
.C(n_245),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_87),
.A2(n_164),
.B1(n_242),
.B2(n_305),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_89),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_91),
.A2(n_95),
.B1(n_96),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_94),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_94),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_95),
.A2(n_96),
.B1(n_172),
.B2(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_96),
.B(n_167),
.C(n_172),
.Y(n_166)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_115),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_113),
.C(n_114),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_103),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_102),
.B(n_228),
.C(n_233),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_102),
.A2(n_103),
.B1(n_228),
.B2(n_229),
.Y(n_268)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_103),
.B(n_121),
.C(n_127),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_123),
.Y(n_122)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_109),
.Y(n_112)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_128),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_117),
.B(n_118),
.C(n_128),
.Y(n_467)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_121),
.A2(n_122),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_121),
.A2(n_122),
.B1(n_151),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_204),
.C(n_208),
.Y(n_203)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_126),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_129),
.B(n_134),
.C(n_136),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_131),
.Y(n_136)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_144),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_139),
.B(n_142),
.CI(n_144),
.CON(n_217),
.SN(n_217)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_166),
.C(n_178),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_160),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_146),
.B(n_150),
.Y(n_289)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_157),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_151),
.Y(n_474)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_157),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_156),
.Y(n_258)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_160),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_178),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_168),
.B(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_168),
.A2(n_193),
.B1(n_276),
.B2(n_277),
.Y(n_347)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_170),
.Y(n_385)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_171),
.Y(n_376)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_176),
.Y(n_273)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_177),
.Y(n_371)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_217),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_183),
.B(n_217),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_184),
.B(n_186),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_188),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_202),
.C(n_214),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_189),
.B(n_291),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.C(n_200),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_190),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_194),
.B(n_200),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_202),
.B(n_214),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.C(n_212),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_208),
.Y(n_283)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_210),
.Y(n_262)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g489 ( 
.A(n_217),
.Y(n_489)
);

AOI221xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_353),
.B1(n_453),
.B2(n_458),
.C(n_459),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_293),
.C(n_297),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_220),
.A2(n_454),
.B(n_457),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_286),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_221),
.B(n_286),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_263),
.C(n_265),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_222),
.B(n_263),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_248),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_223),
.B(n_249),
.C(n_260),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.C(n_240),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_225),
.B(n_241),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_227),
.B(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_232),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_233),
.B(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_260),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_256),
.C(n_259),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_285),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_250),
.A2(n_252),
.B(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_259),
.Y(n_285)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_265),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_280),
.C(n_284),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_266),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.C(n_274),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_267),
.B(n_349),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_269),
.A2(n_274),
.B1(n_275),
.B2(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_270),
.B(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_290),
.C(n_292),
.Y(n_294)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_293),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_294),
.B(n_295),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_324),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_298),
.A2(n_455),
.B(n_456),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_322),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_299),
.B(n_322),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_320),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_320),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.C(n_311),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_306),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_308),
.B(n_390),
.Y(n_389)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_327),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.C(n_316),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_312),
.A2(n_313),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_351),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_325),
.B(n_351),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.C(n_348),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_326),
.B(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_328),
.B(n_348),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.C(n_346),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_329),
.B(n_444),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_332),
.A2(n_346),
.B1(n_347),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_332),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_338),
.C(n_343),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_333),
.A2(n_334),
.B1(n_343),
.B2(n_344),
.Y(n_432)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_338),
.B(n_432),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_448),
.B(n_452),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_434),
.B(n_447),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_421),
.B(n_433),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_397),
.B(n_420),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_387),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_358),
.B(n_387),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_372),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_359),
.B(n_373),
.C(n_380),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_366),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_360),
.B(n_367),
.C(n_369),
.Y(n_430)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_380),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_377),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_375),
.Y(n_409)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_381),
.Y(n_386)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.C(n_392),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_389),
.A2(n_392),
.B1(n_393),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_414),
.B(n_419),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_407),
.B(n_413),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_400),
.B(n_406),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_406),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_404),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_404),
.Y(n_415)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_405),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_416),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_423),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_429),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_430),
.C(n_431),
.Y(n_446)
);

BUFx24_ASAP7_75t_SL g488 ( 
.A(n_424),
.Y(n_488)
);

FAx1_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_427),
.CI(n_428),
.CON(n_424),
.SN(n_424)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_427),
.C(n_428),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_446),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_446),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_443),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_437),
.B(n_440),
.C(n_443),
.Y(n_449)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_441),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_449),
.B(n_450),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_486),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_466),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_475),
.B1(n_476),
.B2(n_485),
.Y(n_470)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_471),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_477),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_478),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_480),
.Y(n_479)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);


endmodule