module real_jpeg_18146_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_448),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_0),
.B(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_1),
.A2(n_44),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_1),
.A2(n_134),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_1),
.Y(n_164)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_1),
.A2(n_112),
.A3(n_175),
.B1(n_177),
.B2(n_180),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_1),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_1),
.B(n_137),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_1),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_1),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_2),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_3),
.A2(n_23),
.B1(n_59),
.B2(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_3),
.A2(n_62),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_L g220 ( 
.A1(n_3),
.A2(n_62),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_3),
.A2(n_62),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_4),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_4),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_5),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_6),
.A2(n_47),
.B1(n_234),
.B2(n_344),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_7),
.A2(n_54),
.B1(n_90),
.B2(n_93),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_7),
.A2(n_54),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_7),
.A2(n_54),
.B1(n_347),
.B2(n_349),
.Y(n_346)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_8),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_8),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_8),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_9),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_9),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_9),
.Y(n_179)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_10),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_12),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_145),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_144),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_55),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_19),
.B(n_55),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_32),
.B1(n_41),
.B2(n_51),
.Y(n_19)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_20),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_21),
.A2(n_32),
.B1(n_58),
.B2(n_63),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_21),
.A2(n_32),
.B1(n_58),
.B2(n_63),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_21),
.B(n_32),
.Y(n_374)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B(n_32),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_22),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_25),
.Y(n_22)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_32),
.A2(n_41),
.B(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_32),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_32)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_34),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_34),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_34),
.Y(n_331)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_38),
.Y(n_123)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_47),
.A2(n_105),
.B1(n_181),
.B2(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_48),
.B(n_64),
.Y(n_332)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_138),
.C(n_142),
.Y(n_55)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_56),
.B(n_138),
.CI(n_142),
.CON(n_165),
.SN(n_165)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_69),
.C(n_97),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_57),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_57),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_57),
.B(n_204),
.C(n_341),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_57),
.A2(n_154),
.B1(n_204),
.B2(n_226),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_57),
.B(n_299),
.C(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_57),
.A2(n_154),
.B1(n_299),
.B2(n_305),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_64),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_65),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_65),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_69),
.A2(n_98),
.B1(n_99),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_69),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_69),
.B(n_159),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_89),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_79),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_71),
.A2(n_79),
.B(n_316),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_71),
.A2(n_360),
.B(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2x1p5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_81),
.Y(n_80)
);

AO22x2_ASAP7_75t_L g212 ( 
.A1(n_72),
.A2(n_80),
.B1(n_213),
.B2(n_220),
.Y(n_212)
);

AO22x1_ASAP7_75t_L g230 ( 
.A1(n_72),
.A2(n_80),
.B1(n_213),
.B2(n_220),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_72),
.B(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_72),
.A2(n_89),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_75),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_76),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_76),
.Y(n_235)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_76),
.Y(n_237)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_76),
.Y(n_273)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_76),
.Y(n_348)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_80),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_84),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_84),
.Y(n_363)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_96),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_96),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_96),
.Y(n_225)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_109),
.B1(n_130),
.B2(n_137),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_100),
.A2(n_109),
.B1(n_137),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_101),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_124),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_110),
.A2(n_124),
.B1(n_161),
.B2(n_205),
.Y(n_204)
);

OA22x2_ASAP7_75t_L g299 ( 
.A1(n_110),
.A2(n_124),
.B1(n_161),
.B2(n_205),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_110),
.A2(n_124),
.B(n_161),
.Y(n_390)
);

NAND2x1p5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_124),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_119),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_124)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_127),
.Y(n_223)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_140),
.B(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_166),
.B(n_446),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_165),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_148),
.B(n_165),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.C(n_157),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_150),
.A2(n_158),
.B1(n_429),
.B2(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_150),
.Y(n_437)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_158),
.C(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_155),
.B(n_226),
.C(n_315),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_155),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_155),
.Y(n_429)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_156),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_156),
.A2(n_317),
.B1(n_389),
.B2(n_390),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_157),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_158),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g451 ( 
.A(n_165),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_425),
.B(n_443),
.Y(n_166)
);

AO221x1_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_336),
.B1(n_338),
.B2(n_418),
.C(n_424),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_309),
.B(n_335),
.Y(n_168)
);

AOI21x1_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_292),
.B(n_308),
.Y(n_169)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_241),
.B(n_291),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_228),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_172),
.B(n_228),
.Y(n_291)
);

XOR2x2_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_203),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_173),
.B(n_212),
.C(n_226),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_183),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_174),
.B(n_183),
.Y(n_295)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_191),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_184),
.A2(n_232),
.B1(n_233),
.B2(n_238),
.Y(n_231)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_185),
.B(n_192),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_214),
.B(n_217),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g371 ( 
.A(n_191),
.B(n_346),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_192),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g279 ( 
.A1(n_199),
.A2(n_233),
.B(n_280),
.Y(n_279)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_202),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_212),
.B1(n_226),
.B2(n_227),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_204),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_204),
.A2(n_226),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_211),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_212),
.A2(n_227),
.B1(n_244),
.B2(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_212),
.B(n_384),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_212),
.A2(n_227),
.B1(n_384),
.B2(n_411),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_213),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_213),
.B(n_358),
.Y(n_368)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_245),
.A3(n_249),
.B1(n_251),
.B2(n_256),
.Y(n_244)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.C(n_240),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_229),
.A2(n_230),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_229),
.B(n_295),
.C(n_297),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_229),
.A2(n_230),
.B1(n_342),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_240),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_230),
.B(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_231),
.B(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_231),
.B(n_282),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_231),
.A2(n_263),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_232),
.A2(n_343),
.B1(n_346),
.B2(n_352),
.Y(n_342)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI21x1_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_266),
.B(n_290),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_262),
.Y(n_242)
);

NOR2xp67_ASAP7_75t_SL g290 ( 
.A(n_243),
.B(n_262),
.Y(n_290)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_244),
.Y(n_288)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_263),
.B(n_322),
.Y(n_401)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_285),
.B(n_289),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_281),
.B(n_284),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_279),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_286),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_299),
.C(n_303),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_280),
.A2(n_343),
.B(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_307),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_307),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_297),
.B1(n_298),
.B2(n_306),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_305),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_299),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_299),
.A2(n_357),
.B(n_364),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_299),
.B(n_357),
.Y(n_364)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_311),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_312),
.B(n_319),
.C(n_320),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_402),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_391),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_376),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_339),
.B(n_376),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_355),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_340),
.B(n_356),
.C(n_365),
.Y(n_439)
);

XNOR2x1_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_378),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_342),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx12f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_365),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_364),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_364),
.A2(n_428),
.B1(n_432),
.B2(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_372),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_369),
.A2(n_370),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_370),
.A2(n_371),
.B1(n_373),
.B2(n_375),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_370),
.A2(n_375),
.B(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_373),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.C(n_382),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_379),
.Y(n_393)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_388),
.C(n_389),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_396),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_384),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_391),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_394),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_397),
.C(n_400),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_398),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_401),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_414),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_405),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_410),
.C(n_412),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_412),
.B2(n_413),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_414),
.B(n_421),
.Y(n_420)
);

NAND2x1_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_417),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_420),
.B(n_422),
.C(n_423),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_438),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_426),
.A2(n_444),
.B(n_445),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_435),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_435),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_432),
.C(n_433),
.Y(n_427)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_428),
.Y(n_442)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_441),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_440),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);


endmodule