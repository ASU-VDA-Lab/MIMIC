module real_aes_7605_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g177 ( .A1(n_0), .A2(n_178), .B(n_181), .C(n_185), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_1), .B(n_169), .Y(n_188) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_3), .B(n_179), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_4), .A2(n_142), .B(n_145), .C(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_5), .A2(n_137), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_6), .A2(n_137), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_7), .B(n_169), .Y(n_555) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_8), .A2(n_171), .B(n_243), .Y(n_242) );
AOI222xp33_ASAP7_75t_L g457 ( .A1(n_9), .A2(n_458), .B1(n_746), .B2(n_747), .C1(n_750), .C2(n_753), .Y(n_457) );
AND2x6_ASAP7_75t_L g142 ( .A(n_10), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_11), .A2(n_142), .B(n_145), .C(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g515 ( .A(n_12), .Y(n_515) );
INVx1_ASAP7_75t_L g107 ( .A(n_13), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_13), .B(n_40), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_14), .B(n_184), .Y(n_526) );
INVx1_ASAP7_75t_L g163 ( .A(n_15), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_16), .B(n_179), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_17), .B(n_454), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_18), .A2(n_180), .B(n_535), .C(n_537), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_19), .B(n_169), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_20), .B(n_157), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_21), .A2(n_145), .B(n_148), .C(n_156), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_22), .A2(n_183), .B(n_251), .C(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_23), .B(n_184), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_24), .B(n_184), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_25), .Y(n_496) );
INVx1_ASAP7_75t_L g476 ( .A(n_26), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_27), .A2(n_145), .B(n_156), .C(n_246), .Y(n_245) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_28), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_29), .Y(n_522) );
INVx1_ASAP7_75t_L g490 ( .A(n_30), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_31), .A2(n_137), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g140 ( .A(n_32), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_33), .A2(n_195), .B(n_196), .C(n_200), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_34), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_35), .A2(n_183), .B(n_552), .C(n_554), .Y(n_551) );
INVxp67_ASAP7_75t_L g491 ( .A(n_36), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_37), .B(n_248), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_38), .A2(n_145), .B(n_156), .C(n_475), .Y(n_474) );
CKINVDCx14_ASAP7_75t_R g550 ( .A(n_39), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_40), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_41), .A2(n_185), .B(n_513), .C(n_514), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_42), .B(n_136), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_43), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_44), .B(n_179), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_45), .B(n_137), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_46), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_47), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_48), .A2(n_195), .B(n_200), .C(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g182 ( .A(n_49), .Y(n_182) );
INVx1_ASAP7_75t_L g226 ( .A(n_50), .Y(n_226) );
INVx1_ASAP7_75t_L g563 ( .A(n_51), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_52), .B(n_137), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_53), .Y(n_165) );
CKINVDCx14_ASAP7_75t_R g511 ( .A(n_54), .Y(n_511) );
INVx1_ASAP7_75t_L g143 ( .A(n_55), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_56), .B(n_137), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_57), .B(n_169), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_58), .A2(n_155), .B(n_211), .C(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g162 ( .A(n_59), .Y(n_162) );
INVx1_ASAP7_75t_SL g553 ( .A(n_60), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_61), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_62), .B(n_179), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_63), .A2(n_102), .B1(n_113), .B2(n_757), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_64), .B(n_169), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_65), .B(n_180), .Y(n_261) );
INVx1_ASAP7_75t_L g499 ( .A(n_66), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_67), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_68), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_69), .A2(n_145), .B(n_200), .C(n_209), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_70), .Y(n_235) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_72), .A2(n_137), .B(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_73), .A2(n_93), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_73), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_74), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_75), .A2(n_137), .B(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_76), .A2(n_100), .B1(n_748), .B2(n_749), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_76), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_77), .A2(n_136), .B(n_486), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_78), .Y(n_473) );
INVx1_ASAP7_75t_L g533 ( .A(n_79), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_80), .B(n_153), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_81), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_82), .A2(n_137), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g536 ( .A(n_83), .Y(n_536) );
INVx2_ASAP7_75t_L g160 ( .A(n_84), .Y(n_160) );
INVx1_ASAP7_75t_L g525 ( .A(n_85), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_86), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_87), .B(n_184), .Y(n_262) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_88), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g449 ( .A(n_88), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g461 ( .A(n_88), .B(n_451), .Y(n_461) );
INVx2_ASAP7_75t_L g465 ( .A(n_88), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_89), .A2(n_145), .B(n_200), .C(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_90), .B(n_137), .Y(n_193) );
INVx1_ASAP7_75t_L g197 ( .A(n_91), .Y(n_197) );
INVxp67_ASAP7_75t_L g238 ( .A(n_92), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_93), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_94), .B(n_171), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_95), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g210 ( .A(n_96), .Y(n_210) );
INVx1_ASAP7_75t_L g257 ( .A(n_97), .Y(n_257) );
INVx2_ASAP7_75t_L g566 ( .A(n_98), .Y(n_566) );
AND2x2_ASAP7_75t_L g228 ( .A(n_99), .B(n_159), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_100), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_105), .Y(n_758) );
OR2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
AND2x2_ASAP7_75t_L g451 ( .A(n_109), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_456), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g756 ( .A(n_115), .Y(n_756) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_447), .B(n_453), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B1(n_124), .B2(n_125), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_124), .A2(n_459), .B1(n_462), .B2(n_466), .Y(n_458) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_125), .A2(n_459), .B1(n_754), .B2(n_755), .Y(n_753) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_402), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_337), .Y(n_126) );
NAND4xp25_ASAP7_75t_SL g127 ( .A(n_128), .B(n_282), .C(n_306), .D(n_329), .Y(n_127) );
AOI221xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_219), .B1(n_253), .B2(n_266), .C(n_269), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_189), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_131), .A2(n_167), .B1(n_220), .B2(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_131), .B(n_190), .Y(n_340) );
AND2x2_ASAP7_75t_L g359 ( .A(n_131), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_131), .B(n_343), .Y(n_429) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_167), .Y(n_131) );
AND2x2_ASAP7_75t_L g297 ( .A(n_132), .B(n_190), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_132), .B(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g320 ( .A(n_132), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g325 ( .A(n_132), .B(n_168), .Y(n_325) );
INVx2_ASAP7_75t_L g357 ( .A(n_132), .Y(n_357) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_132), .Y(n_401) );
AND2x2_ASAP7_75t_L g418 ( .A(n_132), .B(n_295), .Y(n_418) );
INVx5_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g336 ( .A(n_133), .B(n_295), .Y(n_336) );
AND2x4_ASAP7_75t_L g350 ( .A(n_133), .B(n_167), .Y(n_350) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_133), .Y(n_354) );
AND2x2_ASAP7_75t_L g374 ( .A(n_133), .B(n_289), .Y(n_374) );
AND2x2_ASAP7_75t_L g424 ( .A(n_133), .B(n_191), .Y(n_424) );
AND2x2_ASAP7_75t_L g434 ( .A(n_133), .B(n_168), .Y(n_434) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_164), .Y(n_133) );
AOI21xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_144), .B(n_157), .Y(n_134) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g258 ( .A(n_138), .B(n_142), .Y(n_258) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g155 ( .A(n_139), .Y(n_155) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx1_ASAP7_75t_L g252 ( .A(n_140), .Y(n_252) );
INVx1_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_141), .Y(n_151) );
INVx3_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
INVx1_ASAP7_75t_L g248 ( .A(n_141), .Y(n_248) );
BUFx3_ASAP7_75t_L g156 ( .A(n_142), .Y(n_156) );
INVx4_ASAP7_75t_SL g187 ( .A(n_142), .Y(n_187) );
INVx5_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx3_ASAP7_75t_L g186 ( .A(n_146), .Y(n_186) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_146), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .B(n_154), .Y(n_148) );
INVx2_ASAP7_75t_L g153 ( .A(n_150), .Y(n_153) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g196 ( .A1(n_153), .A2(n_197), .B(n_198), .C(n_199), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_153), .A2(n_199), .B(n_226), .C(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_153), .A2(n_499), .B(n_500), .C(n_501), .Y(n_498) );
O2A1O1Ixp5_ASAP7_75t_L g524 ( .A1(n_153), .A2(n_501), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_154), .A2(n_179), .B(n_476), .C(n_477), .Y(n_475) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_155), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_158), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g166 ( .A(n_159), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_159), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_159), .A2(n_223), .B(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_159), .A2(n_258), .B(n_473), .C(n_474), .Y(n_472) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_159), .A2(n_509), .B(n_516), .Y(n_508) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AND2x2_ASAP7_75t_L g172 ( .A(n_160), .B(n_161), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_166), .A2(n_521), .B(n_527), .Y(n_520) );
AND2x2_ASAP7_75t_L g290 ( .A(n_167), .B(n_190), .Y(n_290) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_167), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_167), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g380 ( .A(n_167), .Y(n_380) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g268 ( .A(n_168), .B(n_205), .Y(n_268) );
AND2x2_ASAP7_75t_L g295 ( .A(n_168), .B(n_206), .Y(n_295) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_173), .B(n_188), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_170), .B(n_202), .Y(n_201) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_170), .A2(n_207), .B(n_217), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_170), .B(n_218), .Y(n_217) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_170), .A2(n_256), .B(n_263), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_170), .B(n_479), .Y(n_478) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_170), .A2(n_495), .B(n_502), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_170), .B(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_171), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_171), .A2(n_244), .B(n_245), .Y(n_243) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g265 ( .A(n_172), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_187), .Y(n_174) );
INVx2_ASAP7_75t_L g195 ( .A(n_176), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_176), .A2(n_187), .B(n_235), .C(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_176), .A2(n_187), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_176), .A2(n_187), .B(n_511), .C(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_176), .A2(n_187), .B(n_533), .C(n_534), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_176), .A2(n_187), .B(n_550), .C(n_551), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_SL g562 ( .A1(n_176), .A2(n_187), .B(n_563), .C(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_179), .B(n_238), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_179), .A2(n_212), .B1(n_490), .B2(n_491), .Y(n_489) );
INVx5_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_180), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_183), .B(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g513 ( .A(n_184), .Y(n_513) );
INVx2_ASAP7_75t_L g501 ( .A(n_185), .Y(n_501) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_186), .Y(n_199) );
INVx1_ASAP7_75t_L g537 ( .A(n_186), .Y(n_537) );
INVx1_ASAP7_75t_L g200 ( .A(n_187), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_189), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_203), .Y(n_189) );
OR2x2_ASAP7_75t_L g321 ( .A(n_190), .B(n_204), .Y(n_321) );
AND2x2_ASAP7_75t_L g358 ( .A(n_190), .B(n_268), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_190), .B(n_289), .Y(n_369) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_190), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_190), .B(n_325), .Y(n_442) );
INVx5_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
BUFx2_ASAP7_75t_L g267 ( .A(n_191), .Y(n_267) );
AND2x2_ASAP7_75t_L g276 ( .A(n_191), .B(n_204), .Y(n_276) );
AND2x2_ASAP7_75t_L g392 ( .A(n_191), .B(n_287), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_191), .B(n_325), .Y(n_414) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_201), .Y(n_191) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_204), .Y(n_360) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_205), .Y(n_312) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
BUFx2_ASAP7_75t_L g289 ( .A(n_206), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_216), .Y(n_207) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_213), .C(n_214), .Y(n_209) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_212), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_212), .B(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g554 ( .A(n_215), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_229), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_220), .B(n_302), .Y(n_421) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_221), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g273 ( .A(n_221), .B(n_274), .Y(n_273) );
INVx5_ASAP7_75t_SL g281 ( .A(n_221), .Y(n_281) );
OR2x2_ASAP7_75t_L g304 ( .A(n_221), .B(n_274), .Y(n_304) );
OR2x2_ASAP7_75t_L g314 ( .A(n_221), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g377 ( .A(n_221), .B(n_231), .Y(n_377) );
AND2x2_ASAP7_75t_SL g415 ( .A(n_221), .B(n_230), .Y(n_415) );
NOR4xp25_ASAP7_75t_L g436 ( .A(n_221), .B(n_357), .C(n_437), .D(n_438), .Y(n_436) );
AND2x2_ASAP7_75t_L g446 ( .A(n_221), .B(n_278), .Y(n_446) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_228), .Y(n_221) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g271 ( .A(n_230), .B(n_267), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_230), .B(n_273), .Y(n_440) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_240), .Y(n_230) );
OR2x2_ASAP7_75t_L g280 ( .A(n_231), .B(n_281), .Y(n_280) );
INVx3_ASAP7_75t_L g287 ( .A(n_231), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_231), .B(n_255), .Y(n_299) );
INVxp67_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_231), .B(n_274), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_231), .B(n_241), .Y(n_368) );
AND2x2_ASAP7_75t_L g383 ( .A(n_231), .B(n_278), .Y(n_383) );
OR2x2_ASAP7_75t_L g412 ( .A(n_231), .B(n_241), .Y(n_412) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_239), .Y(n_231) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_232), .A2(n_531), .B(n_538), .Y(n_530) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_232), .A2(n_548), .B(n_555), .Y(n_547) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_232), .A2(n_561), .B(n_567), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_240), .B(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_240), .B(n_281), .Y(n_420) );
OR2x2_ASAP7_75t_L g441 ( .A(n_240), .B(n_318), .Y(n_441) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g254 ( .A(n_241), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g278 ( .A(n_241), .B(n_274), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_241), .B(n_255), .Y(n_293) );
AND2x2_ASAP7_75t_L g363 ( .A(n_241), .B(n_287), .Y(n_363) );
AND2x2_ASAP7_75t_L g397 ( .A(n_241), .B(n_281), .Y(n_397) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_242), .B(n_281), .Y(n_300) );
AND2x2_ASAP7_75t_L g328 ( .A(n_242), .B(n_255), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B(n_250), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_250), .A2(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_253), .B(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_254), .A2(n_343), .B1(n_379), .B2(n_396), .C(n_398), .Y(n_395) );
INVx5_ASAP7_75t_SL g274 ( .A(n_255), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_259), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_258), .A2(n_496), .B(n_497), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_258), .A2(n_522), .B(n_523), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g484 ( .A(n_265), .Y(n_484) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
OAI33xp33_ASAP7_75t_L g294 ( .A1(n_267), .A2(n_295), .A3(n_296), .B1(n_298), .B2(n_301), .B3(n_305), .Y(n_294) );
OR2x2_ASAP7_75t_L g310 ( .A(n_267), .B(n_311), .Y(n_310) );
AOI322xp5_ASAP7_75t_L g419 ( .A1(n_267), .A2(n_336), .A3(n_343), .B1(n_420), .B2(n_421), .C1(n_422), .C2(n_425), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_267), .B(n_295), .Y(n_437) );
A2O1A1Ixp33_ASAP7_75t_SL g443 ( .A1(n_267), .A2(n_295), .B(n_444), .C(n_446), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g282 ( .A1(n_268), .A2(n_283), .B1(n_288), .B2(n_291), .C(n_294), .Y(n_282) );
INVx1_ASAP7_75t_L g375 ( .A(n_268), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_268), .B(n_424), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_272), .B1(n_275), .B2(n_277), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g352 ( .A(n_273), .B(n_287), .Y(n_352) );
AND2x2_ASAP7_75t_L g410 ( .A(n_273), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g318 ( .A(n_274), .B(n_281), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_274), .B(n_287), .Y(n_346) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_276), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_276), .B(n_354), .Y(n_408) );
OAI321xp33_ASAP7_75t_L g427 ( .A1(n_276), .A2(n_349), .A3(n_428), .B1(n_429), .B2(n_430), .C(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g394 ( .A(n_277), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_278), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g333 ( .A(n_278), .B(n_281), .Y(n_333) );
AOI321xp33_ASAP7_75t_L g391 ( .A1(n_278), .A2(n_295), .A3(n_392), .B1(n_393), .B2(n_394), .C(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g308 ( .A(n_280), .B(n_293), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_281), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_281), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_281), .B(n_367), .Y(n_404) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g327 ( .A(n_285), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g292 ( .A(n_286), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g400 ( .A(n_287), .Y(n_400) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_290), .B(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g323 ( .A(n_295), .Y(n_323) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_297), .B(n_332), .Y(n_381) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
OR2x2_ASAP7_75t_L g345 ( .A(n_300), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g390 ( .A(n_300), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_301), .A2(n_348), .B1(n_351), .B2(n_353), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g445 ( .A(n_304), .B(n_368), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B1(n_313), .B2(n_319), .C(n_322), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g343 ( .A(n_312), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_SL g389 ( .A(n_315), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_317), .B(n_367), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_317), .A2(n_385), .B(n_387), .Y(n_384) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g430 ( .A(n_318), .B(n_412), .Y(n_430) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_SL g332 ( .A(n_321), .Y(n_332) );
AOI21xp33_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g376 ( .A(n_328), .B(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g438 ( .A(n_328), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B(n_334), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_332), .B(n_350), .Y(n_386) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g407 ( .A(n_336), .Y(n_407) );
NAND5xp2_ASAP7_75t_L g337 ( .A(n_338), .B(n_355), .C(n_364), .D(n_384), .E(n_391), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B(n_344), .C(n_347), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g379 ( .A(n_343), .Y(n_379) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_351), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
OAI21xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_359), .B(n_361), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_356), .A2(n_410), .B1(n_413), .B2(n_415), .C(n_416), .Y(n_409) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AOI321xp33_ASAP7_75t_L g364 ( .A1(n_357), .A2(n_365), .A3(n_369), .B1(n_370), .B2(n_376), .C(n_378), .Y(n_364) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g435 ( .A(n_369), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_371), .B(n_375), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g387 ( .A(n_372), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NOR2xp67_ASAP7_75t_SL g399 ( .A(n_373), .B(n_380), .Y(n_399) );
AOI321xp33_ASAP7_75t_SL g431 ( .A1(n_376), .A2(n_432), .A3(n_433), .B1(n_434), .B2(n_435), .C(n_436), .Y(n_431) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B(n_381), .C(n_382), .Y(n_378) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_389), .B(n_397), .Y(n_426) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND3xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .C(n_401), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_427), .C(n_439), .Y(n_402) );
OAI211xp5_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_405), .B(n_409), .C(n_419), .Y(n_403) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_407), .B(n_408), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_408), .A2(n_440), .B1(n_441), .B2(n_442), .C(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g428 ( .A(n_410), .Y(n_428) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g432 ( .A(n_430), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
CKINVDCx14_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g455 ( .A(n_449), .Y(n_455) );
NOR2x2_ASAP7_75t_L g752 ( .A(n_450), .B(n_465), .Y(n_752) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g464 ( .A(n_451), .B(n_465), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g456 ( .A1(n_453), .A2(n_457), .B(n_756), .Y(n_456) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g755 ( .A(n_463), .Y(n_755) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g754 ( .A(n_466), .Y(n_754) );
OR4x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_636), .C(n_683), .D(n_723), .Y(n_466) );
NAND3xp33_ASAP7_75t_SL g467 ( .A(n_468), .B(n_582), .C(n_611), .Y(n_467) );
AOI211xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_504), .B(n_539), .C(n_575), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_469), .A2(n_595), .B(n_612), .C(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_471), .B(n_574), .Y(n_573) );
INVx3_ASAP7_75t_SL g578 ( .A(n_471), .Y(n_578) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_471), .Y(n_590) );
AND2x4_ASAP7_75t_L g594 ( .A(n_471), .B(n_546), .Y(n_594) );
AND2x2_ASAP7_75t_L g605 ( .A(n_471), .B(n_494), .Y(n_605) );
OR2x2_ASAP7_75t_L g629 ( .A(n_471), .B(n_542), .Y(n_629) );
AND2x2_ASAP7_75t_L g642 ( .A(n_471), .B(n_547), .Y(n_642) );
AND2x2_ASAP7_75t_L g682 ( .A(n_471), .B(n_668), .Y(n_682) );
AND2x2_ASAP7_75t_L g689 ( .A(n_471), .B(n_652), .Y(n_689) );
AND2x2_ASAP7_75t_L g719 ( .A(n_471), .B(n_481), .Y(n_719) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_478), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_480), .B(n_646), .Y(n_658) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_493), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_481), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g596 ( .A(n_481), .B(n_493), .Y(n_596) );
BUFx3_ASAP7_75t_L g604 ( .A(n_481), .Y(n_604) );
OR2x2_ASAP7_75t_L g625 ( .A(n_481), .B(n_507), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_481), .B(n_646), .Y(n_736) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_485), .B(n_492), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_483), .A2(n_543), .B(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g543 ( .A(n_485), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_492), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_493), .B(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g589 ( .A(n_493), .Y(n_589) );
AND2x2_ASAP7_75t_L g652 ( .A(n_493), .B(n_547), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_493), .A2(n_655), .B1(n_657), .B2(n_659), .C(n_660), .Y(n_654) );
AND2x2_ASAP7_75t_L g668 ( .A(n_493), .B(n_542), .Y(n_668) );
AND2x2_ASAP7_75t_L g694 ( .A(n_493), .B(n_578), .Y(n_694) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g574 ( .A(n_494), .B(n_547), .Y(n_574) );
BUFx2_ASAP7_75t_L g708 ( .A(n_494), .Y(n_708) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OAI32xp33_ASAP7_75t_L g674 ( .A1(n_505), .A2(n_635), .A3(n_649), .B1(n_675), .B2(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .Y(n_505) );
AND2x2_ASAP7_75t_L g615 ( .A(n_506), .B(n_559), .Y(n_615) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g597 ( .A(n_507), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_507), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g669 ( .A(n_507), .B(n_559), .Y(n_669) );
AND2x2_ASAP7_75t_L g680 ( .A(n_507), .B(n_572), .Y(n_680) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g581 ( .A(n_508), .B(n_560), .Y(n_581) );
AND2x2_ASAP7_75t_L g585 ( .A(n_508), .B(n_560), .Y(n_585) );
AND2x2_ASAP7_75t_L g620 ( .A(n_508), .B(n_571), .Y(n_620) );
AND2x2_ASAP7_75t_L g627 ( .A(n_508), .B(n_529), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_508), .A2(n_578), .B(n_589), .C(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g686 ( .A(n_508), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_508), .B(n_519), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_517), .B(n_569), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_517), .B(n_585), .Y(n_675) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g580 ( .A(n_518), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_529), .Y(n_518) );
AND2x2_ASAP7_75t_L g572 ( .A(n_519), .B(n_530), .Y(n_572) );
OR2x2_ASAP7_75t_L g587 ( .A(n_519), .B(n_530), .Y(n_587) );
AND2x2_ASAP7_75t_L g610 ( .A(n_519), .B(n_571), .Y(n_610) );
INVx1_ASAP7_75t_L g614 ( .A(n_519), .Y(n_614) );
AND2x2_ASAP7_75t_L g633 ( .A(n_519), .B(n_570), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_519), .A2(n_598), .B1(n_644), .B2(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_519), .B(n_686), .Y(n_710) );
AND2x2_ASAP7_75t_L g725 ( .A(n_519), .B(n_585), .Y(n_725) );
INVx4_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx3_ASAP7_75t_L g557 ( .A(n_520), .Y(n_557) );
AND2x2_ASAP7_75t_L g599 ( .A(n_520), .B(n_530), .Y(n_599) );
AND2x2_ASAP7_75t_L g601 ( .A(n_520), .B(n_559), .Y(n_601) );
AND3x2_ASAP7_75t_L g663 ( .A(n_520), .B(n_627), .C(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g698 ( .A(n_529), .B(n_570), .Y(n_698) );
INVx1_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g559 ( .A(n_530), .B(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_530), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_530), .B(n_569), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_530), .B(n_610), .C(n_686), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_556), .B1(n_568), .B2(n_573), .Y(n_539) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_545), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_542), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g650 ( .A(n_542), .Y(n_650) );
OAI31xp33_ASAP7_75t_L g666 ( .A1(n_545), .A2(n_667), .A3(n_668), .B(n_669), .Y(n_666) );
AND2x2_ASAP7_75t_L g691 ( .A(n_545), .B(n_578), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_545), .B(n_604), .Y(n_737) );
AND2x2_ASAP7_75t_L g646 ( .A(n_546), .B(n_578), .Y(n_646) );
AND2x2_ASAP7_75t_L g707 ( .A(n_546), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g577 ( .A(n_547), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g635 ( .A(n_547), .Y(n_635) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
CKINVDCx16_ASAP7_75t_R g656 ( .A(n_557), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_558), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AOI221x1_ASAP7_75t_SL g623 ( .A1(n_559), .A2(n_624), .B1(n_626), .B2(n_628), .C(n_630), .Y(n_623) );
INVx2_ASAP7_75t_L g571 ( .A(n_560), .Y(n_571) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_560), .Y(n_665) );
INVx1_ASAP7_75t_L g653 ( .A(n_568), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_569), .B(n_586), .Y(n_678) );
INVx1_ASAP7_75t_SL g741 ( .A(n_569), .Y(n_741) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g659 ( .A(n_572), .B(n_585), .Y(n_659) );
INVx1_ASAP7_75t_L g727 ( .A(n_573), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_573), .B(n_656), .Y(n_740) );
INVx2_ASAP7_75t_SL g579 ( .A(n_574), .Y(n_579) );
AND2x2_ASAP7_75t_L g622 ( .A(n_574), .B(n_578), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_574), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_574), .B(n_649), .Y(n_676) );
AOI21xp33_ASAP7_75t_SL g575 ( .A1(n_576), .A2(n_579), .B(n_580), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_577), .B(n_649), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_577), .B(n_604), .Y(n_745) );
OR2x2_ASAP7_75t_L g617 ( .A(n_578), .B(n_596), .Y(n_617) );
AND2x2_ASAP7_75t_L g716 ( .A(n_578), .B(n_707), .Y(n_716) );
OAI22xp5_ASAP7_75t_SL g591 ( .A1(n_579), .A2(n_592), .B1(n_597), .B2(n_600), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_579), .B(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g639 ( .A(n_581), .B(n_587), .Y(n_639) );
INVx1_ASAP7_75t_L g703 ( .A(n_581), .Y(n_703) );
AOI311xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_588), .A3(n_590), .B(n_591), .C(n_602), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_586), .A2(n_718), .B1(n_730), .B2(n_733), .C(n_735), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_586), .B(n_741), .Y(n_743) );
INVx2_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g640 ( .A(n_588), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_589), .A2(n_631), .B(n_632), .C(n_634), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_SL g699 ( .A1(n_593), .A2(n_595), .B(n_700), .C(n_701), .Y(n_699) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_594), .B(n_668), .Y(n_734) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_597), .A2(n_617), .B1(n_618), .B2(n_621), .C(n_623), .Y(n_616) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g619 ( .A(n_599), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g702 ( .A(n_599), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_603), .A2(n_661), .B(n_662), .C(n_666), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_604), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_604), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g626 ( .A(n_610), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_614), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g728 ( .A(n_617), .Y(n_728) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_620), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g655 ( .A(n_620), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g732 ( .A(n_620), .Y(n_732) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g673 ( .A(n_622), .B(n_649), .Y(n_673) );
INVx1_ASAP7_75t_SL g667 ( .A(n_629), .Y(n_667) );
INVx1_ASAP7_75t_L g644 ( .A(n_635), .Y(n_644) );
NAND3xp33_ASAP7_75t_SL g636 ( .A(n_637), .B(n_654), .C(n_670), .Y(n_636) );
AOI322xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .A3(n_641), .B1(n_643), .B2(n_647), .C1(n_651), .C2(n_653), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g690 ( .A1(n_638), .A2(n_691), .B(n_692), .C(n_699), .Y(n_690) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_641), .A2(n_662), .B1(n_693), .B2(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g651 ( .A(n_649), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g688 ( .A(n_649), .B(n_689), .Y(n_688) );
AOI32xp33_ASAP7_75t_L g739 ( .A1(n_649), .A2(n_740), .A3(n_741), .B1(n_742), .B2(n_744), .Y(n_739) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g661 ( .A(n_652), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_652), .A2(n_705), .B1(n_709), .B2(n_711), .C(n_714), .Y(n_704) );
AND2x2_ASAP7_75t_L g718 ( .A(n_652), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g721 ( .A(n_656), .B(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g731 ( .A(n_656), .B(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g722 ( .A(n_665), .B(n_686), .Y(n_722) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .B(n_674), .C(n_677), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI211xp5_ASAP7_75t_SL g683 ( .A1(n_684), .A2(n_687), .B(n_690), .C(n_704), .Y(n_683) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_698), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g713 ( .A(n_710), .Y(n_713) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B(n_720), .Y(n_714) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OAI211xp5_ASAP7_75t_SL g723 ( .A1(n_724), .A2(n_726), .B(n_729), .C(n_739), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI21xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
endmodule