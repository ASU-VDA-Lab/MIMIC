module fake_jpeg_19919_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_60),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_48),
.B1(n_56),
.B2(n_55),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_43),
.B(n_44),
.C(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_49),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_38),
.B1(n_45),
.B2(n_44),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_46),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_81),
.B1(n_86),
.B2(n_5),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_65),
.B1(n_63),
.B2(n_62),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_53),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_2),
.C(n_3),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_51),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_1),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_88),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_99)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_20),
.A3(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_90)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_17),
.A3(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_96),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_87),
.B1(n_8),
.B2(n_7),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_99),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_105),
.B(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_79),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_103),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_76),
.B(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_109),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_106),
.B1(n_108),
.B2(n_91),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_111),
.B(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_114),
.B(n_94),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_12),
.B(n_13),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_15),
.C(n_18),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_21),
.B(n_25),
.C(n_26),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_27),
.Y(n_119)
);


endmodule