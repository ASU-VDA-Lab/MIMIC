module fake_netlist_1_1308_n_703 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_703);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_703;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g77 ( .A(n_76), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_46), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_34), .Y(n_79) );
BUFx3_ASAP7_75t_L g80 ( .A(n_59), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_54), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_47), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_35), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_13), .Y(n_84) );
CKINVDCx14_ASAP7_75t_R g85 ( .A(n_30), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_28), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_74), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_43), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_20), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_67), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_66), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_61), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_37), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_55), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_50), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_18), .Y(n_97) );
BUFx2_ASAP7_75t_SL g98 ( .A(n_49), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_23), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_12), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_60), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_14), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_42), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_70), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_68), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_40), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_65), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_27), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_56), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_8), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_38), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_25), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_39), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_26), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_12), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_36), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_14), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_71), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_21), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_69), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_16), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_72), .Y(n_124) );
INVxp33_ASAP7_75t_L g125 ( .A(n_20), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_117), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_78), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_78), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_117), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_112), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_77), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_84), .B(n_0), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_84), .B(n_1), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_125), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
BUFx8_ASAP7_75t_L g141 ( .A(n_95), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_89), .B(n_1), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_96), .B(n_2), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_80), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_95), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_86), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_102), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_91), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_91), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_102), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_86), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_92), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_89), .B(n_2), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_92), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_94), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_97), .B(n_3), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_97), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_101), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_100), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_101), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_96), .B(n_3), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_104), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_104), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_105), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_105), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_106), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_161), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
AND3x1_ASAP7_75t_L g173 ( .A(n_133), .B(n_100), .C(n_103), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_126), .B(n_114), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_126), .B(n_85), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
OR2x6_ASAP7_75t_L g177 ( .A(n_145), .B(n_98), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
AO22x2_ASAP7_75t_L g179 ( .A1(n_138), .A2(n_109), .B1(n_110), .B2(n_122), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_139), .A2(n_123), .B1(n_121), .B2(n_119), .Y(n_180) );
INVx4_ASAP7_75t_SL g181 ( .A(n_135), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_135), .Y(n_183) );
INVx4_ASAP7_75t_L g184 ( .A(n_135), .Y(n_184) );
NAND2x1p5_ASAP7_75t_L g185 ( .A(n_132), .B(n_109), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_130), .B(n_119), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_161), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_132), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_128), .B(n_124), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_162), .B(n_123), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_128), .B(n_88), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
BUFx4f_ASAP7_75t_L g196 ( .A(n_129), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_162), .B(n_121), .Y(n_197) );
NAND2x1_ASAP7_75t_L g198 ( .A(n_132), .B(n_122), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_146), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_146), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_161), .Y(n_204) );
BUFx10_ASAP7_75t_L g205 ( .A(n_129), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_159), .B(n_103), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_161), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_163), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
OAI22x1_ASAP7_75t_L g210 ( .A1(n_164), .A2(n_108), .B1(n_118), .B2(n_106), .Y(n_210) );
INVx8_ASAP7_75t_L g211 ( .A(n_140), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_133), .A2(n_169), .B1(n_168), .B2(n_167), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_131), .B(n_115), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_131), .B(n_134), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_134), .B(n_90), .Y(n_217) );
OAI21xp33_ASAP7_75t_L g218 ( .A1(n_142), .A2(n_87), .B(n_118), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_145), .B(n_98), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_140), .B(n_108), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_140), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_150), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_150), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_165), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_142), .B(n_93), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
INVx4_ASAP7_75t_L g229 ( .A(n_150), .Y(n_229) );
AND2x6_ASAP7_75t_L g230 ( .A(n_143), .B(n_110), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_165), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
OR2x6_ASAP7_75t_L g233 ( .A(n_137), .B(n_107), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_205), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_205), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_177), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_216), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_179), .A2(n_141), .B1(n_168), .B2(n_167), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_216), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_177), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_206), .Y(n_243) );
INVx5_ASAP7_75t_L g244 ( .A(n_205), .Y(n_244) );
NOR2xp33_ASAP7_75t_SL g245 ( .A(n_211), .B(n_81), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_211), .Y(n_246) );
BUFx12f_ASAP7_75t_L g247 ( .A(n_177), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_222), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_211), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_174), .B(n_141), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_222), .B(n_141), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_222), .B(n_141), .Y(n_252) );
BUFx12f_ASAP7_75t_L g253 ( .A(n_177), .Y(n_253) );
AO22x1_ASAP7_75t_L g254 ( .A1(n_206), .A2(n_116), .B1(n_111), .B2(n_113), .Y(n_254) );
INVx4_ASAP7_75t_L g255 ( .A(n_211), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_185), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_185), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_233), .A2(n_120), .B1(n_137), .B2(n_144), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_233), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_179), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_213), .B(n_169), .Y(n_261) );
INVx4_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_185), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_206), .B(n_166), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_233), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_196), .B(n_166), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_179), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_175), .B(n_148), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_179), .A2(n_148), .B1(n_160), .B2(n_143), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_220), .Y(n_270) );
AO22x1_ASAP7_75t_L g271 ( .A1(n_219), .A2(n_155), .B1(n_144), .B2(n_158), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_219), .B(n_155), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_233), .B(n_160), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_220), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_192), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_183), .Y(n_276) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_192), .B(n_158), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_173), .A2(n_153), .B1(n_157), .B2(n_156), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_183), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_220), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_190), .Y(n_281) );
INVx3_ASAP7_75t_L g282 ( .A(n_198), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_230), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_196), .B(n_157), .Y(n_284) );
BUFx4f_ASAP7_75t_L g285 ( .A(n_230), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_189), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_198), .Y(n_287) );
OR2x6_ASAP7_75t_L g288 ( .A(n_210), .B(n_156), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_195), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_182), .B(n_154), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_189), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_201), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_230), .Y(n_293) );
NOR2x1p5_ASAP7_75t_L g294 ( .A(n_197), .B(n_154), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_189), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_217), .B(n_153), .Y(n_296) );
AND2x4_ASAP7_75t_L g297 ( .A(n_197), .B(n_147), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_226), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_218), .B(n_99), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_186), .B(n_147), .Y(n_301) );
BUFx8_ASAP7_75t_SL g302 ( .A(n_186), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_189), .Y(n_303) );
INVxp67_ASAP7_75t_L g304 ( .A(n_275), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_260), .Y(n_305) );
AND2x6_ASAP7_75t_L g306 ( .A(n_263), .B(n_171), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_302), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_272), .B(n_172), .Y(n_308) );
BUFx2_ASAP7_75t_R g309 ( .A(n_302), .Y(n_309) );
OAI222xp33_ASAP7_75t_L g310 ( .A1(n_258), .A2(n_180), .B1(n_178), .B2(n_191), .C1(n_194), .C2(n_214), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_243), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_238), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_272), .A2(n_210), .B1(n_227), .B2(n_231), .C(n_196), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_240), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_260), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_235), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_259), .A2(n_230), .B1(n_184), .B2(n_107), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_244), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_255), .B(n_181), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_235), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_267), .A2(n_184), .B1(n_136), .B2(n_149), .Y(n_321) );
BUFx8_ASAP7_75t_L g322 ( .A(n_247), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_290), .A2(n_127), .B(n_136), .C(n_147), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_235), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_259), .A2(n_230), .B1(n_184), .B2(n_127), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_246), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_265), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_244), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_255), .B(n_181), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_265), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_241), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_267), .A2(n_230), .B1(n_163), .B2(n_136), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_263), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_255), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_272), .B(n_181), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_294), .A2(n_127), .B1(n_149), .B2(n_152), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_248), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_244), .B(n_149), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_263), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_244), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_297), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_256), .A2(n_152), .B1(n_229), .B2(n_224), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_248), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_297), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_257), .A2(n_152), .B1(n_229), .B2(n_224), .Y(n_346) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_245), .A2(n_151), .B1(n_229), .B2(n_224), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_247), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_263), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_246), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_301), .Y(n_351) );
INVxp67_ASAP7_75t_SL g352 ( .A(n_235), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_277), .B(n_151), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_253), .A2(n_151), .B1(n_199), .B2(n_187), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_301), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_270), .A2(n_151), .B1(n_199), .B2(n_234), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_301), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_334), .B(n_274), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_304), .A2(n_253), .B1(n_242), .B2(n_237), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_305), .A2(n_242), .B1(n_237), .B2(n_269), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_305), .A2(n_280), .B1(n_249), .B2(n_273), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_308), .B(n_271), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_313), .A2(n_268), .B(n_296), .C(n_250), .Y(n_363) );
INVx4_ASAP7_75t_SL g364 ( .A(n_306), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_311), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_308), .B(n_264), .Y(n_367) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_310), .A2(n_254), .B1(n_261), .B2(n_239), .C1(n_298), .C2(n_299), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_338), .B(n_278), .Y(n_369) );
NOR2xp33_ASAP7_75t_SL g370 ( .A(n_309), .B(n_285), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_323), .A2(n_193), .B(n_176), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_315), .B(n_288), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_312), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_330), .B(n_288), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g375 ( .A1(n_323), .A2(n_282), .B(n_287), .C(n_292), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_315), .A2(n_249), .B1(n_285), .B2(n_288), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_316), .Y(n_377) );
AOI21xp5_ASAP7_75t_SL g378 ( .A1(n_316), .A2(n_283), .B(n_236), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_327), .A2(n_288), .B1(n_300), .B2(n_284), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_334), .B(n_244), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_335), .A2(n_236), .B(n_252), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_316), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_306), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_337), .A2(n_236), .B(n_251), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_322), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_342), .A2(n_281), .B1(n_289), .B2(n_284), .C(n_266), .Y(n_386) );
NAND2x1p5_ASAP7_75t_L g387 ( .A(n_320), .B(n_246), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_345), .A2(n_266), .B1(n_287), .B2(n_282), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_318), .B(n_236), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_314), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_320), .Y(n_391) );
AOI222xp33_ASAP7_75t_L g392 ( .A1(n_367), .A2(n_307), .B1(n_322), .B2(n_355), .C1(n_351), .C2(n_357), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_368), .A2(n_322), .B1(n_353), .B2(n_331), .Y(n_393) );
OAI21xp5_ASAP7_75t_SL g394 ( .A1(n_360), .A2(n_332), .B(n_317), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_373), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_385), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_385), .Y(n_397) );
OA21x2_ASAP7_75t_L g398 ( .A1(n_375), .A2(n_212), .B(n_176), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_363), .A2(n_324), .B(n_320), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_372), .A2(n_362), .B1(n_374), .B2(n_379), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_390), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_370), .A2(n_325), .B1(n_336), .B2(n_285), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_365), .A2(n_347), .B1(n_348), .B2(n_321), .C(n_353), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_377), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_369), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_372), .A2(n_306), .B1(n_339), .B2(n_320), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_359), .A2(n_343), .B1(n_354), .B2(n_332), .C(n_339), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_374), .A2(n_339), .B1(n_306), .B2(n_282), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_380), .A2(n_306), .B1(n_287), .B2(n_337), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_358), .A2(n_306), .B1(n_324), .B2(n_318), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_361), .A2(n_328), .B1(n_341), .B2(n_324), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_358), .B(n_328), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_380), .A2(n_344), .B1(n_341), .B2(n_350), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_380), .A2(n_344), .B1(n_350), .B2(n_326), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_386), .A2(n_326), .B1(n_333), .B2(n_349), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_358), .A2(n_349), .B1(n_340), .B2(n_333), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_376), .A2(n_324), .B1(n_283), .B2(n_246), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_346), .B1(n_356), .B2(n_248), .C(n_293), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_381), .A2(n_151), .B1(n_349), .B2(n_340), .C(n_333), .Y(n_419) );
CKINVDCx6p67_ASAP7_75t_R g420 ( .A(n_383), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_393), .A2(n_383), .B1(n_387), .B2(n_389), .Y(n_421) );
OAI322xp33_ASAP7_75t_L g422 ( .A1(n_405), .A2(n_151), .A3(n_170), .B1(n_234), .B2(n_7), .C1(n_8), .C2(n_9), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_396), .B(n_340), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_420), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_405), .B(n_371), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_395), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_395), .B(n_371), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_404), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_392), .A2(n_400), .B1(n_403), .B2(n_407), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_397), .B(n_389), .Y(n_431) );
OR2x6_ASAP7_75t_L g432 ( .A(n_394), .B(n_378), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_401), .A2(n_371), .B1(n_384), .B2(n_170), .C(n_389), .Y(n_433) );
AO31x2_ASAP7_75t_L g434 ( .A1(n_399), .A2(n_377), .A3(n_382), .B(n_193), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_404), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
NAND4xp25_ASAP7_75t_L g437 ( .A(n_394), .B(n_188), .C(n_200), .D(n_203), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_398), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_408), .B(n_382), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_412), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_398), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_420), .B(n_366), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_411), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_398), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_398), .B(n_366), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_418), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_419), .B(n_391), .C(n_366), .Y(n_447) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_415), .A2(n_387), .B1(n_352), .B2(n_276), .C(n_279), .Y(n_448) );
OAI221xp5_ASAP7_75t_SL g449 ( .A1(n_402), .A2(n_378), .B1(n_215), .B2(n_188), .C(n_200), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_406), .A2(n_364), .B1(n_279), .B2(n_276), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_410), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_413), .A2(n_187), .B1(n_221), .B2(n_207), .C(n_204), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_416), .B(n_391), .C(n_228), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_417), .Y(n_454) );
INVx5_ASAP7_75t_L g455 ( .A(n_409), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_414), .A2(n_364), .B1(n_391), .B2(n_319), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_430), .A2(n_187), .B1(n_221), .B2(n_207), .C(n_204), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_428), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_429), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_426), .B(n_436), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g462 ( .A1(n_424), .A2(n_387), .B1(n_364), .B2(n_329), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_428), .B(n_364), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_422), .A2(n_221), .B1(n_207), .B2(n_204), .C(n_202), .Y(n_464) );
OAI31xp33_ASAP7_75t_L g465 ( .A1(n_424), .A2(n_329), .A3(n_319), .B(n_6), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_423), .B(n_203), .C(n_212), .D(n_215), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_424), .A2(n_329), .B1(n_319), .B2(n_283), .Y(n_467) );
OAI33xp33_ASAP7_75t_L g468 ( .A1(n_426), .A2(n_223), .A3(n_228), .B1(n_6), .B2(n_7), .B3(n_9), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_436), .B(n_4), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_440), .B(n_4), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_437), .B(n_223), .C(n_189), .Y(n_471) );
NAND4xp25_ASAP7_75t_L g472 ( .A(n_431), .B(n_5), .C(n_10), .D(n_11), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_432), .A2(n_283), .B1(n_262), .B2(n_293), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_435), .B(n_5), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_425), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_432), .B(n_10), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_427), .Y(n_479) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_437), .B(n_202), .C(n_208), .Y(n_480) );
AOI33xp33_ASAP7_75t_L g481 ( .A1(n_451), .A2(n_11), .A3(n_13), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_481) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_451), .B(n_202), .C(n_208), .Y(n_482) );
NAND2xp33_ASAP7_75t_SL g483 ( .A(n_442), .B(n_262), .Y(n_483) );
AOI222xp33_ASAP7_75t_L g484 ( .A1(n_446), .A2(n_15), .B1(n_17), .B2(n_18), .C1(n_19), .C2(n_21), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_442), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_455), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_446), .B(n_19), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_445), .Y(n_488) );
AOI32xp33_ASAP7_75t_L g489 ( .A1(n_421), .A2(n_293), .A3(n_262), .B1(n_32), .B2(n_33), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_445), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_438), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_443), .B(n_232), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_432), .B(n_22), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_439), .B(n_232), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_455), .B(n_232), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_438), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_432), .B(n_31), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_432), .B(n_41), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_441), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_441), .B(n_44), .Y(n_500) );
AOI33xp33_ASAP7_75t_L g501 ( .A1(n_456), .A2(n_303), .A3(n_295), .B1(n_291), .B2(n_286), .B3(n_53), .Y(n_501) );
AOI211xp5_ASAP7_75t_SL g502 ( .A1(n_422), .A2(n_45), .B(n_48), .C(n_51), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_444), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_455), .A2(n_202), .B1(n_232), .B2(n_209), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_444), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_455), .B(n_52), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_458), .B(n_455), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_458), .B(n_434), .Y(n_508) );
OAI21xp5_ASAP7_75t_SL g509 ( .A1(n_472), .A2(n_450), .B(n_447), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_490), .B(n_455), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_474), .B(n_434), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_474), .B(n_434), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_477), .B(n_434), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_481), .B(n_449), .C(n_433), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_490), .B(n_434), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_477), .B(n_454), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_460), .Y(n_517) );
INVx5_ASAP7_75t_L g518 ( .A(n_486), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_491), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_476), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_488), .B(n_454), .Y(n_521) );
BUFx2_ASAP7_75t_L g522 ( .A(n_486), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_485), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_469), .B(n_453), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_479), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_489), .A2(n_453), .B1(n_448), .B2(n_452), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_488), .B(n_57), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_491), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_463), .B(n_62), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_499), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_499), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_475), .Y(n_532) );
AOI31xp33_ASAP7_75t_SL g533 ( .A1(n_484), .A2(n_63), .A3(n_64), .B(n_73), .Y(n_533) );
AOI21xp5_ASAP7_75t_SL g534 ( .A1(n_480), .A2(n_75), .B(n_202), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_503), .Y(n_535) );
OAI31xp33_ASAP7_75t_L g536 ( .A1(n_465), .A2(n_286), .A3(n_291), .B(n_295), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_486), .B(n_208), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_475), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_463), .B(n_208), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_503), .B(n_208), .Y(n_540) );
NAND4xp25_ASAP7_75t_L g541 ( .A(n_465), .B(n_303), .C(n_209), .D(n_232), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_496), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_459), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_496), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_469), .B(n_209), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_459), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_461), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_505), .B(n_209), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_506), .B(n_209), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_505), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_461), .B(n_478), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_478), .B(n_493), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_493), .B(n_498), .Y(n_553) );
CKINVDCx16_ASAP7_75t_R g554 ( .A(n_483), .Y(n_554) );
NOR3xp33_ASAP7_75t_L g555 ( .A(n_470), .B(n_468), .C(n_487), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_497), .B(n_498), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_497), .B(n_506), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_494), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_500), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_500), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_495), .B(n_473), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_480), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_501), .B(n_504), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_471), .B(n_502), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_482), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_520), .B(n_489), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_519), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_523), .B(n_471), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_551), .B(n_482), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_519), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_517), .B(n_462), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_559), .B(n_466), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_551), .B(n_464), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_515), .B(n_457), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_528), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_515), .B(n_467), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_555), .B(n_466), .C(n_509), .D(n_556), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_522), .B(n_518), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_541), .A2(n_565), .B(n_534), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_507), .B(n_510), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_518), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_507), .B(n_510), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_521), .B(n_508), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_530), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_538), .B(n_532), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_530), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_521), .B(n_508), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_531), .B(n_535), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_525), .B(n_552), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_516), .B(n_511), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_522), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_531), .B(n_535), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_542), .B(n_544), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_516), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_543), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_544), .B(n_550), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_550), .B(n_511), .Y(n_599) );
NOR2xp67_ASAP7_75t_SL g600 ( .A(n_534), .B(n_554), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_512), .B(n_513), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_558), .B(n_553), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_514), .B(n_563), .C(n_564), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_543), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_546), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_512), .B(n_513), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_553), .B(n_524), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_529), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_546), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_547), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_547), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_560), .B(n_557), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_540), .Y(n_613) );
OR2x6_ASAP7_75t_L g614 ( .A(n_557), .B(n_549), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_561), .B(n_540), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_561), .B(n_539), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_579), .B(n_518), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_603), .B(n_564), .Y(n_618) );
OAI31xp33_ASAP7_75t_L g619 ( .A1(n_578), .A2(n_565), .A3(n_536), .B(n_526), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_590), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_590), .Y(n_621) );
INVx4_ASAP7_75t_L g622 ( .A(n_579), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_594), .Y(n_623) );
OAI211xp5_ASAP7_75t_L g624 ( .A1(n_580), .A2(n_529), .B(n_518), .C(n_562), .Y(n_624) );
OAI321xp33_ASAP7_75t_L g625 ( .A1(n_567), .A2(n_549), .A3(n_563), .B1(n_539), .B2(n_545), .C(n_562), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_579), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_591), .B(n_518), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_585), .B(n_566), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_594), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_581), .B(n_518), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_568), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_568), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_585), .B(n_566), .Y(n_633) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_593), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_589), .B(n_548), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_582), .B(n_549), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_571), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_581), .B(n_527), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_582), .B(n_537), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_589), .B(n_548), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_601), .B(n_537), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_587), .Y(n_642) );
NAND4xp25_ASAP7_75t_L g643 ( .A(n_572), .B(n_533), .C(n_537), .D(n_573), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_607), .Y(n_644) );
XNOR2x2_ASAP7_75t_L g645 ( .A(n_569), .B(n_602), .Y(n_645) );
XOR2xp5_ASAP7_75t_L g646 ( .A(n_612), .B(n_592), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_595), .Y(n_647) );
AOI211x1_ASAP7_75t_L g648 ( .A1(n_600), .A2(n_601), .B(n_606), .C(n_583), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_571), .Y(n_649) );
XOR2x2_ASAP7_75t_L g650 ( .A(n_583), .B(n_574), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_606), .B(n_596), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_576), .Y(n_652) );
AOI211xp5_ASAP7_75t_SL g653 ( .A1(n_608), .A2(n_600), .B(n_574), .C(n_570), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_577), .A2(n_575), .B(n_570), .C(n_613), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_614), .A2(n_613), .B1(n_616), .B2(n_577), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g656 ( .A1(n_575), .A2(n_615), .B(n_599), .C(n_586), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_599), .B(n_584), .Y(n_657) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_604), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g659 ( .A1(n_615), .A2(n_598), .B(n_595), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_584), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_597), .B(n_611), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_597), .B(n_611), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_605), .B(n_609), .Y(n_663) );
XNOR2xp5_ASAP7_75t_L g664 ( .A(n_614), .B(n_598), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_588), .Y(n_665) );
AOI221x1_ASAP7_75t_L g666 ( .A1(n_605), .A2(n_603), .B1(n_578), .B2(n_580), .C(n_555), .Y(n_666) );
A2O1A1Ixp33_ASAP7_75t_L g667 ( .A1(n_610), .A2(n_580), .B(n_556), .C(n_600), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_614), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_614), .B(n_601), .Y(n_669) );
OAI22x1_ASAP7_75t_L g670 ( .A1(n_617), .A2(n_622), .B1(n_646), .B2(n_639), .Y(n_670) );
NOR4xp25_ASAP7_75t_L g671 ( .A(n_618), .B(n_667), .C(n_642), .D(n_656), .Y(n_671) );
OAI222xp33_ASAP7_75t_L g672 ( .A1(n_622), .A2(n_617), .B1(n_655), .B2(n_664), .C1(n_639), .C2(n_618), .Y(n_672) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_658), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_622), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_663), .Y(n_675) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_666), .A2(n_619), .B(n_648), .C(n_653), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_630), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_650), .A2(n_624), .B(n_625), .Y(n_678) );
O2A1O1Ixp33_ASAP7_75t_L g679 ( .A1(n_643), .A2(n_634), .B(n_659), .C(n_644), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_636), .A2(n_627), .B(n_663), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_654), .A2(n_633), .B1(n_628), .B2(n_623), .C(n_620), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_633), .A2(n_628), .B1(n_621), .B2(n_629), .C(n_651), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_671), .A2(n_627), .B1(n_647), .B2(n_669), .C(n_668), .Y(n_683) );
AOI311xp33_ASAP7_75t_L g684 ( .A1(n_672), .A2(n_645), .A3(n_649), .B(n_631), .C(n_632), .Y(n_684) );
NAND4xp25_ASAP7_75t_SL g685 ( .A(n_676), .B(n_626), .C(n_645), .D(n_641), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_670), .A2(n_636), .B(n_662), .Y(n_686) );
OAI211xp5_ASAP7_75t_SL g687 ( .A1(n_678), .A2(n_657), .B(n_661), .C(n_662), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_674), .A2(n_635), .B1(n_640), .B2(n_638), .Y(n_688) );
OA22x2_ASAP7_75t_L g689 ( .A1(n_678), .A2(n_635), .B1(n_640), .B2(n_661), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_684), .A2(n_679), .B1(n_680), .B2(n_681), .C(n_673), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_689), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_683), .A2(n_682), .B(n_677), .C(n_675), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_688), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_686), .B1(n_685), .B2(n_687), .Y(n_694) );
XOR2xp5_ASAP7_75t_L g695 ( .A(n_691), .B(n_652), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_690), .A2(n_665), .B1(n_637), .B2(n_660), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_695), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_696), .Y(n_698) );
INVx2_ASAP7_75t_SL g699 ( .A(n_697), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_698), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_699), .Y(n_701) );
OAI21xp5_ASAP7_75t_SL g702 ( .A1(n_701), .A2(n_700), .B(n_699), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_702), .A2(n_694), .B(n_692), .Y(n_703) );
endmodule