module real_jpeg_11623_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

INVx4_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_70),
.B1(n_72),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_3),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_132),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_42),
.B1(n_47),
.B2(n_132),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_132),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_5),
.A2(n_42),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_5),
.A2(n_53),
.B1(n_59),
.B2(n_60),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_6),
.A2(n_38),
.B1(n_70),
.B2(n_72),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_38),
.B1(n_42),
.B2(n_47),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_6),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_7),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_7),
.B(n_78),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_7),
.B(n_30),
.C(n_46),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_7),
.A2(n_42),
.B1(n_47),
.B2(n_152),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_7),
.A2(n_35),
.B1(n_86),
.B2(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_7),
.B(n_108),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_11),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_11),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_11),
.A2(n_59),
.B1(n_60),
.B2(n_76),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_11),
.A2(n_42),
.B1(n_47),
.B2(n_76),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_76),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_12),
.A2(n_70),
.B1(n_72),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_12),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_12),
.A2(n_42),
.B1(n_47),
.B2(n_161),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_161),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_13),
.A2(n_42),
.B1(n_47),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_13),
.A2(n_50),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_14),
.A2(n_32),
.B1(n_59),
.B2(n_60),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_14),
.A2(n_32),
.B1(n_42),
.B2(n_47),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_32),
.B1(n_70),
.B2(n_72),
.Y(n_96)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_19),
.B(n_111),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_80),
.B2(n_81),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.C(n_66),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_22),
.A2(n_23),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_26),
.A2(n_35),
.B(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_28),
.B(n_35),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_29),
.A2(n_30),
.B1(n_44),
.B2(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_29),
.B(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_33),
.A2(n_34),
.B1(n_122),
.B2(n_148),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_33),
.A2(n_37),
.B(n_124),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_33),
.A2(n_34),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_35),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_35),
.B(n_152),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_35),
.A2(n_86),
.B1(n_236),
.B2(n_244),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_36),
.A2(n_86),
.B(n_238),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_39),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_40),
.A2(n_52),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_40),
.A2(n_89),
.B(n_103),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_40),
.A2(n_101),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_40),
.A2(n_51),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_40),
.A2(n_51),
.B1(n_210),
.B2(n_233),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_41)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

OA22x2_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_47),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_42),
.A2(n_57),
.B(n_205),
.C(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_42),
.B(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_SL g46 ( 
.A(n_44),
.Y(n_46)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_47),
.B(n_56),
.C(n_60),
.Y(n_206)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_48),
.A2(n_105),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_49),
.A2(n_51),
.B(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_51),
.B(n_152),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_66),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_61),
.Y(n_54)
);

AND2x4_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_55),
.B(n_63),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_55),
.A2(n_155),
.B1(n_156),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_55),
.A2(n_156),
.B1(n_173),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_65)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_58),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_73),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_59),
.B(n_72),
.C(n_73),
.Y(n_153)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_60),
.A2(n_69),
.B(n_151),
.C(n_153),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g205 ( 
.A(n_60),
.B(n_152),
.CON(n_205),
.SN(n_205)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_64),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_64),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_64),
.A2(n_108),
.B1(n_182),
.B2(n_205),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_75),
.B(n_77),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_67),
.A2(n_74),
.B1(n_75),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_67),
.A2(n_74),
.B1(n_131),
.B2(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_68)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_70),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g151 ( 
.A(n_72),
.B(n_152),
.CON(n_151),
.SN(n_151)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_78),
.A2(n_94),
.B1(n_151),
.B2(n_160),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_98),
.B2(n_99),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_88),
.B1(n_97),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_121),
.B(n_123),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_106),
.B(n_110),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_106),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_127),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_118),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.C(n_129),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_120),
.B(n_125),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_126),
.A2(n_129),
.B1(n_130),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_165),
.B(n_278),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_162),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_137),
.B(n_162),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_138),
.B(n_141),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_143),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_154),
.C(n_158),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_145),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_158),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B(n_157),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_193),
.B(n_273),
.C(n_277),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_186),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_176),
.C(n_179),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_168),
.B(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_171),
.C(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_185),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_187),
.B(n_191),
.C(n_192),
.Y(n_274)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_267),
.B(n_272),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_222),
.B(n_266),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_212),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_198),
.B(n_212),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.C(n_208),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_199),
.A2(n_200),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_207),
.B(n_208),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_213),
.B(n_218),
.C(n_220),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_260),
.B(n_265),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_250),
.B(n_259),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_239),
.B(n_249),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_234),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_245),
.B(n_248),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_257),
.C(n_258),
.Y(n_264)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_264),
.Y(n_265)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_271),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);


endmodule