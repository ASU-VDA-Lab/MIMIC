module real_jpeg_5432_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_0),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_0),
.A2(n_279),
.B1(n_374),
.B2(n_376),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_0),
.A2(n_87),
.B1(n_279),
.B2(n_408),
.Y(n_407)
);

OAI22xp33_ASAP7_75t_L g469 ( 
.A1(n_0),
.A2(n_279),
.B1(n_344),
.B2(n_470),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_1),
.A2(n_55),
.B1(n_100),
.B2(n_104),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_1),
.A2(n_55),
.B1(n_185),
.B2(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_1),
.A2(n_55),
.B1(n_422),
.B2(n_424),
.Y(n_421)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_2),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_2),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_2),
.Y(n_237)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_2),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_2),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_2),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_2),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_3),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_3),
.A2(n_49),
.B1(n_109),
.B2(n_112),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_49),
.B1(n_144),
.B2(n_147),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_3),
.A2(n_49),
.B1(n_315),
.B2(n_354),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_4),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_4),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_4),
.Y(n_443)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_4),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_5),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_5),
.B(n_140),
.C(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_5),
.B(n_88),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_5),
.B(n_201),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_5),
.B(n_142),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_5),
.B(n_111),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_6),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_6),
.A2(n_186),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g369 ( 
.A1(n_6),
.A2(n_186),
.B1(n_305),
.B2(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_6),
.A2(n_186),
.B1(n_344),
.B2(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_7),
.Y(n_336)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_8),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_9),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_9),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_9),
.A2(n_173),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_9),
.A2(n_173),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_9),
.A2(n_48),
.B1(n_173),
.B2(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_10),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_11),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_12),
.Y(n_135)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_12),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_13),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_13),
.A2(n_72),
.B1(n_314),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_13),
.A2(n_72),
.B1(n_399),
.B2(n_401),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_13),
.A2(n_72),
.B1(n_455),
.B2(n_457),
.Y(n_454)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_14),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_15),
.A2(n_40),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_15),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_15),
.A2(n_67),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_15),
.A2(n_67),
.B1(n_211),
.B2(n_395),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_15),
.A2(n_67),
.B1(n_270),
.B2(n_413),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_16),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_16),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_16),
.A2(n_212),
.B1(n_230),
.B2(n_233),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_16),
.A2(n_212),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_16),
.A2(n_65),
.B1(n_212),
.B2(n_442),
.Y(n_441)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_18),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_547),
.B(n_549),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_58),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_50),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_24),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_24),
.B(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_25)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_26),
.Y(n_338)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_33),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_33),
.Y(n_271)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_36),
.A2(n_361),
.B(n_362),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_36),
.B(n_364),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_50)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_48),
.Y(n_366)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_48),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_50),
.B(n_60),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_56),
.B1(n_64),
.B2(n_68),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_51),
.A2(n_52),
.B1(n_56),
.B2(n_68),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_51),
.A2(n_363),
.B(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_51),
.A2(n_56),
.B1(n_416),
.B2(n_441),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_51),
.A2(n_56),
.B1(n_64),
.B2(n_519),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_56),
.B(n_168),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_56),
.A2(n_441),
.B(n_473),
.Y(n_483)
);

AO21x1_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_155),
.B(n_546),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_151),
.C(n_152),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_61),
.A2(n_62),
.B1(n_542),
.B2(n_543),
.Y(n_541)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_73),
.C(n_116),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_63),
.B(n_534),
.Y(n_533)
);

OAI21xp33_ASAP7_75t_SL g361 ( 
.A1(n_65),
.A2(n_168),
.B(n_341),
.Y(n_361)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_73),
.A2(n_116),
.B1(n_117),
.B2(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_73),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_99),
.B1(n_107),
.B2(n_108),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_74),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_74),
.A2(n_107),
.B1(n_301),
.B2(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_74),
.A2(n_107),
.B1(n_407),
.B2(n_412),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_74),
.A2(n_99),
.B1(n_107),
.B2(n_523),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_88),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_80),
.B1(n_84),
.B2(n_86),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_83),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_83),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_83),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_SL g290 ( 
.A(n_84),
.B(n_146),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_88),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_88),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

AOI22x1_ASAP7_75t_L g444 ( 
.A1(n_88),
.A2(n_153),
.B1(n_309),
.B2(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_88),
.A2(n_153),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_96),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g213 ( 
.A(n_90),
.Y(n_213)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_92),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_92),
.Y(n_400)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_94),
.Y(n_375)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_98),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_103),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_103),
.Y(n_414)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_107),
.B(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_107),
.A2(n_301),
.B(n_308),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_115),
.Y(n_265)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_115),
.Y(n_330)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_115),
.Y(n_340)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_115),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_116),
.A2(n_117),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_116),
.B(n_518),
.C(n_521),
.Y(n_529)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_141),
.B(n_143),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_118),
.A2(n_165),
.B(n_169),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_118),
.A2(n_141),
.B1(n_210),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_118),
.A2(n_169),
.B(n_258),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_118),
.A2(n_141),
.B1(n_373),
.B2(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_119),
.B(n_170),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_119),
.A2(n_142),
.B1(n_394),
.B2(n_398),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_119),
.A2(n_142),
.B1(n_398),
.B2(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_119),
.A2(n_142),
.B1(n_421),
.B2(n_460),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_130),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_123),
.Y(n_397)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_SL g211 ( 
.A(n_129),
.Y(n_211)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_130),
.A2(n_210),
.B(n_214),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_133),
.B1(n_136),
.B2(n_139),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_137),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_141),
.A2(n_214),
.B(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_143),
.Y(n_460)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_146),
.Y(n_423)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_149),
.Y(n_286)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_150),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_151),
.B(n_152),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_153),
.A2(n_264),
.B(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_153),
.B(n_309),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_153),
.A2(n_268),
.B(n_486),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_540),
.B(n_545),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_512),
.B(n_537),
.Y(n_156)
);

OAI311xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_379),
.A3(n_488),
.B1(n_506),
.C1(n_511),
.Y(n_157)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_321),
.B(n_378),
.Y(n_158)
);

AO21x1_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_292),
.B(n_320),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_252),
.B(n_291),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_217),
.B(n_251),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_182),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_163),
.B(n_182),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_175),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_164),
.A2(n_175),
.B1(n_176),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_164),
.Y(n_249)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_168),
.A2(n_192),
.B(n_199),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_SL g264 ( 
.A1(n_168),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_168),
.B(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_174),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

INVx3_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_178),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_180),
.Y(n_316)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_207),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_183),
.B(n_208),
.C(n_216),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_192),
.B(n_199),
.Y(n_183)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_191),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_192),
.A2(n_347),
.B1(n_348),
.B2(n_351),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_192),
.A2(n_385),
.B1(n_389),
.B2(n_392),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_192),
.A2(n_392),
.B(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_202),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_193),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_193),
.A2(n_275),
.B1(n_313),
.B2(n_317),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_193),
.A2(n_352),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_205),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_215),
.B2(n_216),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_241),
.B(n_250),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_227),
.B(n_240),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx8_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_239),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_239),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_235),
.B(n_238),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_237),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_274),
.B(n_281),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_248),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_248),
.Y(n_250)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_247),
.Y(n_350)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_247),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_254),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_272),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_262),
.B2(n_263),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_262),
.C(n_272),
.Y(n_293)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI32xp33_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_283),
.A3(n_284),
.B1(n_287),
.B2(n_290),
.Y(n_282)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_271),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_282),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_282),
.Y(n_298)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx8_ASAP7_75t_L g354 ( 
.A(n_278),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_293),
.B(n_294),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_299),
.B2(n_319),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_298),
.C(n_319),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_299),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_310),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_300),
.B(n_311),
.C(n_312),
.Y(n_355)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_304),
.Y(n_456)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_322),
.B(n_323),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_358),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_324)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_345),
.B2(n_346),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_327),
.B(n_345),
.Y(n_484)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_331),
.A3(n_334),
.B1(n_337),
.B2(n_341),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_355),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_355),
.B(n_356),
.C(n_358),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_367),
.B2(n_377),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_359),
.B(n_368),
.C(n_372),
.Y(n_497)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_367),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_372),
.Y(n_367)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_369),
.Y(n_486)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_474),
.Y(n_379)
);

A2O1A1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_380),
.A2(n_474),
.B(n_507),
.C(n_510),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_446),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_381),
.B(n_446),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_418),
.C(n_431),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_382),
.B(n_418),
.CI(n_431),
.CON(n_487),
.SN(n_487)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_405),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_383),
.B(n_406),
.C(n_415),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_393),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_384),
.B(n_393),
.Y(n_480)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_394),
.Y(n_434)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx8_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_415),
.Y(n_405)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_412),
.Y(n_453)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_420),
.B1(n_426),
.B2(n_430),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_420),
.B(n_426),
.Y(n_464)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_426),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_426),
.A2(n_430),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_426),
.A2(n_464),
.B(n_467),
.Y(n_515)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_439),
.C(n_444),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_432),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_435),
.Y(n_496)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_439),
.A2(n_440),
.B1(n_444),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_444),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_447),
.B(n_450),
.C(n_462),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_462),
.B2(n_463),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_458),
.B(n_461),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_459),
.Y(n_461)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_454),
.Y(n_523)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_461),
.B(n_515),
.CI(n_516),
.CON(n_514),
.SN(n_514)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_461),
.B(n_515),
.C(n_516),
.Y(n_536)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_473),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_469),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_471),
.Y(n_470)
);

INVx8_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_487),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_487),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.C(n_481),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_476),
.A2(n_477),
.B1(n_480),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.C(n_485),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_482),
.A2(n_483),
.B1(n_485),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_485),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g553 ( 
.A(n_487),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_501),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_508),
.B(n_509),
.Y(n_507)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_498),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_498),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_495),
.C(n_497),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_504),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_495),
.A2(n_496),
.B1(n_497),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_497),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_503),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_526),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_525),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_525),
.Y(n_538)
);

BUFx24_ASAP7_75t_SL g555 ( 
.A(n_514),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_518),
.B1(n_520),
.B2(n_524),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_517),
.A2(n_518),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_517),
.B(n_528),
.C(n_532),
.Y(n_544)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_520),
.Y(n_524)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_526),
.A2(n_538),
.B(n_539),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_527),
.B(n_536),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_536),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_528),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_544),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_541),
.B(n_544),
.Y(n_545)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx13_ASAP7_75t_L g551 ( 
.A(n_548),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_552),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);


endmodule