module fake_jpeg_21200_n_324 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_11),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_18),
.B1(n_14),
.B2(n_20),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_27),
.B1(n_33),
.B2(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_56),
.Y(n_67)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_54),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_26),
.B(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_43),
.B1(n_27),
.B2(n_35),
.Y(n_70)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_45),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_48),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_59),
.Y(n_76)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_70),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_36),
.B1(n_42),
.B2(n_40),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_36),
.B1(n_55),
.B2(n_39),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_60),
.B1(n_57),
.B2(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_52),
.C(n_53),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_39),
.B1(n_36),
.B2(n_29),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_78),
.B1(n_72),
.B2(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_53),
.Y(n_89)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_38),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_86),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_90),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_53),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_59),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_97),
.Y(n_100)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_59),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_66),
.B1(n_63),
.B2(n_70),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_118),
.B1(n_93),
.B2(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_63),
.B(n_74),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_74),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_76),
.Y(n_114)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_38),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_78),
.B(n_72),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_63),
.B1(n_62),
.B2(n_73),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_63),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_24),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_73),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_91),
.B1(n_55),
.B2(n_75),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_124),
.A2(n_125),
.B1(n_138),
.B2(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_115),
.B1(n_121),
.B2(n_107),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_136),
.B1(n_146),
.B2(n_135),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_87),
.C(n_89),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_133),
.C(n_30),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_87),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_134),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_77),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_132),
.A2(n_144),
.B(n_31),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_75),
.B1(n_36),
.B2(n_55),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_75),
.B1(n_88),
.B2(n_46),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_46),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_16),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_46),
.Y(n_142)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_60),
.B1(n_68),
.B2(n_57),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_48),
.B(n_101),
.C(n_44),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_45),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_98),
.A2(n_17),
.B1(n_16),
.B2(n_22),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_49),
.B1(n_54),
.B2(n_46),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_54),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_156),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_41),
.B1(n_49),
.B2(n_60),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_20),
.B1(n_31),
.B2(n_32),
.Y(n_180)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_41),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_57),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_117),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_161),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_139),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_119),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_164),
.B(n_177),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_179),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_119),
.B1(n_120),
.B2(n_113),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_174),
.B1(n_178),
.B2(n_183),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_171),
.B(n_143),
.C(n_45),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_SL g171 ( 
.A1(n_152),
.A2(n_101),
.B(n_45),
.C(n_31),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_144),
.B(n_132),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_175),
.C(n_184),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_30),
.B1(n_18),
.B2(n_17),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_131),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_30),
.B1(n_18),
.B2(n_20),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_154),
.B1(n_147),
.B2(n_153),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_136),
.A2(n_18),
.B1(n_16),
.B2(n_22),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_31),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_24),
.C(n_45),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_187),
.C(n_45),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_25),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_126),
.A2(n_22),
.B1(n_13),
.B2(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_128),
.Y(n_191)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_141),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_205),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_126),
.B(n_148),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_197),
.B1(n_168),
.B2(n_171),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_206),
.B1(n_207),
.B2(n_12),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_32),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_209),
.B(n_44),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_132),
.C(n_144),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_161),
.C(n_159),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_143),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_179),
.A2(n_15),
.B1(n_44),
.B2(n_13),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_176),
.B1(n_168),
.B2(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_212),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_19),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_44),
.B1(n_32),
.B2(n_25),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_237),
.Y(n_251)
);

OAI22x1_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_171),
.B1(n_184),
.B2(n_187),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_206),
.B1(n_211),
.B2(n_193),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_229),
.B1(n_207),
.B2(n_198),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_24),
.C(n_11),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_230),
.C(n_11),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_24),
.C(n_11),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_233),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_13),
.B1(n_12),
.B2(n_15),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_235),
.Y(n_247)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_25),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_201),
.B1(n_213),
.B2(n_200),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_239),
.A2(n_246),
.B1(n_231),
.B2(n_230),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_214),
.B(n_210),
.Y(n_241)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_244),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_218),
.A2(n_199),
.B1(n_202),
.B2(n_204),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_219),
.A2(n_212),
.B1(n_197),
.B2(n_203),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_254),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_256),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_19),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_255),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_9),
.B(n_10),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_9),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_216),
.A2(n_15),
.B1(n_44),
.B2(n_19),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_227),
.B1(n_222),
.B2(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_267),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_237),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_264),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_215),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_228),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_269),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_232),
.B1(n_217),
.B2(n_229),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_21),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_221),
.Y(n_269)
);

AOI221xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_44),
.B1(n_7),
.B2(n_8),
.C(n_5),
.Y(n_271)
);

NOR3xp33_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_254),
.C(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_282),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_284),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_239),
.C(n_238),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_280),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_270),
.A2(n_245),
.B(n_246),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_258),
.Y(n_281)
);

XOR2x2_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_5),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_242),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_256),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_285),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_257),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_272),
.A2(n_15),
.B1(n_6),
.B2(n_10),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_5),
.B(n_8),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_261),
.C(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_292),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_273),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

AOI221xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_282),
.B1(n_6),
.B2(n_8),
.C(n_4),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_21),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_298),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_21),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_23),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_21),
.Y(n_298)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_308),
.B(n_3),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_6),
.B1(n_21),
.B2(n_23),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_21),
.C(n_23),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_309),
.C(n_289),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_23),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_289),
.B(n_1),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_312),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_0),
.C(n_1),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_306),
.B(n_304),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_315),
.A2(n_300),
.B(n_3),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_316),
.B(n_317),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_3),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_3),
.C(n_4),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_4),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_4),
.B(n_306),
.Y(n_324)
);


endmodule