module fake_jpeg_26371_n_82 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_82);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_82;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx4_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_22),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_19),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_20),
.C(n_21),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_20),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_17),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_18),
.B1(n_22),
.B2(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_36),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_37),
.B1(n_23),
.B2(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

OAI32xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_40),
.A3(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_27),
.C(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_8),
.B1(n_14),
.B2(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

OA21x2_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_12),
.B(n_14),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_51),
.B1(n_39),
.B2(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_49),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_11),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AO22x2_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_60),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_34),
.C(n_50),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_42),
.B1(n_46),
.B2(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_56),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_46),
.B(n_51),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_57),
.B(n_56),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_72),
.B1(n_48),
.B2(n_54),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_62),
.B1(n_63),
.B2(n_37),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_1),
.C(n_2),
.Y(n_76)
);

OAI31xp33_ASAP7_75t_L g78 ( 
.A1(n_74),
.A2(n_75),
.A3(n_1),
.B(n_2),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_40),
.Y(n_75)
);

MAJx2_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_73),
.C(n_7),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_78),
.C(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_4),
.Y(n_81)
);

AOI321xp33_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_78),
.C(n_13),
.Y(n_82)
);


endmodule