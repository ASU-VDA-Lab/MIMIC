module fake_jpeg_27531_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_44),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_46),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_24),
.Y(n_67)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_31),
.B(n_2),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_29),
.B(n_3),
.C(n_4),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_61),
.B1(n_69),
.B2(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_63),
.Y(n_76)
);

OA21x2_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_27),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_15),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_28),
.B1(n_30),
.B2(n_27),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_69),
.B1(n_0),
.B2(n_3),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_15),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_30),
.B1(n_23),
.B2(n_25),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_74),
.B1(n_6),
.B2(n_7),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_38),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_75),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_41),
.A2(n_32),
.B1(n_20),
.B2(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_34),
.B(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_86),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_90),
.Y(n_110)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_29),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_91),
.B1(n_58),
.B2(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_0),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_4),
.C(n_5),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_6),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_5),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_98),
.B1(n_66),
.B2(n_52),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_9),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_11),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_97),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_6),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_58),
.A3(n_65),
.B1(n_51),
.B2(n_57),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_107),
.B1(n_112),
.B2(n_94),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_71),
.B1(n_57),
.B2(n_73),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_108),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_131)
);

XOR2x2_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_62),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_115),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_73),
.B1(n_62),
.B2(n_68),
.Y(n_114)
);

OAI22x1_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_66),
.B1(n_64),
.B2(n_53),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_13),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_122),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_79),
.B(n_90),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_132),
.B(n_134),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_124),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_78),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_81),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_89),
.C(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_95),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_115),
.C(n_104),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_94),
.B(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_111),
.B1(n_114),
.B2(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_137),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_106),
.B(n_83),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_142),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_129),
.C(n_120),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_124),
.A2(n_112),
.B1(n_83),
.B2(n_99),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_132),
.B1(n_133),
.B2(n_121),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_103),
.B1(n_77),
.B2(n_92),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_151),
.C(n_154),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_140),
.B1(n_136),
.B2(n_85),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_156),
.Y(n_161)
);

NAND2x1_ASAP7_75t_SL g153 ( 
.A(n_138),
.B(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_64),
.B(n_13),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_125),
.C(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_143),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_160),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_150),
.A2(n_153),
.B1(n_142),
.B2(n_155),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_151),
.B(n_147),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_148),
.Y(n_166)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_167),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_161),
.B(n_154),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_159),
.B(n_162),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_171),
.B1(n_163),
.B2(n_14),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_160),
.B(n_161),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_164),
.Y(n_172)
);

AOI21x1_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_159),
.B(n_163),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_174),
.C(n_170),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_14),
.C(n_64),
.Y(n_176)
);


endmodule