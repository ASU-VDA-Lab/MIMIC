module real_jpeg_7350_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_323;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_0),
.A2(n_90),
.B1(n_92),
.B2(n_94),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_0),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_0),
.A2(n_94),
.B1(n_127),
.B2(n_131),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_0),
.A2(n_94),
.B1(n_416),
.B2(n_417),
.Y(n_415)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_1),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_1),
.Y(n_223)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_1),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_1),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_1),
.Y(n_449)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_2),
.Y(n_143)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_2),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_2),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_3),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_3),
.A2(n_54),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_3),
.A2(n_54),
.B1(n_420),
.B2(n_421),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_3),
.A2(n_54),
.B1(n_92),
.B2(n_430),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_4),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_4),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_4),
.A2(n_154),
.B1(n_226),
.B2(n_304),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_4),
.A2(n_154),
.B1(n_399),
.B2(n_401),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_4),
.A2(n_154),
.B1(n_293),
.B2(n_428),
.Y(n_427)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_180),
.B1(n_183),
.B2(n_187),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_6),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_6),
.B(n_197),
.C(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_6),
.B(n_74),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_6),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_6),
.B(n_125),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_6),
.B(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_7),
.Y(n_533)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_8),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_9),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_9),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_9),
.A2(n_87),
.B1(n_139),
.B2(n_144),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_9),
.A2(n_87),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_9),
.A2(n_87),
.B1(n_420),
.B2(n_437),
.Y(n_436)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_11),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_12),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_12),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_12),
.A2(n_210),
.B1(n_235),
.B2(n_257),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_12),
.A2(n_235),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_12),
.A2(n_51),
.B1(n_235),
.B2(n_453),
.Y(n_452)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_15),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_16),
.A2(n_204),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_16),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_16),
.A2(n_195),
.B1(n_208),
.B2(n_283),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_16),
.A2(n_91),
.B1(n_208),
.B2(n_298),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_16),
.A2(n_51),
.B1(n_53),
.B2(n_208),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_17),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_17),
.A2(n_62),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_17),
.A2(n_62),
.B1(n_206),
.B2(n_344),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_17),
.A2(n_62),
.B1(n_131),
.B2(n_424),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_18),
.A2(n_110),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_18),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_18),
.A2(n_190),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_18),
.A2(n_85),
.B1(n_190),
.B2(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_18),
.A2(n_190),
.B1(n_388),
.B2(n_393),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_532),
.B(n_534),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_169),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_167),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_145),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_23),
.B(n_145),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_132),
.B2(n_133),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_63),
.C(n_95),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_26),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_27),
.A2(n_55),
.B1(n_57),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_27),
.A2(n_50),
.B1(n_55),
.B2(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_27),
.A2(n_391),
.B(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_27),
.A2(n_55),
.B1(n_432),
.B2(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_28),
.A2(n_387),
.B(n_390),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_28),
.B(n_392),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g364 ( 
.A(n_32),
.Y(n_364)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B1(n_44),
.B2(n_48),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_39),
.Y(n_366)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_42),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_43),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_43),
.Y(n_290)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_43),
.Y(n_299)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_43),
.Y(n_337)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_47),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_47),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_53),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_55),
.B(n_187),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_55),
.A2(n_452),
.B(n_477),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_56),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_56),
.B(n_153),
.Y(n_476)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_59),
.Y(n_373)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_63),
.A2(n_95),
.B1(n_96),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_64),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_64),
.A2(n_82),
.B1(n_88),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_64),
.A2(n_88),
.B1(n_332),
.B2(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_64),
.A2(n_88),
.B1(n_427),
.B2(n_429),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_70),
.Y(n_314)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_70),
.Y(n_321)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_74),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g456 ( 
.A1(n_74),
.A2(n_135),
.B1(n_339),
.B2(n_457),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_74),
.A2(n_135),
.B1(n_162),
.B2(n_465),
.Y(n_464)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_74)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_76),
.Y(n_400)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_77),
.Y(n_234)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_77),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_77),
.Y(n_283)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_78),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

INVx6_ASAP7_75t_L g439 ( 
.A(n_79),
.Y(n_439)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_88),
.B(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_88),
.A2(n_332),
.B(n_338),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g308 ( 
.A1(n_91),
.A2(n_292),
.A3(n_309),
.B1(n_311),
.B2(n_315),
.Y(n_308)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_93),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_95),
.B(n_151),
.C(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_95),
.A2(n_96),
.B1(n_159),
.B2(n_160),
.Y(n_521)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_124),
.B(n_126),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_97),
.A2(n_179),
.B(n_188),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_97),
.A2(n_124),
.B1(n_233),
.B2(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_97),
.A2(n_188),
.B(n_282),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_97),
.A2(n_124),
.B1(n_398),
.B2(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_98),
.B(n_189),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_98),
.A2(n_125),
.B1(n_419),
.B2(n_423),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_98),
.A2(n_125),
.B1(n_423),
.B2(n_436),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_98),
.A2(n_125),
.B1(n_436),
.B2(n_468),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_106),
.B2(n_110),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_114),
.B1(n_118),
.B2(n_121),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_112),
.Y(n_402)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_113),
.A2(n_233),
.B(n_239),
.Y(n_232)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_116),
.Y(n_345)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_116),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_120),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_120),
.Y(n_305)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_124),
.A2(n_239),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_125),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_126),
.Y(n_468)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_129),
.Y(n_195)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_135),
.A2(n_286),
.B(n_295),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_135),
.B(n_339),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_135),
.A2(n_295),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_157),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_527)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_150),
.A2(n_151),
.B1(n_521),
.B2(n_522),
.Y(n_520)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_155),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_157),
.A2(n_158),
.B1(n_526),
.B2(n_527),
.Y(n_525)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_516),
.B(n_529),
.Y(n_170)
);

OAI311xp33_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_405),
.A3(n_492),
.B1(n_510),
.C1(n_515),
.Y(n_171)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_351),
.B(n_404),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_323),
.B(n_350),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_276),
.B(n_322),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_242),
.B(n_275),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_201),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_177),
.B(n_201),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_192),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_178),
.A2(n_192),
.B1(n_193),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_178),
.Y(n_273)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_182),
.Y(n_424)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_186),
.Y(n_310)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_186),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_187),
.A2(n_214),
.B(n_221),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g286 ( 
.A1(n_187),
.A2(n_287),
.B(n_291),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_187),
.B(n_371),
.Y(n_370)
);

OAI21xp33_ASAP7_75t_SL g387 ( 
.A1(n_187),
.A2(n_370),
.B(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_191),
.Y(n_420)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_230),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_202),
.B(n_231),
.C(n_241),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_214),
.B(n_221),
.Y(n_202)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_206),
.Y(n_413)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx4_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_214),
.A2(n_376),
.B1(n_377),
.B2(n_379),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_214),
.A2(n_411),
.B1(n_414),
.B2(n_415),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_214),
.A2(n_347),
.B(n_415),
.Y(n_440)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_215),
.B(n_224),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_215),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_215),
.A2(n_303),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_215),
.A2(n_380),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_229),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_240),
.B2(n_241),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_234),
.Y(n_422)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_266),
.B(n_274),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_254),
.B(n_265),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_253),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_252),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_252),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_264),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_260),
.B(n_263),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_263),
.A2(n_302),
.B(n_306),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_272),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_272),
.Y(n_274)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_278),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_300),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_284),
.B2(n_285),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_281),
.B(n_284),
.C(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_299),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_308),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_308),
.Y(n_329)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_324),
.B(n_325),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_330),
.B2(n_349),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_329),
.C(n_349),
.Y(n_352)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_330),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_340),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_331),
.B(n_341),
.C(n_342),
.Y(n_381)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_352),
.B(n_353),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_384),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_354)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_374),
.B2(n_375),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_357),
.B(n_374),
.Y(n_488)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_361),
.A3(n_363),
.B1(n_365),
.B2(n_370),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_381),
.B(n_382),
.C(n_384),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_386),
.B1(n_394),
.B2(n_403),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_385),
.B(n_395),
.C(n_397),
.Y(n_501)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_394),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_397),
.Y(n_394)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_478),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g510 ( 
.A1(n_406),
.A2(n_478),
.B(n_511),
.C(n_514),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_458),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_407),
.B(n_458),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_433),
.C(n_442),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g491 ( 
.A(n_408),
.B(n_433),
.CI(n_442),
.CON(n_491),
.SN(n_491)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_425),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_409),
.B(n_426),
.C(n_431),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_418),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_410),
.B(n_418),
.Y(n_484)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_419),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_431),
.Y(n_425)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_427),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_429),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_440),
.B2(n_441),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_435),
.B(n_440),
.Y(n_472)
);

INVx3_ASAP7_75t_SL g437 ( 
.A(n_438),
.Y(n_437)
);

INVx8_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_440),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_440),
.A2(n_441),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_440),
.A2(n_472),
.B(n_475),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_450),
.C(n_456),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_443),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_444),
.B(n_446),
.Y(n_500)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_450),
.A2(n_451),
.B1(n_456),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx8_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_456),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_459),
.B(n_462),
.C(n_470),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_462),
.B1(n_470),
.B2(n_471),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_466),
.B(n_469),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_467),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

FAx1_ASAP7_75t_SL g518 ( 
.A(n_469),
.B(n_519),
.CI(n_520),
.CON(n_518),
.SN(n_518)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_469),
.B(n_519),
.C(n_520),
.Y(n_528)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_491),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_479),
.B(n_491),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_484),
.C(n_485),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_480),
.A2(n_481),
.B1(n_484),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_484),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_503),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_488),
.C(n_489),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_486),
.A2(n_487),
.B1(n_489),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_489),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_491),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_493),
.B(n_505),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_494),
.A2(n_512),
.B(n_513),
.Y(n_511)
);

NOR2x1_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_502),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_502),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_499),
.C(n_501),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_508),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_499),
.A2(n_500),
.B1(n_501),
.B2(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_507),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_507),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_524),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_518),
.B(n_523),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_523),
.Y(n_530)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_518),
.Y(n_538)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_521),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_524),
.A2(n_530),
.B(n_531),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_525),
.B(n_528),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_528),
.Y(n_531)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx13_ASAP7_75t_L g535 ( 
.A(n_533),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_536),
.Y(n_534)
);


endmodule