module fake_jpeg_19304_n_324 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_11),
.B(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_27),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_34)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_25),
.A2(n_17),
.B1(n_15),
.B2(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_31),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_25),
.A2(n_16),
.B1(n_11),
.B2(n_23),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_25),
.B1(n_16),
.B2(n_18),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_11),
.B1(n_25),
.B2(n_24),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_24),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_60),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g64 ( 
.A1(n_55),
.A2(n_43),
.B1(n_34),
.B2(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_11),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_59),
.B1(n_37),
.B2(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_39),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_63),
.B(n_18),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_40),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_45),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_32),
.B(n_42),
.C(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_32),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_12),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_83),
.B(n_84),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_64),
.B(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_52),
.B1(n_60),
.B2(n_47),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_100),
.B1(n_103),
.B2(n_73),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_51),
.C(n_55),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_55),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_55),
.B1(n_48),
.B2(n_53),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_58),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_97),
.Y(n_104)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_71),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_102),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_63),
.A2(n_36),
.B1(n_37),
.B2(n_35),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g105 ( 
.A(n_86),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_80),
.B(n_72),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_113),
.B(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_81),
.B1(n_76),
.B2(n_64),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_117),
.B1(n_37),
.B2(n_36),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_78),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_111),
.B(n_22),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_122),
.B1(n_98),
.B2(n_49),
.Y(n_133)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_129),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_116),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_64),
.B1(n_77),
.B2(n_70),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_83),
.B(n_85),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_11),
.B(n_23),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_75),
.A3(n_71),
.B1(n_79),
.B2(n_26),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_26),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_79),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_120),
.Y(n_147)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_48),
.B1(n_71),
.B2(n_46),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_103),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_67),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_43),
.B(n_22),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_94),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_65),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_85),
.B1(n_100),
.B2(n_98),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_133),
.B1(n_140),
.B2(n_154),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_135),
.A2(n_157),
.B1(n_163),
.B2(n_19),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_137),
.A2(n_160),
.B(n_161),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_12),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_138),
.B(n_142),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_67),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_156),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_108),
.B1(n_109),
.B2(n_107),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_12),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_12),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_98),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_151),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_74),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_104),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_37),
.B1(n_66),
.B2(n_43),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_66),
.B1(n_43),
.B2(n_16),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_163),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_113),
.A2(n_43),
.B1(n_17),
.B2(n_18),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_74),
.B(n_23),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_128),
.A2(n_74),
.B(n_23),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_162),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_16),
.B1(n_15),
.B2(n_18),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_111),
.C(n_118),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_21),
.C(n_33),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_161),
.Y(n_214)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_121),
.B1(n_106),
.B2(n_14),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_157),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_173),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_R g172 ( 
.A(n_158),
.B(n_22),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_172),
.B(n_159),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_22),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_146),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_132),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_33),
.C(n_29),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_188),
.C(n_154),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_185),
.B1(n_138),
.B2(n_142),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_19),
.B1(n_17),
.B2(n_21),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_19),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_19),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_17),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_193),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_148),
.B1(n_143),
.B2(n_166),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_33),
.C(n_29),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_19),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_0),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_199),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_196),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_204),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_136),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_220),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_216),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_210),
.C(n_217),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_135),
.C(n_146),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_211),
.A2(n_168),
.B1(n_200),
.B2(n_174),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_162),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_218),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_221),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_144),
.B(n_150),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_150),
.C(n_144),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_12),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_213),
.B1(n_219),
.B2(n_215),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_196),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_227),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_179),
.C(n_188),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_234),
.C(n_240),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_207),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_192),
.C(n_190),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_237),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_169),
.C(n_168),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_174),
.B1(n_185),
.B2(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

AOI22x1_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_170),
.B1(n_172),
.B2(n_186),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_244),
.B1(n_240),
.B2(n_224),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_187),
.C(n_170),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_187),
.C(n_180),
.Y(n_240)
);

XOR2x2_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_26),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_225),
.B(n_233),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_29),
.C(n_33),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_218),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_204),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_254),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_238),
.B1(n_236),
.B2(n_226),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_199),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_250),
.B(n_243),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_8),
.B(n_9),
.Y(n_275)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_262),
.B1(n_8),
.B2(n_9),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_14),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_258),
.B1(n_259),
.B2(n_14),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_14),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_260),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_14),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_238),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_230),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_246),
.B(n_229),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_271),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_260),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_267),
.A2(n_250),
.B1(n_256),
.B2(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_28),
.C(n_31),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_33),
.C(n_29),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_261),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_274),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_275),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_28),
.B1(n_30),
.B2(n_10),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_8),
.B1(n_9),
.B2(n_7),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_6),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_8),
.B1(n_7),
.B2(n_6),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_287),
.B1(n_289),
.B2(n_4),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_280),
.B(n_13),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_262),
.B(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_285),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_257),
.B(n_7),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_14),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_33),
.B1(n_29),
.B2(n_13),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_6),
.B(n_2),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_268),
.B(n_3),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_291),
.A2(n_270),
.B1(n_268),
.B2(n_263),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_292),
.B(n_297),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_29),
.C(n_33),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_300),
.C(n_303),
.Y(n_306)
);

AOI321xp33_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_14),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_1),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_301),
.B(n_302),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_1),
.B(n_3),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_279),
.B(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_29),
.C(n_13),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_14),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_295),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_308),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_298),
.A2(n_283),
.B(n_286),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_312),
.B(n_300),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_13),
.C(n_20),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_297),
.Y(n_312)
);

OAI321xp33_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_312),
.A3(n_304),
.B1(n_311),
.B2(n_306),
.C(n_5),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_20),
.B(n_5),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

OAI321xp33_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_20),
.A3(n_315),
.B1(n_316),
.B2(n_298),
.C(n_296),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_20),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_320),
.B(n_20),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_20),
.B(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_20),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_20),
.B(n_45),
.Y(n_324)
);


endmodule