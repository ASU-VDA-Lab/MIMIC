module real_jpeg_1293_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_1),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_1),
.A2(n_37),
.B1(n_39),
.B2(n_93),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_93),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_93),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_2),
.B(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_2),
.B(n_42),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_2),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_2),
.A2(n_30),
.B(n_81),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_2),
.B(n_48),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_2),
.A2(n_39),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_2),
.B(n_62),
.C(n_65),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_149),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_2),
.B(n_75),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_2),
.B(n_104),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_77),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_5),
.A2(n_37),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_45),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_5),
.A2(n_45),
.B1(n_65),
.B2(n_66),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_71),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_11),
.A2(n_27),
.B1(n_37),
.B2(n_39),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_11),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_11),
.A2(n_27),
.B1(n_65),
.B2(n_66),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_12),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_12),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_12),
.A2(n_41),
.B1(n_65),
.B2(n_66),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_13),
.A2(n_37),
.B1(n_39),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_55),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_13),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_14),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_15),
.A2(n_37),
.B1(n_39),
.B2(n_68),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_127),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_106),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_22),
.B(n_106),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_78),
.C(n_95),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_23),
.B(n_95),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_56),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_43),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_25),
.B(n_43),
.C(n_56),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_40),
.B2(n_42),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_28),
.A2(n_35),
.A3(n_39),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_33),
.B(n_37),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_36),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_36),
.A2(n_91),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_36),
.A2(n_91),
.B1(n_92),
.B2(n_161),
.Y(n_160)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_39),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_37),
.B(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_39),
.A2(n_50),
.A3(n_51),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_54),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_47),
.A2(n_88),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_47),
.A2(n_88),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_47),
.A2(n_87),
.B1(n_88),
.B2(n_135),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_47),
.A2(n_88),
.B1(n_134),
.B2(n_182),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_49),
.B(n_52),
.Y(n_150)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_50),
.B(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_69),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_57),
.B(n_69),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_64),
.B2(n_67),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_59),
.A2(n_64),
.B1(n_144),
.B2(n_185),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_103),
.B1(n_104),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_60),
.A2(n_104),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_60),
.A2(n_104),
.B1(n_145),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_60),
.A2(n_104),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_60),
.A2(n_104),
.B1(n_173),
.B2(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_65),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_65),
.B(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_74),
.B(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_72),
.A2(n_74),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_72),
.A2(n_74),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_75),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_75),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_73),
.A2(n_75),
.B1(n_84),
.B2(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_73),
.A2(n_75),
.B1(n_153),
.B2(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_73),
.A2(n_75),
.B1(n_149),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_73),
.A2(n_75),
.B1(n_203),
.B2(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_78),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_86),
.C(n_90),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_79),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_80),
.B(n_83),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_86),
.B(n_90),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_105),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_105),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_116),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_125),
.B2(n_126),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

AOI31xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_223),
.A3(n_232),
.B(n_236),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_168),
.B(n_222),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_155),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_131),
.B(n_155),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_142),
.C(n_146),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_132),
.B(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_137),
.C(n_141),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_141),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_142),
.B(n_146),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_157),
.B(n_158),
.C(n_159),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_160),
.B(n_163),
.C(n_167),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_164),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_217),
.B(n_221),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_186),
.B(n_216),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_178),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_175),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_181),
.C(n_184),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_197),
.B(n_215),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_195),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_209),
.B(n_214),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_204),
.B(n_208),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_206),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_213),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_220),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.C(n_231),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_231),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_234),
.Y(n_237)
);


endmodule