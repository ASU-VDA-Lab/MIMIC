module real_jpeg_31420_n_23 (n_17, n_8, n_0, n_21, n_168, n_2, n_10, n_175, n_9, n_12, n_166, n_170, n_6, n_176, n_171, n_169, n_167, n_177, n_11, n_14, n_172, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_1, n_20, n_19, n_16, n_15, n_13, n_23);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_10;
input n_175;
input n_9;
input n_12;
input n_166;
input n_170;
input n_6;
input n_176;
input n_171;
input n_169;
input n_167;
input n_177;
input n_11;
input n_14;
input n_172;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_23;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_0),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_1),
.B(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_2),
.B(n_98),
.Y(n_97)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_2),
.B(n_98),
.CON(n_110),
.SN(n_110)
);

AOI221xp5_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_17),
.B1(n_47),
.B2(n_51),
.C(n_55),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_47),
.C(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_8),
.B(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_8),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_9),
.B(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_12),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_13),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_14),
.B(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_14),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_15),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_15),
.B(n_144),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_16),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_16),
.B(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_19),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_20),
.A2(n_79),
.A3(n_81),
.B1(n_88),
.B2(n_113),
.C1(n_115),
.C2(n_176),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_21),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_21),
.B(n_121),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_22),
.B(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_R g49 ( 
.A(n_31),
.B(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_125),
.B(n_148),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_118),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI31xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_72),
.A3(n_102),
.B(n_108),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_66),
.C(n_67),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_59),
.B(n_65),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_51),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_168),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_63),
.Y(n_71)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_87),
.C(n_97),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_109),
.B(n_112),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_97),
.C(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_172),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

OA21x2_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_96),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_110),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_134),
.C(n_138),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_159),
.C(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI322xp33_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_140),
.A3(n_158),
.B1(n_161),
.B2(n_162),
.C1(n_163),
.C2(n_177),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_149),
.B(n_156),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVxp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_166),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_167),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_169),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_170),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_171),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_173),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_174),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_175),
.Y(n_105)
);


endmodule