module fake_jpeg_22900_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx8_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_40),
.Y(n_42)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_16),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_51),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_26),
.B1(n_16),
.B2(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_58),
.B1(n_32),
.B2(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_26),
.B1(n_28),
.B2(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_62),
.Y(n_79)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_68),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_80),
.B1(n_35),
.B2(n_32),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_78),
.Y(n_90)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_42),
.B(n_40),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_25),
.B1(n_23),
.B2(n_15),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_33),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_17),
.B1(n_21),
.B2(n_22),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_111),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_55),
.C(n_31),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_106),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_57),
.B(n_54),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_102),
.B(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_100),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_68),
.B1(n_35),
.B2(n_71),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_50),
.B(n_25),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_31),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_31),
.C(n_33),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_70),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_35),
.B1(n_39),
.B2(n_38),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_82),
.B1(n_72),
.B2(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_21),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_78),
.Y(n_126)
);

BUFx8_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_115),
.B1(n_137),
.B2(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_112),
.A2(n_70),
.B1(n_68),
.B2(n_74),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_121),
.B1(n_134),
.B2(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_119),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_124),
.B(n_92),
.Y(n_142)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_70),
.B1(n_81),
.B2(n_76),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_76),
.B1(n_82),
.B2(n_23),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_123),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_63),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_132),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_85),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_22),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_38),
.B1(n_77),
.B2(n_72),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_106),
.C(n_102),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_82),
.B1(n_77),
.B2(n_38),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_132),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_95),
.B1(n_131),
.B2(n_135),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_158),
.B(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_155),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_127),
.A2(n_28),
.B(n_22),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_154),
.B(n_130),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_107),
.B1(n_88),
.B2(n_96),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_151),
.B1(n_153),
.B2(n_163),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_107),
.B1(n_88),
.B2(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_161),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_56),
.B1(n_62),
.B2(n_46),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_15),
.B(n_23),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_111),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_129),
.A2(n_104),
.B(n_25),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_128),
.B(n_15),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_116),
.B(n_117),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_134),
.A3(n_114),
.B1(n_137),
.B2(n_115),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_122),
.A2(n_79),
.B(n_45),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_126),
.A2(n_87),
.B1(n_104),
.B2(n_65),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_175),
.B(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_182),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_135),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_187),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_172),
.A2(n_60),
.B1(n_30),
.B2(n_29),
.Y(n_213)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_183),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_75),
.C(n_65),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_185),
.C(n_162),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_75),
.B(n_120),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_159),
.B(n_20),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_186),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_133),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_188),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_37),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_133),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_37),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_89),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_139),
.A2(n_164),
.B(n_154),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_29),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_171),
.B(n_153),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_206),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_208),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_185),
.C(n_168),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_165),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_189),
.A2(n_145),
.B1(n_139),
.B2(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_143),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_133),
.B1(n_24),
.B2(n_27),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_27),
.B1(n_24),
.B2(n_30),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_64),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_18),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_213),
.B(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_64),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_197),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_222),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_225),
.C(n_204),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_179),
.B1(n_175),
.B2(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_188),
.C(n_190),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_187),
.C(n_166),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_170),
.B(n_181),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_230),
.B(n_193),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_183),
.B1(n_165),
.B2(n_177),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_235),
.B1(n_203),
.B2(n_209),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_206),
.A2(n_177),
.B(n_27),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_208),
.Y(n_232)
);

INVxp33_ASAP7_75t_SL g247 ( 
.A(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_0),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_194),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_192),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_246),
.B1(n_250),
.B2(n_234),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_204),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_253),
.C(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_243),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_232),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_215),
.B1(n_227),
.B2(n_216),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_196),
.B1(n_205),
.B2(n_198),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_201),
.CI(n_200),
.CON(n_249),
.SN(n_249)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_249),
.B(n_226),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_198),
.B1(n_214),
.B2(n_194),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_210),
.C(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_264),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_215),
.C(n_216),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_263),
.C(n_265),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_111),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_231),
.C(n_218),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_236),
.B(n_251),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_230),
.B(n_195),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_237),
.A2(n_203),
.B1(n_233),
.B2(n_211),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_270),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_269),
.A2(n_242),
.B1(n_249),
.B2(n_243),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_240),
.C(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_281),
.C(n_282),
.Y(n_286)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_0),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_254),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_280),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_279),
.A2(n_283),
.B1(n_256),
.B2(n_268),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_111),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_67),
.C(n_24),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_67),
.B1(n_30),
.B2(n_18),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_60),
.C(n_10),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_8),
.C(n_14),
.Y(n_291)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_263),
.C(n_258),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_294),
.C(n_14),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_291),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_275),
.A2(n_8),
.B1(n_11),
.B2(n_7),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_289),
.B(n_292),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_278),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_18),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_11),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_278),
.B(n_276),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_293),
.A2(n_295),
.B(n_6),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_18),
.C(n_30),
.Y(n_294)
);

NOR2x1_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_6),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_297),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_41),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_41),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_290),
.A3(n_295),
.B1(n_6),
.B2(n_12),
.C1(n_13),
.C2(n_5),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_304),
.A2(n_305),
.B(n_298),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_13),
.B(n_12),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_308),
.B(n_311),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_303),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_309)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g313 ( 
.A1(n_309),
.A2(n_300),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_41),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_313),
.C(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_314),
.C(n_310),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_3),
.B(n_4),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_4),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_41),
.Y(n_320)
);


endmodule