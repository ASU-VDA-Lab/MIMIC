module fake_aes_6321_n_716 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_716);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_716;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_564;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g81 ( .A(n_6), .Y(n_81) );
INVxp67_ASAP7_75t_L g82 ( .A(n_35), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_5), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_6), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_74), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_19), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_61), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_39), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_62), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_40), .Y(n_90) );
INVx1_ASAP7_75t_SL g91 ( .A(n_9), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_41), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_69), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_44), .Y(n_96) );
BUFx2_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_72), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_26), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_77), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_66), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_80), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_43), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_78), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_64), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_15), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_23), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_52), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_30), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_37), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_49), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_25), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_20), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_32), .Y(n_116) );
CKINVDCx14_ASAP7_75t_R g117 ( .A(n_50), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_59), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_71), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_12), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_58), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_9), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_63), .B(n_65), .Y(n_123) );
INVxp33_ASAP7_75t_SL g124 ( .A(n_47), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_3), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_68), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_23), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_28), .Y(n_128) );
INVxp33_ASAP7_75t_L g129 ( .A(n_76), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_54), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_97), .B(n_0), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_97), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_125), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_125), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_116), .B(n_1), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_106), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_117), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_125), .B(n_1), .Y(n_139) );
NOR2xp33_ASAP7_75t_R g140 ( .A(n_108), .B(n_29), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_127), .B(n_4), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_119), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_127), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_129), .B(n_4), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_106), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
NAND2xp33_ASAP7_75t_R g148 ( .A(n_124), .B(n_31), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_83), .B(n_5), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_83), .B(n_7), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_87), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_82), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_91), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
CKINVDCx8_ASAP7_75t_R g155 ( .A(n_81), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_88), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
XNOR2xp5_ASAP7_75t_L g158 ( .A(n_91), .B(n_7), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_114), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_85), .B(n_34), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_81), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_90), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_81), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_114), .B(n_8), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_98), .Y(n_166) );
NAND2xp33_ASAP7_75t_L g167 ( .A(n_85), .B(n_79), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_81), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_89), .Y(n_169) );
INVxp67_ASAP7_75t_SL g170 ( .A(n_86), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_99), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_111), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_81), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_86), .Y(n_174) );
NOR2xp67_ASAP7_75t_L g175 ( .A(n_92), .B(n_8), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_131), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_168), .Y(n_177) );
AND2x2_ASAP7_75t_L g178 ( .A(n_137), .B(n_110), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_159), .B(n_130), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_169), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_169), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_168), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_152), .B(n_151), .Y(n_186) );
AND2x6_ASAP7_75t_L g187 ( .A(n_139), .B(n_130), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_168), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_169), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_139), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_170), .B(n_107), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_138), .B(n_105), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_145), .Y(n_196) );
INVx5_ASAP7_75t_L g197 ( .A(n_160), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_151), .B(n_105), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
OR2x2_ASAP7_75t_L g200 ( .A(n_146), .B(n_93), .Y(n_200) );
INVx8_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_145), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_141), .Y(n_204) );
OAI22xp33_ASAP7_75t_SL g205 ( .A1(n_133), .A2(n_107), .B1(n_93), .B2(n_110), .Y(n_205) );
AND2x6_ASAP7_75t_L g206 ( .A(n_141), .B(n_109), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_141), .Y(n_208) );
INVxp67_ASAP7_75t_L g209 ( .A(n_132), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_132), .A2(n_84), .B1(n_113), .B2(n_115), .Y(n_210) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_174), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_160), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_143), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_134), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_142), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_143), .Y(n_216) );
AO22x2_ASAP7_75t_L g217 ( .A1(n_154), .A2(n_104), .B1(n_92), .B2(n_96), .Y(n_217) );
OR2x2_ASAP7_75t_L g218 ( .A(n_136), .B(n_122), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_134), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_154), .B(n_113), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_166), .B(n_109), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_135), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_135), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_144), .Y(n_225) );
BUFx8_ASAP7_75t_SL g226 ( .A(n_171), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_149), .A2(n_115), .B1(n_120), .B2(n_122), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_156), .B(n_120), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_144), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_147), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_156), .B(n_103), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_157), .B(n_103), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_161), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_160), .Y(n_235) );
INVx5_ASAP7_75t_L g236 ( .A(n_160), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_160), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_157), .B(n_102), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_160), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_162), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_162), .B(n_102), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_165), .B(n_104), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_196), .B(n_172), .Y(n_243) );
NOR2xp33_ASAP7_75t_R g244 ( .A(n_215), .B(n_163), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_208), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_234), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_193), .B(n_150), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_186), .B(n_164), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_214), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_184), .B(n_165), .Y(n_250) );
BUFx10_ASAP7_75t_L g251 ( .A(n_187), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_196), .B(n_149), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_214), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_187), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_208), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_202), .B(n_150), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
BUFx12f_ASAP7_75t_SL g258 ( .A(n_178), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_209), .A2(n_173), .B1(n_148), .B2(n_175), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_184), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_189), .Y(n_261) );
AOI22x1_ASAP7_75t_L g262 ( .A1(n_235), .A2(n_89), .B1(n_126), .B2(n_128), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_187), .A2(n_175), .B1(n_167), .B2(n_158), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_189), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_193), .B(n_140), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_193), .B(n_101), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_178), .B(n_158), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_229), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_219), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_208), .Y(n_270) );
INVxp67_ASAP7_75t_L g271 ( .A(n_211), .Y(n_271) );
NOR3xp33_ASAP7_75t_SL g272 ( .A(n_194), .B(n_112), .C(n_95), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_193), .B(n_101), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_221), .B(n_100), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_229), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_208), .B(n_118), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_200), .Y(n_277) );
BUFx2_ASAP7_75t_SL g278 ( .A(n_187), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_184), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_205), .A2(n_118), .B(n_94), .C(n_95), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_200), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_218), .B(n_100), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_187), .A2(n_121), .B1(n_94), .B2(n_96), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_218), .B(n_221), .Y(n_285) );
NOR3xp33_ASAP7_75t_SL g286 ( .A(n_222), .B(n_121), .C(n_123), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_181), .B(n_155), .Y(n_287) );
NOR2xp33_ASAP7_75t_R g288 ( .A(n_201), .B(n_155), .Y(n_288) );
AOI211xp5_ASAP7_75t_L g289 ( .A1(n_205), .A2(n_128), .B(n_126), .C(n_89), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_237), .A2(n_239), .B(n_235), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_238), .B(n_187), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_223), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_184), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_187), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_238), .B(n_128), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_228), .B(n_126), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_224), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_228), .B(n_10), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_238), .B(n_10), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_238), .B(n_11), .Y(n_300) );
NOR2xp33_ASAP7_75t_R g301 ( .A(n_201), .B(n_11), .Y(n_301) );
NAND3xp33_ASAP7_75t_SL g302 ( .A(n_210), .B(n_12), .C(n_13), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_206), .B(n_13), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_229), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_226), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_217), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_217), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_206), .B(n_14), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_224), .Y(n_309) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_184), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_206), .B(n_15), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_206), .B(n_16), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_191), .B(n_42), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_217), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_251), .Y(n_315) );
CKINVDCx11_ASAP7_75t_R g316 ( .A(n_246), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_249), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_299), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_253), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_268), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_257), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_269), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_291), .A2(n_207), .B(n_199), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_285), .B(n_206), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_247), .B(n_207), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_254), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_279), .Y(n_327) );
AOI21xp33_ASAP7_75t_L g328 ( .A1(n_277), .A2(n_191), .B(n_192), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_299), .A2(n_206), .B1(n_210), .B2(n_204), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_265), .A2(n_204), .B(n_192), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_247), .B(n_199), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_248), .B(n_206), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_248), .B(n_240), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_245), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_282), .B(n_227), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_268), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_245), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_299), .Y(n_338) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_254), .Y(n_339) );
OR2x6_ASAP7_75t_L g340 ( .A(n_278), .B(n_201), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_247), .B(n_217), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_283), .B(n_240), .Y(n_343) );
INVx3_ASAP7_75t_SL g344 ( .A(n_246), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_275), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_294), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_258), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_294), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_306), .A2(n_242), .B1(n_241), .B2(n_198), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_243), .A2(n_231), .B1(n_232), .B2(n_201), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_L g351 ( .A1(n_281), .A2(n_225), .B(n_233), .C(n_179), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_297), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_251), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_275), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_298), .B(n_239), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_244), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_251), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_266), .B(n_225), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_260), .Y(n_360) );
INVx5_ASAP7_75t_L g361 ( .A(n_304), .Y(n_361) );
O2A1O1Ixp33_ASAP7_75t_L g362 ( .A1(n_307), .A2(n_233), .B(n_179), .C(n_176), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_258), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_309), .A2(n_201), .B(n_239), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_304), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_314), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_250), .A2(n_239), .B(n_237), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_245), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_255), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_255), .Y(n_370) );
OA21x2_ASAP7_75t_L g371 ( .A1(n_317), .A2(n_290), .B(n_262), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_318), .A2(n_298), .B1(n_276), .B2(n_266), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_335), .A2(n_267), .B1(n_264), .B2(n_271), .C(n_252), .Y(n_374) );
OR2x4_ASAP7_75t_L g375 ( .A(n_333), .B(n_302), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_361), .Y(n_376) );
AND2x2_ASAP7_75t_SL g377 ( .A(n_318), .B(n_298), .Y(n_377) );
INVx4_ASAP7_75t_SL g378 ( .A(n_340), .Y(n_378) );
CKINVDCx6p67_ASAP7_75t_R g379 ( .A(n_344), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_319), .Y(n_380) );
CKINVDCx6p67_ASAP7_75t_R g381 ( .A(n_344), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_338), .A2(n_276), .B1(n_266), .B2(n_284), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_320), .Y(n_383) );
NAND3xp33_ASAP7_75t_SL g384 ( .A(n_357), .B(n_244), .C(n_261), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_338), .A2(n_263), .B1(n_259), .B2(n_256), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_329), .A2(n_274), .B1(n_273), .B2(n_300), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_319), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_321), .Y(n_389) );
OA21x2_ASAP7_75t_L g390 ( .A1(n_321), .A2(n_290), .B(n_313), .Y(n_390) );
AO31x2_ASAP7_75t_L g391 ( .A1(n_349), .A2(n_313), .A3(n_295), .B(n_230), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_322), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_343), .A2(n_274), .B1(n_296), .B2(n_289), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_322), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_361), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_341), .A2(n_274), .B1(n_296), .B2(n_255), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_326), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_347), .B(n_305), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_357), .A2(n_301), .B1(n_296), .B2(n_303), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_341), .A2(n_270), .B1(n_287), .B2(n_301), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_324), .A2(n_312), .B1(n_311), .B2(n_308), .Y(n_401) );
AND2x6_ASAP7_75t_L g402 ( .A(n_326), .B(n_270), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_347), .A2(n_363), .B1(n_366), .B2(n_331), .Y(n_403) );
OA21x2_ASAP7_75t_L g404 ( .A1(n_327), .A2(n_286), .B(n_176), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_327), .Y(n_405) );
OAI21x1_ASAP7_75t_SL g406 ( .A1(n_373), .A2(n_362), .B(n_352), .Y(n_406) );
AOI222xp33_ASAP7_75t_L g407 ( .A1(n_374), .A2(n_316), .B1(n_352), .B2(n_342), .C1(n_363), .C2(n_331), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_377), .B(n_342), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_380), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_402), .Y(n_411) );
OAI31xp33_ASAP7_75t_SL g412 ( .A1(n_393), .A2(n_328), .A3(n_331), .B(n_325), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_377), .A2(n_350), .B1(n_359), .B2(n_332), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_387), .A2(n_325), .B1(n_355), .B2(n_330), .Y(n_414) );
NAND2xp33_ASAP7_75t_L g415 ( .A(n_402), .B(n_326), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_382), .A2(n_325), .B1(n_320), .B2(n_336), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_404), .A2(n_316), .B1(n_355), .B2(n_287), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_402), .Y(n_418) );
AOI322xp5_ASAP7_75t_L g419 ( .A1(n_384), .A2(n_272), .A3(n_230), .B1(n_183), .B2(n_190), .C1(n_182), .C2(n_180), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_404), .A2(n_355), .B1(n_368), .B2(n_369), .Y(n_420) );
A2O1A1Ixp33_ASAP7_75t_L g421 ( .A1(n_385), .A2(n_351), .B(n_323), .C(n_365), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_404), .A2(n_368), .B1(n_334), .B2(n_337), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_379), .A2(n_368), .B1(n_365), .B2(n_370), .Y(n_423) );
AO21x2_ASAP7_75t_L g424 ( .A1(n_401), .A2(n_364), .B(n_345), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_379), .A2(n_365), .B1(n_370), .B2(n_270), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_396), .A2(n_354), .B1(n_345), .B2(n_336), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_380), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_381), .A2(n_361), .B1(n_356), .B2(n_346), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_381), .A2(n_361), .B1(n_356), .B2(n_346), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_375), .A2(n_354), .B1(n_180), .B2(n_190), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_405), .B(n_361), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_405), .B(n_183), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_375), .A2(n_340), .B1(n_182), .B2(n_348), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_372), .B(n_326), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_398), .A2(n_250), .B1(n_237), .B2(n_367), .C(n_212), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_408), .B(n_383), .Y(n_436) );
AND2x4_ASAP7_75t_L g437 ( .A(n_418), .B(n_378), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_416), .A2(n_375), .B1(n_388), .B2(n_392), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_410), .B(n_389), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_408), .B(n_394), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_409), .B(n_403), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_408), .B(n_391), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_416), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_427), .B(n_386), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_427), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_434), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_432), .Y(n_448) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_406), .A2(n_391), .B(n_390), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_409), .B(n_386), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_413), .A2(n_400), .B1(n_399), .B2(n_395), .C(n_376), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_432), .Y(n_452) );
NOR4xp25_ASAP7_75t_SL g453 ( .A(n_421), .B(n_378), .C(n_391), .D(n_402), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_411), .Y(n_454) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_422), .A2(n_391), .B(n_390), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_434), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_407), .A2(n_378), .B1(n_376), .B2(n_395), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_430), .B(n_391), .Y(n_458) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_407), .A2(n_397), .B(n_288), .C(n_371), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_424), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_431), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_406), .A2(n_237), .B1(n_397), .B2(n_212), .C(n_348), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_418), .Y(n_464) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_433), .A2(n_378), .B1(n_402), .B2(n_397), .C1(n_212), .C2(n_20), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_411), .Y(n_466) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_430), .A2(n_390), .B(n_371), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_412), .B(n_371), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_414), .A2(n_340), .B1(n_326), .B2(n_339), .Y(n_469) );
NAND2xp33_ASAP7_75t_R g470 ( .A(n_418), .B(n_288), .Y(n_470) );
AO21x2_ASAP7_75t_L g471 ( .A1(n_424), .A2(n_216), .B(n_203), .Y(n_471) );
NOR4xp25_ASAP7_75t_SL g472 ( .A(n_412), .B(n_402), .C(n_17), .D(n_18), .Y(n_472) );
AOI221xp5_ASAP7_75t_SL g473 ( .A1(n_438), .A2(n_417), .B1(n_433), .B2(n_420), .C(n_423), .Y(n_473) );
AOI221xp5_ASAP7_75t_L g474 ( .A1(n_438), .A2(n_426), .B1(n_425), .B2(n_414), .C(n_429), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_462), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_451), .A2(n_424), .B1(n_411), .B2(n_428), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_447), .B(n_418), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_462), .B(n_424), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_447), .B(n_16), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_451), .A2(n_435), .B1(n_415), .B2(n_419), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_443), .A2(n_339), .B1(n_419), .B2(n_340), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_447), .B(n_17), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_448), .B(n_18), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_448), .B(n_19), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_456), .B(n_21), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_452), .B(n_21), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_456), .B(n_22), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_456), .B(n_22), .Y(n_489) );
OR2x6_ASAP7_75t_L g490 ( .A(n_443), .B(n_339), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_444), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_444), .B(n_24), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
INVx4_ASAP7_75t_SL g494 ( .A(n_437), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_437), .B(n_51), .Y(n_495) );
NOR2x1_ASAP7_75t_L g496 ( .A(n_459), .B(n_339), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_459), .A2(n_24), .A3(n_358), .B(n_315), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_442), .B(n_27), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_442), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_439), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_436), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_439), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_436), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_445), .Y(n_505) );
INVx4_ASAP7_75t_L g506 ( .A(n_437), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_440), .Y(n_507) );
INVx4_ASAP7_75t_L g508 ( .A(n_437), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_457), .A2(n_212), .B1(n_339), .B2(n_236), .C(n_197), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_458), .B(n_450), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_458), .B(n_33), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_450), .B(n_36), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_442), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_436), .B(n_38), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_440), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_440), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_452), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_461), .B(n_45), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_464), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_461), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_437), .B(n_46), .Y(n_521) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_441), .A2(n_203), .B1(n_213), .B2(n_216), .C(n_220), .Y(n_522) );
INVx1_ASAP7_75t_SL g523 ( .A(n_466), .Y(n_523) );
AND2x4_ASAP7_75t_SL g524 ( .A(n_506), .B(n_464), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_501), .B(n_465), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_503), .B(n_465), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_505), .B(n_468), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_493), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_500), .B(n_468), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_498), .A2(n_469), .B(n_453), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_506), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_506), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_493), .Y(n_533) );
NOR2xp33_ASAP7_75t_R g534 ( .A(n_500), .B(n_470), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_507), .B(n_468), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_520), .B(n_449), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_483), .B(n_466), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_484), .Y(n_538) );
INVx6_ASAP7_75t_L g539 ( .A(n_494), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_475), .Y(n_540) );
NOR3xp33_ASAP7_75t_SL g541 ( .A(n_485), .B(n_487), .C(n_474), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_513), .B(n_449), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_517), .B(n_449), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_497), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_523), .Y(n_545) );
OAI21xp33_ASAP7_75t_L g546 ( .A1(n_476), .A2(n_460), .B(n_463), .Y(n_546) );
INVxp67_ASAP7_75t_SL g547 ( .A(n_492), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_513), .B(n_449), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_494), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_515), .B(n_460), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_502), .B(n_455), .Y(n_552) );
OAI211xp5_ASAP7_75t_L g553 ( .A1(n_473), .A2(n_472), .B(n_453), .C(n_463), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_508), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_515), .B(n_460), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_510), .B(n_455), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_502), .B(n_455), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_491), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_516), .B(n_455), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_516), .B(n_455), .Y(n_561) );
NAND2xp33_ASAP7_75t_SL g562 ( .A(n_508), .B(n_469), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_479), .Y(n_563) );
NAND5xp2_ASAP7_75t_SL g564 ( .A(n_481), .B(n_467), .C(n_472), .D(n_454), .E(n_471), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_510), .B(n_454), .Y(n_565) );
OAI31xp33_ASAP7_75t_L g566 ( .A1(n_495), .A2(n_454), .A3(n_358), .B(n_315), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_495), .B(n_467), .Y(n_567) );
NAND2xp33_ASAP7_75t_R g568 ( .A(n_495), .B(n_48), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_491), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_504), .B(n_471), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_478), .B(n_471), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_492), .Y(n_572) );
OAI21xp5_ASAP7_75t_L g573 ( .A1(n_480), .A2(n_197), .B(n_236), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_504), .B(n_471), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_479), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_519), .Y(n_576) );
INVxp33_ASAP7_75t_L g577 ( .A(n_521), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_519), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_478), .B(n_53), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_482), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_477), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_508), .B(n_55), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_528), .Y(n_583) );
NOR3xp33_ASAP7_75t_L g584 ( .A(n_553), .B(n_488), .C(n_489), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_528), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_533), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_533), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_568), .A2(n_521), .B1(n_488), .B2(n_489), .Y(n_588) );
AOI32xp33_ASAP7_75t_L g589 ( .A1(n_562), .A2(n_496), .A3(n_521), .B1(n_499), .B2(n_486), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_540), .B(n_486), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_576), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_576), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_578), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_545), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_578), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_558), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_538), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_532), .A2(n_512), .B1(n_518), .B2(n_511), .Y(n_598) );
NAND3xp33_ASAP7_75t_SL g599 ( .A(n_566), .B(n_512), .C(n_518), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_529), .B(n_477), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_529), .B(n_514), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_527), .B(n_490), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_558), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_554), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_569), .Y(n_605) );
AOI21x1_ASAP7_75t_L g606 ( .A1(n_582), .A2(n_514), .B(n_490), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_569), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_544), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_563), .B(n_494), .Y(n_609) );
OAI22xp33_ASAP7_75t_SL g610 ( .A1(n_539), .A2(n_490), .B1(n_494), .B2(n_509), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_575), .B(n_490), .Y(n_611) );
AND2x2_ASAP7_75t_SL g612 ( .A(n_554), .B(n_522), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_580), .B(n_56), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_544), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_542), .B(n_57), .Y(n_615) );
OAI31xp33_ASAP7_75t_L g616 ( .A1(n_562), .A2(n_358), .A3(n_315), .B(n_73), .Y(n_616) );
OAI32xp33_ASAP7_75t_L g617 ( .A1(n_577), .A2(n_67), .A3(n_70), .B1(n_75), .B2(n_213), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g618 ( .A1(n_525), .A2(n_220), .B1(n_185), .B2(n_188), .C(n_195), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_564), .A2(n_212), .B1(n_360), .B2(n_236), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_581), .B(n_360), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_541), .A2(n_360), .B1(n_236), .B2(n_197), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_526), .A2(n_177), .B1(n_185), .B2(n_188), .C(n_195), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_530), .A2(n_360), .B(n_353), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_551), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_549), .A2(n_353), .B1(n_197), .B2(n_236), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_542), .B(n_177), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_581), .B(n_260), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_564), .A2(n_197), .B1(n_260), .B2(n_280), .C(n_293), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_535), .B(n_353), .Y(n_629) );
NOR3xp33_ASAP7_75t_SL g630 ( .A(n_537), .B(n_353), .C(n_280), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_548), .B(n_260), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_538), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_548), .B(n_280), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_583), .Y(n_634) );
NOR4xp25_ASAP7_75t_SL g635 ( .A(n_618), .B(n_567), .C(n_546), .D(n_547), .Y(n_635) );
NOR3xp33_ASAP7_75t_SL g636 ( .A(n_599), .B(n_565), .C(n_543), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_600), .B(n_552), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_585), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_586), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_597), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g641 ( .A(n_618), .B(n_582), .C(n_579), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_604), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_604), .Y(n_643) );
AND3x2_ASAP7_75t_L g644 ( .A(n_584), .B(n_572), .C(n_579), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_587), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_596), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g647 ( .A(n_594), .B(n_536), .C(n_573), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_590), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_603), .B(n_556), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_605), .B(n_552), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_607), .B(n_557), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_632), .B(n_557), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_591), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_608), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_588), .A2(n_539), .B1(n_531), .B2(n_571), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_612), .B(n_539), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_609), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_611), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_592), .B(n_570), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_624), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_593), .B(n_570), .Y(n_662) );
OAI221xp5_ASAP7_75t_SL g663 ( .A1(n_589), .A2(n_571), .B1(n_531), .B2(n_561), .C(n_560), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_610), .B(n_534), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_613), .B(n_574), .C(n_555), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_595), .Y(n_666) );
INVx1_ASAP7_75t_SL g667 ( .A(n_602), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_599), .A2(n_550), .B(n_551), .Y(n_668) );
AOI22xp33_ASAP7_75t_R g669 ( .A1(n_616), .A2(n_559), .B1(n_524), .B2(n_310), .Y(n_669) );
XNOR2xp5_ASAP7_75t_L g670 ( .A(n_664), .B(n_601), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_640), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_634), .Y(n_672) );
OAI322xp33_ASAP7_75t_L g673 ( .A1(n_664), .A2(n_626), .A3(n_598), .B1(n_623), .B2(n_615), .C1(n_629), .C2(n_621), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g674 ( .A1(n_668), .A2(n_630), .B(n_606), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_637), .B(n_633), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_667), .B(n_620), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_663), .A2(n_622), .B1(n_617), .B2(n_628), .C(n_631), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_636), .B(n_628), .Y(n_678) );
XOR2x2_ASAP7_75t_L g679 ( .A(n_644), .B(n_622), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_657), .A2(n_627), .B(n_619), .C(n_625), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_648), .B(n_293), .Y(n_681) );
NOR2x1_ASAP7_75t_L g682 ( .A(n_643), .B(n_310), .Y(n_682) );
INVx2_ASAP7_75t_SL g683 ( .A(n_658), .Y(n_683) );
OAI32xp33_ASAP7_75t_L g684 ( .A1(n_641), .A2(n_310), .A3(n_642), .B1(n_658), .B2(n_659), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_643), .Y(n_685) );
NOR2x1p5_ASAP7_75t_L g686 ( .A(n_649), .B(n_651), .Y(n_686) );
A2O1A1Ixp33_ASAP7_75t_L g687 ( .A1(n_647), .A2(n_669), .B(n_665), .C(n_635), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_678), .A2(n_655), .B(n_654), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_679), .A2(n_662), .B1(n_660), .B2(n_652), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_685), .Y(n_690) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_683), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_687), .A2(n_638), .B1(n_645), .B2(n_646), .C(n_661), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g693 ( .A(n_670), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_687), .B(n_656), .C(n_639), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_684), .A2(n_650), .B1(n_639), .B2(n_653), .C(n_666), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_686), .B(n_666), .Y(n_696) );
AO22x2_ASAP7_75t_L g697 ( .A1(n_685), .A2(n_640), .B1(n_678), .B2(n_674), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_675), .B(n_672), .Y(n_698) );
AOI322xp5_ASAP7_75t_L g699 ( .A1(n_676), .A2(n_680), .A3(n_677), .B1(n_671), .B2(n_679), .C1(n_682), .C2(n_681), .Y(n_699) );
OAI21xp5_ASAP7_75t_SL g700 ( .A1(n_680), .A2(n_681), .B(n_673), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_L g701 ( .A1(n_687), .A2(n_678), .B(n_684), .C(n_664), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_679), .A2(n_678), .B1(n_670), .B2(n_664), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_690), .Y(n_703) );
OAI211xp5_ASAP7_75t_SL g704 ( .A1(n_701), .A2(n_699), .B(n_702), .C(n_692), .Y(n_704) );
AND2x4_ASAP7_75t_L g705 ( .A(n_691), .B(n_696), .Y(n_705) );
INVx3_ASAP7_75t_SL g706 ( .A(n_691), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_698), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_706), .Y(n_708) );
NOR4xp25_ASAP7_75t_L g709 ( .A(n_704), .B(n_694), .C(n_700), .D(n_689), .Y(n_709) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_704), .A2(n_694), .B(n_688), .C(n_695), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_708), .B(n_705), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_711), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_711), .B(n_705), .Y(n_714) );
AOI322xp5_ASAP7_75t_L g715 ( .A1(n_713), .A2(n_712), .A3(n_709), .B1(n_693), .B2(n_703), .C1(n_707), .C2(n_697), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_713), .B(n_714), .Y(n_716) );
endmodule