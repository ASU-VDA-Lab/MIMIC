module fake_jpeg_3268_n_108 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_64),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_69),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_52),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_33),
.B1(n_32),
.B2(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_1),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_50),
.B1(n_32),
.B2(n_3),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_50),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_50),
.C(n_2),
.Y(n_79)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_80),
.Y(n_88)
);

NAND2xp67_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_85),
.Y(n_93)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_28),
.B1(n_10),
.B2(n_12),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_86),
.B(n_4),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_5),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_74),
.B(n_69),
.C(n_71),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_94),
.B1(n_95),
.B2(n_80),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_17),
.C(n_23),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_14),
.C(n_20),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_82),
.B1(n_80),
.B2(n_7),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_88),
.B1(n_93),
.B2(n_87),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_100),
.B1(n_97),
.B2(n_98),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_97),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_9),
.C(n_19),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_18),
.C(n_26),
.Y(n_106)
);

AO21x1_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_5),
.B(n_6),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_6),
.Y(n_108)
);


endmodule