module fake_netlist_1_203_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_10), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_6), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_11), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_13), .B(n_0), .Y(n_19) );
INVx2_ASAP7_75t_SL g20 ( .A(n_15), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_14), .B(n_0), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_16), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_14), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_18), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_19), .A2(n_12), .B1(n_17), .B2(n_1), .Y(n_26) );
INVx3_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_24), .B(n_2), .Y(n_28) );
INVx2_ASAP7_75t_SL g29 ( .A(n_26), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_27), .B(n_25), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_27), .B(n_2), .Y(n_31) );
XOR2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_29), .Y(n_32) );
NAND2xp33_ASAP7_75t_SL g33 ( .A(n_31), .B(n_27), .Y(n_33) );
A2O1A1Ixp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_28), .B(n_3), .C(n_5), .Y(n_34) );
INVx2_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_35), .Y(n_36) );
HB1xp67_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
NAND3xp33_ASAP7_75t_L g39 ( .A(n_38), .B(n_37), .C(n_33), .Y(n_39) );
endmodule