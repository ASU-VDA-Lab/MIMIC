module fake_jpeg_8482_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_40),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_38),
.B1(n_42),
.B2(n_36),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_49),
.B1(n_51),
.B2(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_18),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_21),
.B1(n_33),
.B2(n_16),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_21),
.B1(n_33),
.B2(n_24),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_52),
.B(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_21),
.B1(n_33),
.B2(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_22),
.B(n_30),
.C(n_19),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_27),
.B1(n_28),
.B2(n_18),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_67),
.B1(n_32),
.B2(n_23),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_22),
.B1(n_31),
.B2(n_24),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_70),
.B1(n_26),
.B2(n_25),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_32),
.B1(n_23),
.B2(n_29),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_36),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_83),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_90),
.B1(n_69),
.B2(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_75),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_45),
.Y(n_97)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_70),
.B1(n_66),
.B2(n_56),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_29),
.B(n_26),
.C(n_25),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_25),
.B1(n_46),
.B2(n_47),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_92),
.Y(n_116)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_26),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_51),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_106),
.B1(n_111),
.B2(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_74),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_53),
.C(n_63),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_109),
.C(n_73),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_27),
.Y(n_144)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_81),
.B1(n_71),
.B2(n_94),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_46),
.B1(n_65),
.B2(n_50),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_54),
.C(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_46),
.B1(n_44),
.B2(n_20),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_62),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_44),
.B1(n_18),
.B2(n_20),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_28),
.B(n_20),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_71),
.B(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_44),
.B1(n_18),
.B2(n_20),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_88),
.B1(n_84),
.B2(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_86),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_129),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_96),
.B1(n_97),
.B2(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_132),
.B1(n_95),
.B2(n_98),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_100),
.C(n_109),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_107),
.A2(n_78),
.B1(n_85),
.B2(n_87),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_107),
.B1(n_118),
.B2(n_102),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_138),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_143),
.B(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_94),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_104),
.B(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_15),
.Y(n_171)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_74),
.B1(n_84),
.B2(n_78),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_28),
.B(n_20),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_27),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_108),
.B(n_28),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_28),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_104),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_0),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_148),
.A2(n_151),
.B(n_134),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_156),
.C(n_157),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_143),
.B(n_140),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_152),
.B(n_164),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_141),
.B1(n_132),
.B2(n_145),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_109),
.B1(n_101),
.B2(n_114),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_167),
.B1(n_143),
.B2(n_124),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_101),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_120),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_111),
.B1(n_112),
.B2(n_106),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_158),
.A2(n_162),
.B1(n_168),
.B2(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_159),
.B(n_173),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_107),
.B1(n_68),
.B2(n_60),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_60),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_174),
.C(n_146),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_68),
.B1(n_60),
.B2(n_55),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_27),
.B1(n_80),
.B2(n_79),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_170),
.B(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_162),
.B1(n_151),
.B2(n_168),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_177),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_139),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_136),
.B(n_123),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_190),
.B(n_192),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_184),
.A2(n_194),
.B1(n_199),
.B2(n_158),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_146),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_189),
.C(n_198),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_167),
.B1(n_150),
.B2(n_161),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_122),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_148),
.A2(n_134),
.B(n_135),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_175),
.Y(n_208)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_0),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_169),
.A2(n_142),
.B1(n_130),
.B2(n_138),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_197),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_144),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_142),
.B1(n_133),
.B2(n_130),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_131),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_142),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_80),
.C(n_79),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_202),
.A2(n_210),
.B1(n_196),
.B2(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_208),
.B1(n_187),
.B2(n_178),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_154),
.B1(n_175),
.B2(n_163),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_154),
.B1(n_165),
.B2(n_131),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_212),
.A2(n_213),
.B1(n_220),
.B2(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_163),
.B1(n_171),
.B2(n_174),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_55),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_218),
.C(n_225),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_105),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_217),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_105),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_80),
.B1(n_79),
.B2(n_2),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_193),
.CI(n_184),
.CON(n_227),
.SN(n_227)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_176),
.B1(n_182),
.B2(n_201),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_80),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_79),
.C(n_1),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_190),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_222),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_228),
.A2(n_240),
.B(n_243),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_206),
.C(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_177),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_235),
.B(n_238),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_236),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_196),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_239),
.A2(n_244),
.B1(n_246),
.B2(n_15),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_242),
.B1(n_216),
.B2(n_183),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_207),
.A2(n_178),
.B1(n_195),
.B2(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_227),
.B(n_15),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_249),
.Y(n_277)
);

OAI321xp33_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_213),
.A3(n_208),
.B1(n_209),
.B2(n_203),
.C(n_179),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_206),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_255),
.C(n_258),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_233),
.B(n_229),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_237),
.A2(n_226),
.B1(n_217),
.B2(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_231),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_179),
.B(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_227),
.B1(n_245),
.B2(n_2),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_1),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_14),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_248),
.B(n_14),
.CI(n_1),
.CON(n_274),
.SN(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_0),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_280),
.Y(n_281)
);

AOI211xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_258),
.B(n_4),
.C(n_5),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_1),
.C(n_3),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_259),
.C(n_256),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_262),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_290),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_291),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_252),
.B1(n_260),
.B2(n_253),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_292),
.B1(n_274),
.B2(n_5),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_251),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_287),
.C(n_289),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_255),
.C(n_257),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_263),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_265),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_294),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_269),
.B(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_300),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_267),
.B1(n_272),
.B2(n_269),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_277),
.B(n_6),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_277),
.C(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_6),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_3),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_306),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_307),
.B(n_304),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_293),
.B(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_3),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.C(n_12),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_297),
.B(n_298),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_314),
.C(n_12),
.Y(n_316)
);

A2O1A1O1Ixp25_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_6),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_310),
.B(n_8),
.C(n_10),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_7),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_315),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_7),
.Y(n_320)
);


endmodule