module real_jpeg_2597_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_1),
.A2(n_54),
.B1(n_56),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_1),
.A2(n_68),
.B1(n_69),
.B2(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_2),
.A2(n_36),
.B1(n_38),
.B2(n_59),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_2),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_2),
.A2(n_59),
.B1(n_68),
.B2(n_69),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_4),
.A2(n_54),
.B1(n_56),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_36),
.B1(n_38),
.B2(n_73),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_4),
.A2(n_68),
.B1(n_69),
.B2(n_73),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_5),
.A2(n_68),
.B1(n_69),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_5),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_5),
.A2(n_54),
.B1(n_56),
.B2(n_86),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_25),
.B(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_11),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_11),
.B(n_38),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_11),
.B(n_65),
.C(n_69),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_11),
.A2(n_30),
.B1(n_54),
.B2(n_56),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_11),
.B(n_57),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_11),
.B(n_83),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_11),
.B(n_77),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_11),
.A2(n_38),
.B(n_145),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_40),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_12),
.A2(n_36),
.B1(n_38),
.B2(n_40),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_12),
.A2(n_40),
.B1(n_54),
.B2(n_56),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_12),
.A2(n_40),
.B1(n_68),
.B2(n_69),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_13),
.A2(n_36),
.B1(n_38),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_46),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_13),
.A2(n_46),
.B1(n_54),
.B2(n_56),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_13),
.A2(n_46),
.B1(n_68),
.B2(n_69),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_132),
.B1(n_208),
.B2(n_209),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_18),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_102),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_92),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_21),
.A2(n_22),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_23),
.B(n_42),
.C(n_61),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_35),
.B2(n_39),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_30),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_26),
.B(n_34),
.C(n_38),
.Y(n_91)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_29),
.A2(n_33),
.B(n_36),
.C(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_30),
.A2(n_81),
.B1(n_83),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_31),
.A2(n_35),
.B1(n_39),
.B2(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_35)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_38),
.B1(n_50),
.B2(n_52),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_36),
.B(n_52),
.C(n_56),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_60),
.B2(n_61),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_57),
.B2(n_58),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_45),
.A2(n_48),
.B1(n_53),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_48),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_48),
.A2(n_53),
.B1(n_101),
.B2(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_50),
.A2(n_54),
.B(n_144),
.C(n_146),
.Y(n_143)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_54),
.B(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_57),
.B(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_72),
.B(n_74),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_62),
.A2(n_127),
.B1(n_140),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_63),
.B(n_75),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_63),
.A2(n_139),
.B(n_141),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_63),
.A2(n_77),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_63),
.A2(n_77),
.B1(n_164),
.B2(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_67),
.B(n_72),
.Y(n_141)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_69),
.B(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_78),
.A2(n_92),
.B1(n_93),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_89),
.B2(n_90),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_81),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_81),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_81),
.A2(n_83),
.B1(n_179),
.B2(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_85),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_82),
.B(n_148),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_82),
.A2(n_123),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_96),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_87),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.C(n_100),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_116),
.B2(n_117),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_125),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_125),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_153),
.B(n_207),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_149),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_149),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_142),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_135),
.B(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_138),
.B(n_142),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_143),
.B(n_147),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_202),
.B(n_206),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_192),
.B(n_201),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_173),
.B(n_191),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_165),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_170),
.C(n_172),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_185),
.B(n_190),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_180),
.B(n_184),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_183),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_189),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_193),
.B(n_194),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_205),
.Y(n_206)
);


endmodule