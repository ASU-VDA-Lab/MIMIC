module fake_jpeg_3555_n_186 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_31),
.C(n_26),
.Y(n_70)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_19),
.B1(n_24),
.B2(n_23),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_32),
.Y(n_53)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_6),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_55),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_79),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_64),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_44),
.B1(n_39),
.B2(n_36),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_30),
.Y(n_64)
);

OR2x2_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_30),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_18),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_10),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_72),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_76),
.B1(n_50),
.B2(n_41),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_35),
.A2(n_19),
.B1(n_4),
.B2(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_6),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_19),
.Y(n_79)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_40),
.B1(n_42),
.B2(n_48),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_96),
.B1(n_97),
.B2(n_68),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_102),
.Y(n_114)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_101),
.Y(n_109)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_10),
.Y(n_101)
);

NOR2x1p5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_12),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_98),
.B(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_77),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_80),
.A2(n_71),
.B1(n_56),
.B2(n_73),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_57),
.B1(n_77),
.B2(n_56),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_66),
.C(n_57),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_84),
.C(n_104),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_116),
.B1(n_117),
.B2(n_123),
.Y(n_137)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_68),
.B(n_56),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_89),
.B(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_122),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_139),
.C(n_141),
.Y(n_146)
);

AO22x1_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_85),
.B1(n_87),
.B2(n_97),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_130),
.B(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_103),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_121),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_137),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_107),
.C(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_115),
.C(n_106),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_107),
.B1(n_115),
.B2(n_112),
.Y(n_141)
);

XOR2x1_ASAP7_75t_SL g145 ( 
.A(n_138),
.B(n_113),
.Y(n_145)
);

OAI31xp33_ASAP7_75t_SL g158 ( 
.A1(n_145),
.A2(n_133),
.A3(n_137),
.B(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_106),
.C(n_112),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_150),
.C(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_152),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_118),
.C(n_108),
.Y(n_150)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_108),
.B(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_151),
.B(n_153),
.C(n_161),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_141),
.B1(n_136),
.B2(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_135),
.Y(n_160)
);

OA21x2_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_153),
.B(n_157),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_129),
.B1(n_140),
.B2(n_126),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_158),
.C(n_155),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_164),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_145),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_168),
.B(n_171),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_167),
.B(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_168),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_172),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_176),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_180),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_177),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_179),
.C(n_184),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_179),
.Y(n_186)
);


endmodule