module real_jpeg_16514_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_295;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_127;
wire n_53;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_4),
.B1(n_19),
.B2(n_20),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_1),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_2),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_2),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_2),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_3),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_3),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_3),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_5),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_5),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_5),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_5),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_5),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_6),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_6),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_6),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_6),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_6),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_6),
.B(n_234),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_7),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_8),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_8),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_9),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_9),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_10),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_11),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_11),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_11),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_11),
.B(n_265),
.Y(n_264)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_13),
.B(n_33),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_13),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_13),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_13),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_13),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_13),
.B(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g153 ( 
.A(n_15),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_16),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_16),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_16),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_16),
.B(n_73),
.Y(n_254)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_183),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_182),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_156),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_23),
.B(n_156),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_105),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_69),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_28),
.Y(n_178)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

XNOR2x2_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_57),
.Y(n_43)
);

MAJx2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.C(n_53),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_45),
.B(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_48),
.Y(n_148)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_56),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_65),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_83),
.C(n_96),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_70),
.B(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_79),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

MAJx3_ASAP7_75t_L g144 ( 
.A(n_72),
.B(n_76),
.C(n_79),
.Y(n_144)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_75),
.Y(n_206)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_82),
.B(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_83),
.A2(n_84),
.B1(n_96),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_85),
.A2(n_89),
.B1(n_90),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_85),
.Y(n_170)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.C(n_103),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_97),
.A2(n_103),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_97),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_102),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_103),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_140),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_123),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_111),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_116),
.B(n_122),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_118),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_133),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_124),
.A2(n_125),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_126),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_126),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g226 ( 
.A(n_127),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_128),
.A2(n_133),
.B1(n_134),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_128),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2x2_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_154),
.B(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_164),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_157),
.A2(n_158),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_164),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.C(n_171),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_165),
.B(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_169),
.B(n_171),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.C(n_179),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_172),
.A2(n_173),
.B1(n_179),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_177),
.B(n_277),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_179),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21x1_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_292),
.B(n_298),
.Y(n_184)
);

AOI21x1_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_280),
.B(n_291),
.Y(n_185)
);

OAI21x1_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_256),
.B(n_279),
.Y(n_186)
);

AOI21x1_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_229),
.B(n_255),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_215),
.B(n_228),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_198),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_190),
.B(n_198),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_195),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_209),
.C(n_211),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_200),
.B(n_202),
.Y(n_251)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_224),
.B(n_227),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_223),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_223),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_249),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_251),
.C(n_252),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_245),
.C(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_258),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_273),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_274),
.C(n_276),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_266),
.C(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_266),
.B1(n_271),
.B2(n_272),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_290),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_SL g291 ( 
.A(n_281),
.B(n_290),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_287),
.C(n_288),
.Y(n_297)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_297),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);


endmodule