module real_aes_5206_n_15 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_15);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_15;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_0), .Y(n_26) );
AOI322xp5_ASAP7_75t_SL g32 ( .A1(n_1), .A2(n_7), .A3(n_29), .B1(n_33), .B2(n_34), .C1(n_41), .C2(n_46), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_2), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g40 ( .A(n_2), .B(n_6), .Y(n_40) );
NOR2xp33_ASAP7_75t_R g20 ( .A(n_3), .B(n_21), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_4), .Y(n_27) );
NOR4xp25_ASAP7_75t_SL g18 ( .A(n_5), .B(n_19), .C(n_25), .D(n_26), .Y(n_18) );
NAND2xp33_ASAP7_75t_R g30 ( .A(n_5), .B(n_20), .Y(n_30) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_5), .Y(n_39) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_6), .B(n_18), .Y(n_17) );
NAND2xp33_ASAP7_75t_R g28 ( .A(n_6), .B(n_29), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_6), .Y(n_33) );
NAND3xp33_ASAP7_75t_SL g21 ( .A(n_8), .B(n_22), .C(n_23), .Y(n_21) );
NOR2xp33_ASAP7_75t_R g24 ( .A(n_9), .B(n_10), .Y(n_24) );
NOR3xp33_ASAP7_75t_SL g36 ( .A(n_9), .B(n_37), .C(n_38), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_10), .Y(n_37) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_11), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_12), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_13), .Y(n_23) );
BUFx8_ASAP7_75t_SL g45 ( .A(n_14), .Y(n_45) );
OAI221xp5_ASAP7_75t_R g15 ( .A1(n_16), .A2(n_17), .B1(n_27), .B2(n_28), .C(n_32), .Y(n_15) );
NAND2xp33_ASAP7_75t_R g48 ( .A(n_18), .B(n_33), .Y(n_48) );
NAND2xp33_ASAP7_75t_R g19 ( .A(n_20), .B(n_24), .Y(n_19) );
NAND3xp33_ASAP7_75t_SL g38 ( .A(n_20), .B(n_26), .C(n_39), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_24), .Y(n_31) );
NOR4xp25_ASAP7_75t_SL g29 ( .A(n_25), .B(n_26), .C(n_30), .D(n_31), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_35), .Y(n_34) );
NAND2xp33_ASAP7_75t_R g35 ( .A(n_36), .B(n_40), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g41 ( .A(n_42), .Y(n_41) );
CKINVDCx20_ASAP7_75t_R g42 ( .A(n_43), .Y(n_42) );
CKINVDCx20_ASAP7_75t_R g43 ( .A(n_44), .Y(n_43) );
CKINVDCx20_ASAP7_75t_R g44 ( .A(n_45), .Y(n_44) );
HB1xp67_ASAP7_75t_L g46 ( .A(n_47), .Y(n_46) );
CKINVDCx5p33_ASAP7_75t_R g47 ( .A(n_48), .Y(n_47) );
endmodule