module fake_jpeg_31047_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_13),
.B(n_7),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_15),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_17),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_20),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_73),
.C(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_86),
.Y(n_88)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_0),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_56),
.B1(n_72),
.B2(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_95),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_93),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_66),
.B(n_57),
.C(n_58),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_71),
.B(n_61),
.Y(n_120)
);

NAND2x1_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_77),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_76),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_104),
.A2(n_116),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_117),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_120),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_69),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_67),
.B1(n_84),
.B2(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_63),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_55),
.B(n_59),
.C(n_60),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_3),
.B(n_4),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_69),
.B1(n_75),
.B2(n_64),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_54),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_2),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_102),
.B(n_0),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_1),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_30),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_75),
.B1(n_102),
.B2(n_101),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_142),
.B1(n_9),
.B2(n_10),
.Y(n_154)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_135),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_133),
.Y(n_149)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_3),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_143),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_4),
.B(n_5),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_12),
.B(n_13),
.Y(n_156)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_155),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_119),
.B1(n_118),
.B2(n_11),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_154),
.B1(n_163),
.B2(n_125),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_27),
.C(n_49),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_138),
.C(n_31),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_11),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_159),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_12),
.B(n_14),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_157),
.A2(n_158),
.B(n_129),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_35),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_34),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_161),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_16),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_167),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_147),
.A2(n_124),
.B1(n_134),
.B2(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_168),
.B(n_170),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_29),
.B(n_39),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_160),
.C(n_150),
.Y(n_177)
);

OAI321xp33_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_159),
.A3(n_148),
.B1(n_163),
.B2(n_149),
.C(n_162),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_173),
.B(n_169),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_164),
.C(n_170),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_175),
.B1(n_178),
.B2(n_168),
.Y(n_182)
);

AO32x1_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_176),
.A3(n_175),
.B1(n_156),
.B2(n_157),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_153),
.C(n_172),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_151),
.C(n_42),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_151),
.B1(n_43),
.B2(n_45),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_40),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_50),
.Y(n_188)
);


endmodule