module fake_jpeg_5812_n_188 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_1),
.B(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_1),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_18),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_5),
.Y(n_77)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_21),
.Y(n_49)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_53),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_27),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_54),
.B(n_69),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_46),
.B1(n_30),
.B2(n_41),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_59),
.B1(n_70),
.B2(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_45),
.B(n_16),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_29),
.B(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_60),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_30),
.B1(n_18),
.B2(n_31),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_75),
.B1(n_11),
.B2(n_64),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_29),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_21),
.B(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_23),
.B1(n_14),
.B2(n_20),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_33),
.A2(n_26),
.B1(n_20),
.B2(n_19),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_72),
.B1(n_78),
.B2(n_67),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_26),
.B1(n_20),
.B2(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_4),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_57),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_9),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_10),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_59),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_61),
.C(n_51),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_102),
.Y(n_113)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_99),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_52),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_78),
.B1(n_67),
.B2(n_55),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_73),
.B1(n_68),
.B2(n_74),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_48),
.B1(n_49),
.B2(n_62),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_53),
.B1(n_61),
.B2(n_51),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_124),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_61),
.B1(n_96),
.B2(n_81),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_81),
.B1(n_102),
.B2(n_80),
.Y(n_130)
);

CKINVDCx12_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_119),
.Y(n_133)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_83),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_87),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_61),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_85),
.B1(n_106),
.B2(n_103),
.C(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_92),
.B1(n_95),
.B2(n_88),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_136),
.B1(n_129),
.B2(n_128),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_112),
.C(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_139),
.C(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_86),
.C(n_101),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_116),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_140),
.B(n_141),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_123),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_103),
.C(n_106),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_107),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_148),
.B1(n_126),
.B2(n_107),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_134),
.B1(n_127),
.B2(n_111),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_109),
.B(n_120),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_131),
.B(n_111),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_137),
.C(n_126),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_109),
.B(n_120),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_84),
.B(n_89),
.Y(n_164)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_149),
.B(n_131),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_156),
.A2(n_161),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_163),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_152),
.C(n_148),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_164),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_171),
.B(n_150),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_175),
.C(n_169),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_158),
.A3(n_144),
.B1(n_164),
.B2(n_163),
.C1(n_166),
.C2(n_150),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_172),
.A2(n_158),
.B1(n_160),
.B2(n_165),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_160),
.B(n_170),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_161),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_181),
.B(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_100),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_147),
.B(n_171),
.Y(n_181)
);

OAI321xp33_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_161),
.A3(n_175),
.B1(n_168),
.B2(n_173),
.C(n_142),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_184),
.A2(n_79),
.B(n_133),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_79),
.B(n_94),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_187),
.B1(n_183),
.B2(n_86),
.C(n_99),
.Y(n_188)
);


endmodule