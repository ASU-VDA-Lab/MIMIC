module fake_netlist_6_1605_n_272 (n_52, n_16, n_1, n_46, n_18, n_21, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_5, n_77, n_42, n_8, n_24, n_54, n_0, n_32, n_66, n_78, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_80, n_41, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_272);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_5;
input n_77;
input n_42;
input n_8;
input n_24;
input n_54;
input n_0;
input n_32;
input n_66;
input n_78;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_80;
input n_41;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_272;

wire n_91;
wire n_146;
wire n_163;
wire n_119;
wire n_235;
wire n_256;
wire n_193;
wire n_147;
wire n_269;
wire n_258;
wire n_154;
wire n_191;
wire n_88;
wire n_209;
wire n_98;
wire n_260;
wire n_265;
wire n_113;
wire n_223;
wire n_270;
wire n_148;
wire n_199;
wire n_161;
wire n_138;
wire n_208;
wire n_228;
wire n_226;
wire n_252;
wire n_266;
wire n_166;
wire n_184;
wire n_212;
wire n_268;
wire n_271;
wire n_158;
wire n_216;
wire n_210;
wire n_83;
wire n_206;
wire n_217;
wire n_167;
wire n_101;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_145;
wire n_92;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_131;
wire n_105;
wire n_227;
wire n_132;
wire n_188;
wire n_186;
wire n_102;
wire n_204;
wire n_245;
wire n_87;
wire n_195;
wire n_261;
wire n_189;
wire n_85;
wire n_130;
wire n_99;
wire n_84;
wire n_213;
wire n_257;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_203;
wire n_254;
wire n_142;
wire n_143;
wire n_207;
wire n_242;
wire n_180;
wire n_155;
wire n_219;
wire n_109;
wire n_150;
wire n_233;
wire n_263;
wire n_122;
wire n_264;
wire n_255;
wire n_205;
wire n_140;
wire n_218;
wire n_120;
wire n_234;
wire n_251;
wire n_214;
wire n_82;
wire n_236;
wire n_246;
wire n_110;
wire n_151;
wire n_112;
wire n_172;
wire n_237;
wire n_244;
wire n_181;
wire n_182;
wire n_124;
wire n_238;
wire n_239;
wire n_126;
wire n_202;
wire n_94;
wire n_97;
wire n_108;
wire n_267;
wire n_116;
wire n_211;
wire n_220;
wire n_117;
wire n_118;
wire n_175;
wire n_224;
wire n_231;
wire n_230;
wire n_93;
wire n_141;
wire n_240;
wire n_135;
wire n_196;
wire n_200;
wire n_165;
wire n_139;
wire n_134;
wire n_259;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_95;
wire n_179;
wire n_248;
wire n_243;
wire n_107;
wire n_229;
wire n_253;
wire n_190;
wire n_123;
wire n_262;
wire n_136;
wire n_187;
wire n_89;
wire n_249;
wire n_173;
wire n_201;
wire n_250;
wire n_103;
wire n_111;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_232;
wire n_115;
wire n_128;
wire n_241;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_221;

INVx1_ASAP7_75t_SL g82 ( 
.A(n_28),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

INVxp33_ASAP7_75t_SL g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_57),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_25),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_6),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_35),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_19),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_14),
.Y(n_113)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_0),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_13),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_62),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_1),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

NAND2x1p5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_10),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_84),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

AND3x2_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_1),
.C(n_3),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_4),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_5),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_87),
.B(n_5),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_147)
);

AND2x4_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_7),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_8),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_97),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_113),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_97),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_93),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_125),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_112),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_110),
.B1(n_100),
.B2(n_108),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_126),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_100),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_144),
.B1(n_150),
.B2(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_165),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_152),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_134),
.Y(n_177)
);

AND2x4_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_127),
.Y(n_178)
);

OR2x6_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_147),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_131),
.B(n_83),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_146),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_83),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_82),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_118),
.B(n_123),
.C(n_122),
.Y(n_188)
);

AND2x4_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_138),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_99),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_96),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_104),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_92),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_107),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_115),
.B1(n_102),
.B2(n_105),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_101),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_117),
.B1(n_106),
.B2(n_109),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_159),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_162),
.Y(n_206)
);

O2A1O1Ixp5_ASAP7_75t_SL g207 ( 
.A1(n_195),
.A2(n_168),
.B(n_164),
.C(n_9),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_196),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_119),
.B(n_168),
.C(n_164),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_168),
.B(n_164),
.C(n_15),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_20),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_179),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

OAI21x1_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_185),
.B(n_180),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_207),
.A2(n_177),
.B(n_191),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_194),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

OAI21x1_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_183),
.B(n_26),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_29),
.B(n_36),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_38),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_48),
.B(n_49),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

AO21x2_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_50),
.B(n_51),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_224),
.A2(n_216),
.B1(n_220),
.B2(n_227),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_210),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_218),
.A2(n_205),
.B(n_204),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_217),
.B1(n_202),
.B2(n_205),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_223),
.B(n_225),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_209),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_53),
.Y(n_239)
);

BUFx4f_ASAP7_75t_SL g240 ( 
.A(n_238),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_222),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_231),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_226),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_231),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_233),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

AO21x2_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_232),
.B(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_243),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_246),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_252),
.Y(n_256)
);

OR2x6_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_247),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_R g258 ( 
.A(n_254),
.B(n_250),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_258),
.B(n_250),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_259),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_261),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_260),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

NOR3xp33_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_251),
.C(n_257),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_67),
.B(n_72),
.Y(n_270)
);

AO221x1_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.C(n_80),
.Y(n_271)
);

OA21x2_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_81),
.B(n_253),
.Y(n_272)
);


endmodule