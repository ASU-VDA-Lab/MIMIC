module fake_jpeg_3355_n_195 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_195);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_26),
.Y(n_59)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_46),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_31),
.C(n_29),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_53),
.B1(n_62),
.B2(n_28),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_22),
.B1(n_29),
.B2(n_23),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_31),
.B1(n_24),
.B2(n_20),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_64),
.B1(n_65),
.B2(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_23),
.B1(n_29),
.B2(n_14),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_27),
.B1(n_17),
.B2(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_66),
.B(n_17),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_68),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_27),
.B(n_16),
.C(n_30),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_44),
.B1(n_39),
.B2(n_23),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_71),
.B(n_75),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_77),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_16),
.B1(n_30),
.B2(n_28),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_81),
.B1(n_13),
.B2(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_78),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_8),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_80),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_5),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

OA22x2_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_86),
.B1(n_90),
.B2(n_97),
.Y(n_108)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_5),
.B1(n_1),
.B2(n_3),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_91),
.Y(n_99)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_0),
.B(n_4),
.C(n_10),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_52),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_10),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_86),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_87),
.B1(n_80),
.B2(n_70),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_13),
.C(n_94),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_105),
.B(n_114),
.C(n_106),
.D(n_90),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_13),
.B1(n_74),
.B2(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_113),
.B1(n_69),
.B2(n_73),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_69),
.B1(n_68),
.B2(n_84),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_91),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_77),
.B1(n_84),
.B2(n_90),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_113),
.B(n_108),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_129),
.B1(n_136),
.B2(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_92),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_127),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_69),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_134),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_95),
.B1(n_96),
.B2(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_146),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_145),
.B1(n_147),
.B2(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_109),
.C(n_102),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_128),
.C(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_147),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_111),
.B(n_109),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_110),
.B(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_103),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_122),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_151),
.A2(n_124),
.B1(n_133),
.B2(n_136),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_99),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_158),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_108),
.B1(n_129),
.B2(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_156),
.B1(n_161),
.B2(n_163),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_101),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_160),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_151),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_164),
.B(n_150),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_138),
.C(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_171),
.C(n_172),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_152),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_141),
.C(n_148),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_146),
.C(n_150),
.Y(n_172)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_169),
.B(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_155),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_175),
.A2(n_173),
.B1(n_165),
.B2(n_163),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_178),
.C(n_179),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_157),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_152),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_164),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_167),
.C(n_154),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

OAI21x1_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_176),
.B(n_166),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_185),
.B(n_177),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_186),
.A2(n_183),
.B(n_177),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_189),
.A2(n_181),
.B(n_88),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_190),
.C(n_117),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_82),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_89),
.Y(n_195)
);


endmodule