module fake_aes_4898_n_441 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_441);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_441;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_73;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NOR2xp67_ASAP7_75t_L g64 ( .A(n_61), .B(n_8), .Y(n_64) );
BUFx6f_ASAP7_75t_L g65 ( .A(n_30), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_63), .Y(n_66) );
INVx1_ASAP7_75t_L g67 ( .A(n_45), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_60), .Y(n_68) );
INVxp67_ASAP7_75t_SL g69 ( .A(n_24), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_7), .Y(n_70) );
CKINVDCx5p33_ASAP7_75t_R g71 ( .A(n_17), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_57), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_56), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_27), .Y(n_74) );
INVxp67_ASAP7_75t_L g75 ( .A(n_58), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_10), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_49), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_3), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_1), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_23), .Y(n_80) );
OR2x2_ASAP7_75t_L g81 ( .A(n_55), .B(n_39), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_18), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_36), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_9), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_47), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_28), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_0), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_46), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_38), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g94 ( .A(n_8), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_62), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_12), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_40), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_41), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_21), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_22), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_33), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_94), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_82), .Y(n_104) );
INVx3_ASAP7_75t_L g105 ( .A(n_82), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
NOR2xp33_ASAP7_75t_R g107 ( .A(n_101), .B(n_32), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_67), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_68), .Y(n_109) );
AND2x4_ASAP7_75t_L g110 ( .A(n_70), .B(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_68), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_94), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_101), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_71), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_83), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_71), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_70), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_72), .Y(n_118) );
XNOR2xp5_ASAP7_75t_L g119 ( .A(n_76), .B(n_1), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_65), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_78), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_72), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_110), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_106), .B(n_66), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_110), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_116), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_110), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_110), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_120), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_118), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_118), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_120), .Y(n_134) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_106), .B(n_81), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_115), .B(n_97), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_120), .Y(n_137) );
OAI221xp5_ASAP7_75t_L g138 ( .A1(n_117), .A2(n_79), .B1(n_78), .B2(n_85), .C(n_96), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_108), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_108), .A2(n_79), .B1(n_90), .B2(n_93), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_109), .B(n_80), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_121), .B(n_87), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_114), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_122), .B(n_75), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_123), .B(n_89), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_132), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_133), .Y(n_148) );
NAND2x1_ASAP7_75t_L g149 ( .A(n_124), .B(n_126), .Y(n_149) );
OR2x2_ASAP7_75t_L g150 ( .A(n_127), .B(n_113), .Y(n_150) );
AOI211xp5_ASAP7_75t_L g151 ( .A1(n_138), .A2(n_119), .B(n_113), .C(n_123), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_136), .B(n_109), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_127), .Y(n_153) );
BUFx3_ASAP7_75t_L g154 ( .A(n_135), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
NOR3xp33_ASAP7_75t_SL g156 ( .A(n_144), .B(n_119), .C(n_111), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_135), .B(n_111), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_135), .Y(n_158) );
NOR3xp33_ASAP7_75t_SL g159 ( .A(n_138), .B(n_88), .C(n_69), .Y(n_159) );
BUFx2_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_146), .B(n_105), .Y(n_161) );
INVx3_ASAP7_75t_SL g162 ( .A(n_133), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_124), .A2(n_104), .B1(n_73), .B2(n_74), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_136), .B(n_105), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_126), .A2(n_73), .B1(n_74), .B2(n_77), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_133), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_146), .B(n_105), .Y(n_167) );
NOR2xp67_ASAP7_75t_L g168 ( .A(n_128), .B(n_81), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_146), .B(n_64), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_136), .B(n_84), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_128), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_130), .B(n_107), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_130), .Y(n_176) );
BUFx4f_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g179 ( .A1(n_154), .A2(n_143), .B1(n_142), .B2(n_125), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_157), .B(n_125), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_149), .A2(n_142), .B(n_145), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_154), .B(n_143), .Y(n_182) );
BUFx12f_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_177), .B(n_140), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_158), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_170), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_176), .A2(n_141), .B1(n_100), .B2(n_77), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_177), .B(n_160), .Y(n_188) );
BUFx12f_ASAP7_75t_L g189 ( .A(n_160), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_176), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_170), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_173), .A2(n_99), .B(n_100), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_152), .B(n_86), .Y(n_195) );
INVx1_ASAP7_75t_SL g196 ( .A(n_162), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_173), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_177), .B(n_103), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_174), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_153), .B(n_112), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_174), .B(n_65), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_152), .B(n_174), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_174), .B(n_91), .Y(n_204) );
OAI22xp5_ASAP7_75t_SL g205 ( .A1(n_151), .A2(n_92), .B1(n_95), .B2(n_98), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_161), .B(n_102), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_150), .B(n_2), .Y(n_207) );
AND2x4_ASAP7_75t_SL g208 ( .A(n_147), .B(n_65), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_183), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_179), .A2(n_168), .B1(n_165), .B2(n_163), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_183), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_181), .A2(n_149), .B(n_168), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_186), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_191), .B(n_147), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_193), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_183), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_207), .Y(n_217) );
OAI221xp5_ASAP7_75t_L g218 ( .A1(n_205), .A2(n_150), .B1(n_156), .B2(n_172), .C(n_159), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_205), .A2(n_161), .B1(n_167), .B2(n_171), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_179), .A2(n_165), .B1(n_163), .B2(n_169), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_183), .B(n_167), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_191), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g223 ( .A1(n_207), .A2(n_164), .B1(n_169), .B2(n_167), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_189), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_184), .B(n_167), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_207), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_188), .B(n_161), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_205), .A2(n_161), .B1(n_171), .B2(n_166), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_180), .A2(n_166), .B1(n_171), .B2(n_148), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_180), .A2(n_166), .B1(n_171), .B2(n_148), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_186), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_182), .A2(n_166), .B1(n_175), .B2(n_155), .Y(n_232) );
OAI211xp5_ASAP7_75t_L g233 ( .A1(n_194), .A2(n_155), .B(n_65), .C(n_120), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_182), .B(n_155), .Y(n_234) );
OAI22xp33_ASAP7_75t_L g235 ( .A1(n_221), .A2(n_207), .B1(n_189), .B2(n_185), .Y(n_235) );
AOI222xp33_ASAP7_75t_L g236 ( .A1(n_218), .A2(n_200), .B1(n_198), .B2(n_184), .C1(n_195), .C2(n_189), .Y(n_236) );
AOI221xp5_ASAP7_75t_L g237 ( .A1(n_210), .A2(n_200), .B1(n_195), .B2(n_206), .C(n_182), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_221), .Y(n_238) );
CKINVDCx8_ASAP7_75t_R g239 ( .A(n_209), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_219), .A2(n_200), .B1(n_182), .B2(n_184), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_209), .Y(n_242) );
AOI222xp33_ASAP7_75t_L g243 ( .A1(n_228), .A2(n_200), .B1(n_198), .B2(n_184), .C1(n_189), .C2(n_182), .Y(n_243) );
NAND2xp33_ASAP7_75t_R g244 ( .A(n_211), .B(n_198), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_223), .A2(n_185), .B1(n_182), .B2(n_193), .Y(n_245) );
NAND3xp33_ASAP7_75t_L g246 ( .A(n_212), .B(n_186), .C(n_197), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_220), .A2(n_185), .B1(n_198), .B2(n_188), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
AOI22xp33_ASAP7_75t_SL g249 ( .A1(n_216), .A2(n_185), .B1(n_188), .B2(n_208), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_221), .Y(n_250) );
AOI21x1_ASAP7_75t_L g251 ( .A1(n_217), .A2(n_201), .B(n_197), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_226), .B(n_188), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_214), .Y(n_253) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_213), .A2(n_181), .B(n_197), .Y(n_254) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_213), .A2(n_193), .B(n_201), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_221), .B(n_193), .Y(n_256) );
OAI31xp33_ASAP7_75t_L g257 ( .A1(n_235), .A2(n_216), .A3(n_214), .B(n_225), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_237), .A2(n_206), .B1(n_187), .B2(n_227), .C(n_230), .Y(n_258) );
AO221x2_ASAP7_75t_L g259 ( .A1(n_245), .A2(n_229), .B1(n_231), .B2(n_224), .C(n_211), .Y(n_259) );
OR2x6_ASAP7_75t_L g260 ( .A(n_253), .B(n_214), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_241), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_241), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_248), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_248), .B(n_231), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_253), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_236), .A2(n_224), .B1(n_227), .B2(n_206), .Y(n_266) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_246), .A2(n_233), .B(n_234), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_248), .B(n_227), .Y(n_268) );
NAND4xp25_ASAP7_75t_L g269 ( .A(n_236), .B(n_206), .C(n_187), .D(n_232), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_253), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_254), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_243), .A2(n_178), .B1(n_204), .B2(n_191), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_254), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_254), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_255), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_246), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_273), .Y(n_278) );
NAND4xp25_ASAP7_75t_L g279 ( .A(n_266), .B(n_243), .C(n_240), .D(n_247), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_263), .B(n_256), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_263), .B(n_256), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_271), .Y(n_282) );
NAND3xp33_ASAP7_75t_SL g283 ( .A(n_257), .B(n_239), .C(n_242), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_261), .B(n_252), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_260), .Y(n_285) );
OAI31xp33_ASAP7_75t_SL g286 ( .A1(n_269), .A2(n_249), .A3(n_196), .B(n_244), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_263), .B(n_255), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_266), .B(n_239), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_264), .B(n_238), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_269), .A2(n_238), .B1(n_202), .B2(n_250), .C(n_204), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_271), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_261), .B(n_250), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_264), .B(n_251), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_262), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_265), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_277), .B(n_178), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_265), .Y(n_300) );
AOI33xp33_ASAP7_75t_L g301 ( .A1(n_272), .A2(n_204), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_9), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_260), .A2(n_208), .B1(n_222), .B2(n_191), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_277), .B(n_178), .Y(n_303) );
NOR2xp67_ASAP7_75t_L g304 ( .A(n_283), .B(n_265), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_279), .B(n_289), .Y(n_305) );
NOR4xp25_ASAP7_75t_SL g306 ( .A(n_285), .B(n_257), .C(n_258), .D(n_259), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_290), .B(n_270), .Y(n_308) );
NOR2xp33_ASAP7_75t_R g309 ( .A(n_298), .B(n_265), .Y(n_309) );
OAI21xp5_ASAP7_75t_SL g310 ( .A1(n_286), .A2(n_291), .B(n_279), .Y(n_310) );
OAI33xp33_ASAP7_75t_L g311 ( .A1(n_296), .A2(n_273), .A3(n_276), .B1(n_275), .B2(n_10), .B3(n_11), .Y(n_311) );
AOI33xp33_ASAP7_75t_L g312 ( .A1(n_291), .A2(n_268), .A3(n_273), .B1(n_6), .B2(n_11), .B3(n_12), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_290), .B(n_270), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_293), .Y(n_314) );
NAND2xp33_ASAP7_75t_R g315 ( .A(n_298), .B(n_260), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_294), .B(n_276), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_298), .B(n_270), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_293), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_275), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_281), .B(n_268), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_294), .B(n_276), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_288), .B(n_259), .Y(n_322) );
NOR2xp33_ASAP7_75t_R g323 ( .A(n_298), .B(n_222), .Y(n_323) );
INVx6_ASAP7_75t_L g324 ( .A(n_299), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_292), .B(n_275), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_278), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_297), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_278), .Y(n_328) );
NOR2x1_ASAP7_75t_L g329 ( .A(n_302), .B(n_267), .Y(n_329) );
OAI221xp5_ASAP7_75t_L g330 ( .A1(n_284), .A2(n_202), .B1(n_65), .B2(n_178), .C(n_196), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_284), .B(n_259), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_292), .B(n_267), .Y(n_332) );
OAI21xp5_ASAP7_75t_SL g333 ( .A1(n_302), .A2(n_208), .B(n_222), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_295), .B(n_267), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_287), .B(n_278), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_299), .A2(n_196), .B(n_178), .C(n_203), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_307), .B(n_287), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_333), .A2(n_208), .B(n_300), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_310), .A2(n_303), .B(n_301), .C(n_178), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_320), .B(n_4), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_308), .B(n_4), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_332), .Y(n_342) );
INVx1_ASAP7_75t_SL g343 ( .A(n_309), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_313), .B(n_5), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_335), .B(n_13), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_324), .B(n_14), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_318), .B(n_14), .Y(n_348) );
OAI22xp33_ASAP7_75t_L g349 ( .A1(n_315), .A2(n_191), .B1(n_251), .B2(n_203), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_305), .B(n_331), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g351 ( .A1(n_305), .A2(n_15), .B1(n_16), .B2(n_17), .C(n_18), .Y(n_351) );
NOR2x1_ASAP7_75t_L g352 ( .A(n_304), .B(n_191), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_319), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_316), .B(n_15), .Y(n_354) );
NAND3xp33_ASAP7_75t_L g355 ( .A(n_306), .B(n_129), .C(n_131), .Y(n_355) );
OAI211xp5_ASAP7_75t_L g356 ( .A1(n_323), .A2(n_309), .B(n_336), .C(n_330), .Y(n_356) );
OAI32xp33_ASAP7_75t_L g357 ( .A1(n_315), .A2(n_16), .A3(n_20), .B1(n_192), .B2(n_199), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_316), .B(n_20), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_321), .B(n_25), .Y(n_359) );
NAND2x1_ASAP7_75t_L g360 ( .A(n_324), .B(n_329), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_321), .B(n_26), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_327), .B(n_29), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_322), .B(n_31), .Y(n_363) );
NOR3xp33_ASAP7_75t_SL g364 ( .A(n_311), .B(n_34), .C(n_35), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_323), .B(n_203), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_312), .A2(n_203), .B(n_199), .C(n_190), .Y(n_366) );
AO22x2_ASAP7_75t_L g367 ( .A1(n_332), .A2(n_190), .B1(n_199), .B2(n_192), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
OAI21xp5_ASAP7_75t_SL g369 ( .A1(n_317), .A2(n_203), .B(n_190), .Y(n_369) );
OAI21xp33_ASAP7_75t_L g370 ( .A1(n_312), .A2(n_137), .B(n_129), .Y(n_370) );
OAI221xp5_ASAP7_75t_L g371 ( .A1(n_328), .A2(n_203), .B1(n_190), .B2(n_155), .C(n_192), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_326), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_372), .Y(n_373) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_351), .B(n_325), .C(n_326), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_364), .A2(n_325), .B(n_328), .Y(n_375) );
XNOR2x1_ASAP7_75t_L g376 ( .A(n_340), .B(n_37), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_350), .B(n_42), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_341), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_345), .Y(n_379) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_339), .A2(n_43), .B(n_44), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_353), .Y(n_381) );
OR2x6_ASAP7_75t_L g382 ( .A(n_338), .B(n_203), .Y(n_382) );
NAND3xp33_ASAP7_75t_L g383 ( .A(n_360), .B(n_203), .C(n_134), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_347), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_342), .B(n_48), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_343), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_344), .B(n_50), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_342), .B(n_51), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_337), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_368), .B(n_52), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_354), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
NOR3xp33_ASAP7_75t_SL g393 ( .A(n_356), .B(n_53), .C(n_54), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_346), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
NOR2x1_ASAP7_75t_L g396 ( .A(n_356), .B(n_203), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_367), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_367), .Y(n_398) );
INVx1_ASAP7_75t_SL g399 ( .A(n_365), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_377), .A2(n_339), .B(n_351), .Y(n_400) );
INVx1_ASAP7_75t_SL g401 ( .A(n_386), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_395), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_391), .A2(n_357), .B1(n_366), .B2(n_370), .C(n_363), .Y(n_403) );
NAND4xp75_ASAP7_75t_L g404 ( .A(n_396), .B(n_352), .C(n_338), .D(n_361), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_389), .B(n_366), .Y(n_405) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_383), .B(n_369), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_381), .B(n_359), .Y(n_407) );
CKINVDCx14_ASAP7_75t_R g408 ( .A(n_378), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_392), .A2(n_349), .B1(n_362), .B2(n_371), .C(n_355), .Y(n_409) );
XOR2x2_ASAP7_75t_L g410 ( .A(n_376), .B(n_371), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_379), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
XNOR2x1_ASAP7_75t_L g413 ( .A(n_394), .B(n_192), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_397), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_393), .B(n_399), .Y(n_415) );
NOR2x1p5_ASAP7_75t_L g416 ( .A(n_398), .B(n_192), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_382), .A2(n_155), .B1(n_131), .B2(n_134), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_384), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_414), .A2(n_374), .B1(n_380), .B2(n_375), .C(n_387), .Y(n_419) );
NAND2xp33_ASAP7_75t_SL g420 ( .A(n_415), .B(n_388), .Y(n_420) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_405), .A2(n_401), .B(n_406), .Y(n_421) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_410), .A2(n_382), .B(n_385), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_418), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_412), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_417), .B(n_390), .Y(n_425) );
AOI321xp33_ASAP7_75t_L g426 ( .A1(n_403), .A2(n_129), .A3(n_131), .B1(n_134), .B2(n_409), .C(n_407), .Y(n_426) );
AOI322xp5_ASAP7_75t_L g427 ( .A1(n_411), .A2(n_305), .A3(n_401), .B1(n_408), .B2(n_350), .C1(n_402), .C2(n_414), .Y(n_427) );
AND4x1_ASAP7_75t_L g428 ( .A(n_416), .B(n_393), .C(n_406), .D(n_396), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_413), .A2(n_305), .B1(n_400), .B2(n_410), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_406), .A2(n_396), .B(n_404), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_424), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_428), .B(n_425), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_421), .B(n_427), .Y(n_433) );
OAI221xp5_ASAP7_75t_SL g434 ( .A1(n_433), .A2(n_422), .B1(n_429), .B2(n_426), .C(n_419), .Y(n_434) );
NOR4xp25_ASAP7_75t_L g435 ( .A(n_433), .B(n_430), .C(n_429), .D(n_423), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_431), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_436), .B(n_432), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_434), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_437), .Y(n_439) );
OR3x2_ASAP7_75t_L g440 ( .A(n_439), .B(n_438), .C(n_435), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_440), .A2(n_432), .B(n_420), .Y(n_441) );
endmodule