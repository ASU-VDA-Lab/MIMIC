module fake_jpeg_7637_n_252 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_16),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_42),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_32),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_46),
.B(n_27),
.C(n_22),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

HAxp5_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_16),
.CON(n_46),
.SN(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_59),
.Y(n_86)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_51),
.B(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_56),
.A2(n_66),
.B1(n_67),
.B2(n_10),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_18),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_21),
.B1(n_23),
.B2(n_19),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_34),
.B1(n_30),
.B2(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_32),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_25),
.B1(n_24),
.B2(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_29),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_28),
.B1(n_34),
.B2(n_30),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_28),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_79),
.B(n_101),
.Y(n_126)
);

OR2x6_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_28),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_35),
.B(n_33),
.C(n_23),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_104),
.B1(n_75),
.B2(n_68),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_93),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_34),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_13),
.B1(n_14),
.B2(n_85),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_41),
.C(n_34),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_69),
.C(n_48),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_107),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_62),
.A2(n_30),
.B1(n_34),
.B2(n_2),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_50),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_11),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_109),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_11),
.B1(n_4),
.B2(n_6),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_0),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_76),
.B(n_8),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_12),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_114),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_57),
.B1(n_75),
.B2(n_69),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_116),
.A2(n_135),
.B1(n_107),
.B2(n_87),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_94),
.C(n_78),
.Y(n_141)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_122),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_109),
.Y(n_145)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_79),
.A2(n_54),
.B(n_53),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_133),
.B(n_108),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_108),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_15),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_15),
.B(n_8),
.C(n_9),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_134),
.B1(n_99),
.B2(n_85),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_6),
.B(n_12),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_129),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_139),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_140),
.B(n_142),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_161),
.C(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_146),
.B1(n_118),
.B2(n_131),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_148),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_78),
.B1(n_93),
.B2(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_157),
.B(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_128),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_77),
.B1(n_95),
.B2(n_90),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_135),
.B1(n_110),
.B2(n_127),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_150),
.C(n_141),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_123),
.B(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_90),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_168),
.C(n_170),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_174),
.C(n_156),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_166),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_126),
.C(n_110),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_127),
.B1(n_118),
.B2(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_131),
.B1(n_134),
.B2(n_110),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_111),
.B(n_124),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_157),
.B(n_137),
.Y(n_190)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_161),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_186),
.C(n_195),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_121),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_187),
.B(n_191),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_196),
.B1(n_180),
.B2(n_172),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_173),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_148),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_146),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_178),
.A2(n_142),
.B1(n_149),
.B2(n_143),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_122),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_198),
.Y(n_204)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_151),
.B(n_133),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_178),
.B1(n_169),
.B2(n_175),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_145),
.C(n_111),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_186),
.C(n_174),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_174),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_207),
.C(n_211),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_199),
.B(n_185),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_210),
.A2(n_196),
.B1(n_193),
.B2(n_200),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_183),
.C(n_182),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_168),
.B1(n_167),
.B2(n_183),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_212),
.A2(n_214),
.B(n_215),
.Y(n_218)
);

XNOR2x2_ASAP7_75t_SL g213 ( 
.A(n_189),
.B(n_181),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_190),
.B(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_167),
.B1(n_182),
.B2(n_179),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_176),
.B1(n_170),
.B2(n_177),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_222),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_220),
.B(n_226),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_200),
.B(n_188),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_224),
.B(n_199),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_195),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_176),
.C(n_191),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_225),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_165),
.C(n_163),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_206),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_219),
.A2(n_213),
.B(n_212),
.C(n_204),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_233),
.B1(n_217),
.B2(n_138),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_221),
.A2(n_208),
.B(n_203),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_232),
.B(n_229),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_215),
.B1(n_214),
.B2(n_203),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_120),
.Y(n_235)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

OAI221xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_225),
.B1(n_223),
.B2(n_211),
.C(n_217),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_240),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_228),
.A2(n_100),
.B1(n_83),
.B2(n_95),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_238),
.B(n_120),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_239),
.A2(n_234),
.B(n_231),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_222),
.C(n_205),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_14),
.B(n_105),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_237),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_243),
.CI(n_231),
.CON(n_245),
.SN(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

INVxp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_249),
.A2(n_247),
.B1(n_100),
.B2(n_83),
.Y(n_250)
);

AOI321xp33_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_88),
.A3(n_102),
.B1(n_105),
.B2(n_248),
.C(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_88),
.Y(n_252)
);


endmodule