module fake_jpeg_1088_n_426 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_1),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_54),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_51),
.B(n_82),
.Y(n_115)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_63),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_58),
.Y(n_133)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_61),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_65),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_1),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_17),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_25),
.B1(n_39),
.B2(n_31),
.Y(n_97)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_84),
.Y(n_138)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_4),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_24),
.B(n_14),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_5),
.Y(n_140)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_44),
.A2(n_17),
.B1(n_36),
.B2(n_41),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_92),
.A2(n_136),
.B1(n_49),
.B2(n_60),
.Y(n_156)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_99),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_97),
.A2(n_139),
.B1(n_37),
.B2(n_9),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_98),
.Y(n_149)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_65),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_74),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_114),
.B(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_132),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_27),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_36),
.C(n_40),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_71),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_66),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_122),
.B(n_6),
.Y(n_182)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_45),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_134),
.B(n_6),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_56),
.A2(n_30),
.B1(n_40),
.B2(n_22),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_72),
.A2(n_22),
.B1(n_16),
.B2(n_40),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_5),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_142),
.A2(n_191),
.B(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_67),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_143),
.B(n_158),
.Y(n_202)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_136),
.A2(n_69),
.B1(n_83),
.B2(n_79),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_145),
.A2(n_154),
.B1(n_156),
.B2(n_159),
.Y(n_204)
);

AOI32xp33_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_59),
.A3(n_47),
.B1(n_86),
.B2(n_46),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_153),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_78),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_92),
.A2(n_68),
.B1(n_55),
.B2(n_77),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_53),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_118),
.A2(n_103),
.B1(n_117),
.B2(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_103),
.B(n_22),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_176),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_165),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_89),
.Y(n_166)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_98),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_169),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_16),
.B1(n_37),
.B2(n_7),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_168),
.A2(n_175),
.B1(n_187),
.B2(n_14),
.Y(n_224)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_121),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_182),
.Y(n_220)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_70),
.B1(n_62),
.B2(n_16),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_174),
.A2(n_145),
.B(n_170),
.C(n_166),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_37),
.B1(n_9),
.B2(n_10),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_117),
.B(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_178),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_94),
.B(n_95),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_179),
.B(n_180),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_130),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

NAND2x1p5_ASAP7_75t_L g185 ( 
.A(n_107),
.B(n_37),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_96),
.B(n_6),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_12),
.Y(n_217)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_189),
.Y(n_225)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_91),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_104),
.B(n_9),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_104),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_113),
.B1(n_110),
.B2(n_105),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_200),
.B1(n_212),
.B2(n_214),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_113),
.B1(n_110),
.B2(n_105),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_126),
.B1(n_100),
.B2(n_96),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_155),
.B1(n_174),
.B2(n_192),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_142),
.B(n_126),
.C(n_90),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_206),
.C(n_235),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_142),
.B(n_90),
.C(n_100),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_37),
.B(n_11),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_232),
.B(n_174),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_160),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_141),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_217),
.B(n_212),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_143),
.B(n_13),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_236),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_184),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_163),
.A2(n_14),
.B(n_147),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_226),
.A2(n_229),
.B(n_199),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_157),
.A2(n_185),
.B(n_159),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_174),
.B1(n_189),
.B2(n_172),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_174),
.A2(n_152),
.B(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_148),
.B(n_162),
.C(n_171),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_149),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_239),
.A2(n_242),
.B1(n_249),
.B2(n_271),
.Y(n_307)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_240),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_152),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_270),
.C(n_228),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_177),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g302 ( 
.A(n_245),
.B(n_254),
.C(n_262),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_211),
.A2(n_144),
.B1(n_181),
.B2(n_188),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_247),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_193),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_250),
.B(n_267),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_150),
.B1(n_164),
.B2(n_161),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_178),
.B(n_153),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_258),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_198),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_206),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_255),
.B(n_259),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_203),
.Y(n_256)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_198),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_257),
.B(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_209),
.B(n_205),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_204),
.A2(n_193),
.B1(n_202),
.B2(n_232),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_213),
.B(n_220),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_204),
.A2(n_202),
.B1(n_234),
.B2(n_197),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_263),
.A2(n_269),
.B1(n_274),
.B2(n_222),
.Y(n_289)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_272),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_224),
.A2(n_230),
.B1(n_229),
.B2(n_221),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_266),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_223),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_216),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_220),
.B(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_227),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_235),
.B1(n_194),
.B2(n_195),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_196),
.B(n_195),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_194),
.A2(n_203),
.B1(n_225),
.B2(n_210),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_233),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_273),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_227),
.B1(n_228),
.B2(n_233),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_218),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_219),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_292),
.C(n_300),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_278),
.B(n_309),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_284),
.B(n_259),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_262),
.B(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_293),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_291),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_248),
.A2(n_237),
.B(n_222),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_287),
.A2(n_255),
.B(n_247),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_289),
.A2(n_306),
.B1(n_256),
.B2(n_273),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_274),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_238),
.B(n_237),
.C(n_199),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_266),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_275),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_296),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_245),
.B(n_257),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_238),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_271),
.Y(n_301)
);

INVx11_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_240),
.B(n_264),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

NOR2x1_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_249),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_305),
.A2(n_250),
.B(n_267),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_263),
.A2(n_244),
.B1(n_248),
.B2(n_242),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_260),
.Y(n_309)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g357 ( 
.A1(n_313),
.A2(n_326),
.B(n_332),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_251),
.B1(n_239),
.B2(n_253),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_333),
.B1(n_301),
.B2(n_283),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_314),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_325),
.Y(n_356)
);

NOR3xp33_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_254),
.C(n_276),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_334),
.C(n_335),
.Y(n_347)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_279),
.A2(n_255),
.B(n_259),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_255),
.C(n_259),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_329),
.C(n_299),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_304),
.Y(n_324)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_327),
.B(n_338),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_258),
.C(n_246),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_281),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_331),
.B(n_336),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_297),
.A2(n_261),
.B(n_251),
.Y(n_332)
);

OAI322xp33_ASAP7_75t_L g334 ( 
.A1(n_308),
.A2(n_256),
.A3(n_293),
.B1(n_296),
.B2(n_282),
.C1(n_295),
.C2(n_290),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_286),
.B(n_278),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_SL g336 ( 
.A(n_290),
.B(n_282),
.C(n_309),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_280),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_350),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_315),
.A2(n_306),
.B1(n_289),
.B2(n_283),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_340),
.A2(n_351),
.B1(n_361),
.B2(n_321),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_358),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_317),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_348),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_330),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_349),
.A2(n_355),
.B1(n_313),
.B2(n_328),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_284),
.C(n_299),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_318),
.A2(n_298),
.B1(n_285),
.B2(n_291),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_318),
.B(n_280),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_327),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_333),
.A2(n_279),
.B1(n_305),
.B2(n_287),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_316),
.B(n_322),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_337),
.A2(n_305),
.B1(n_281),
.B2(n_302),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_359),
.A2(n_326),
.B(n_320),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_311),
.B(n_277),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_329),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_328),
.A2(n_303),
.B1(n_310),
.B2(n_332),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_352),
.A2(n_331),
.B1(n_324),
.B2(n_321),
.Y(n_362)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_356),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_366),
.Y(n_386)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_364),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_365),
.A2(n_367),
.B1(n_361),
.B2(n_352),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_356),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_355),
.A2(n_323),
.B1(n_311),
.B2(n_335),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_377),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_357),
.A2(n_334),
.B(n_323),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_370),
.A2(n_371),
.B(n_373),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_372),
.A2(n_345),
.B1(n_347),
.B2(n_343),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_357),
.A2(n_336),
.B(n_321),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_375),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_358),
.B(n_325),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_380),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_338),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_350),
.C(n_339),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_340),
.A2(n_310),
.B1(n_312),
.B2(n_359),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_381),
.B(n_382),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_354),
.C(n_360),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_363),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_388),
.A2(n_366),
.B(n_367),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_390),
.B(n_393),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_391),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_376),
.C(n_379),
.Y(n_393)
);

AOI21xp33_ASAP7_75t_L g397 ( 
.A1(n_394),
.A2(n_371),
.B(n_365),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_373),
.A2(n_345),
.B(n_341),
.Y(n_395)
);

OAI21x1_ASAP7_75t_SL g400 ( 
.A1(n_395),
.A2(n_384),
.B(n_389),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_400),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_399),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_387),
.A2(n_370),
.B(n_380),
.Y(n_399)
);

OAI221xp5_ASAP7_75t_L g401 ( 
.A1(n_394),
.A2(n_377),
.B1(n_369),
.B2(n_376),
.C(n_343),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_404),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_310),
.C(n_381),
.Y(n_404)
);

NAND4xp25_ASAP7_75t_SL g405 ( 
.A(n_392),
.B(n_386),
.C(n_395),
.D(n_390),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_385),
.Y(n_407)
);

OAI21x1_ASAP7_75t_SL g406 ( 
.A1(n_392),
.A2(n_389),
.B(n_385),
.Y(n_406)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_406),
.A2(n_384),
.B(n_386),
.Y(n_411)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_407),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_404),
.B(n_382),
.C(n_383),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_402),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_383),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_410),
.A2(n_411),
.B(n_414),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_388),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_415),
.B(n_416),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_387),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_409),
.B(n_405),
.C(n_413),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_418),
.B(n_413),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_419),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_420),
.B(n_417),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_421),
.A2(n_418),
.B(n_412),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_L g425 ( 
.A1(n_423),
.A2(n_424),
.B(n_422),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_416),
.Y(n_426)
);


endmodule