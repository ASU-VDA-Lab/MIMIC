module fake_jpeg_8866_n_109 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_0),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_12),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_13),
.B1(n_27),
.B2(n_26),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_12),
.B1(n_24),
.B2(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_31),
.B(n_25),
.C(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_53),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_18),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_47),
.B(n_59),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_13),
.B1(n_18),
.B2(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_52),
.B1(n_21),
.B2(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_23),
.B1(n_16),
.B2(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_26),
.B(n_28),
.Y(n_60)
);

FAx1_ASAP7_75t_SL g59 ( 
.A(n_32),
.B(n_27),
.CI(n_26),
.CON(n_59),
.SN(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_59),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_46),
.B(n_59),
.C(n_51),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_28),
.B1(n_21),
.B2(n_4),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_47),
.B1(n_44),
.B2(n_58),
.Y(n_77)
);

AOI221xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_77),
.B1(n_78),
.B2(n_69),
.C(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_80),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_79),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_52),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_81),
.C(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_4),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_46),
.C(n_45),
.Y(n_81)
);

NOR2xp67_ASAP7_75t_R g82 ( 
.A(n_65),
.B(n_45),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_60),
.C(n_3),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.C(n_85),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_68),
.C(n_72),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_62),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_1),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_77),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_82),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_92),
.B(n_93),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_98),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_87),
.C(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_67),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_102),
.C(n_66),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_70),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_90),
.B(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_100),
.B(n_70),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_105),
.B1(n_66),
.B2(n_6),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_10),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_106),
.Y(n_109)
);


endmodule