module fake_jpeg_15291_n_61 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_61);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_61;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_9),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_5),
.B(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_1),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_41),
.C(n_42),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_3),
.B1(n_6),
.B2(n_11),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_3),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_20),
.B1(n_34),
.B2(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_27),
.B(n_25),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_50)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_49),
.A2(n_43),
.B1(n_38),
.B2(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_51),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_55),
.B(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_28),
.Y(n_61)
);


endmodule