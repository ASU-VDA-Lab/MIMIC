module fake_ibex_1011_n_1537 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_285, n_139, n_247, n_274, n_288, n_55, n_130, n_275, n_291, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_273, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_287, n_110, n_193, n_293, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_278, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_282, n_14, n_0, n_239, n_289, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_294, n_150, n_286, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_284, n_80, n_172, n_215, n_250, n_279, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_281, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_280, n_269, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_283, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_270, n_295, n_230, n_96, n_185, n_271, n_241, n_68, n_117, n_292, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_290, n_218, n_259, n_132, n_174, n_276, n_277, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_272, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1537);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_285;
input n_139;
input n_247;
input n_274;
input n_288;
input n_55;
input n_130;
input n_275;
input n_291;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_273;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_287;
input n_110;
input n_193;
input n_293;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_278;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_282;
input n_14;
input n_0;
input n_239;
input n_289;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_294;
input n_150;
input n_286;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_284;
input n_80;
input n_172;
input n_215;
input n_250;
input n_279;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_281;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_280;
input n_269;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_283;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_270;
input n_295;
input n_230;
input n_96;
input n_185;
input n_271;
input n_241;
input n_68;
input n_117;
input n_292;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_290;
input n_218;
input n_259;
input n_132;
input n_174;
input n_276;
input n_277;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_272;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1537;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_737;
wire n_606;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_303;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1433;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1397;
wire n_1211;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_143),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_2),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_167),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_65),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_175),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_120),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_223),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_99),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_75),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_237),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_239),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_26),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_62),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_200),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_233),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_125),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_280),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_71),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_184),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_236),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_135),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_193),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_248),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_85),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_88),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_27),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_232),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_59),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_1),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_6),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_285),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_9),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_165),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_85),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_32),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_172),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_36),
.B(n_0),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_61),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_269),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_137),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_43),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_39),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_189),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_244),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_88),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_163),
.B(n_99),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_152),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_204),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_194),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_93),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_192),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_131),
.B(n_262),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_201),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_207),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_162),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_141),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_268),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_29),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_15),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_156),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_190),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_1),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_159),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_82),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_139),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_33),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_47),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_263),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_155),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_27),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_153),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_46),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_33),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_35),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_118),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_4),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_45),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_272),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_294),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_56),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_206),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_6),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_238),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_235),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_78),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_75),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_73),
.B(n_116),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_28),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_29),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_183),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_72),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_158),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_256),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_253),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_126),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_250),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_19),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_164),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_59),
.Y(n_398)
);

INVxp33_ASAP7_75t_SL g399 ( 
.A(n_259),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_170),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_291),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_279),
.B(n_276),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_21),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_74),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_95),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_282),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_46),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_81),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_78),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_0),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_71),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_264),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_103),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_129),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_258),
.B(n_187),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_278),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_275),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_185),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_68),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_246),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_83),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_171),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_195),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_142),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_295),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_149),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_147),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_229),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_224),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_179),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_289),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_69),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_28),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_178),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_4),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_260),
.Y(n_436)
);

BUFx10_ASAP7_75t_L g437 ( 
.A(n_254),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_242),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_114),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_128),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_181),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_261),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_136),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_102),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_182),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_271),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_226),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_130),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_231),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_227),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_210),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_157),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_120),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_252),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_110),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_216),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_288),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_98),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_2),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_150),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_205),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_198),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_73),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_188),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_191),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_292),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_106),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_274),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_95),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_211),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_251),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_199),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_42),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_31),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_217),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_160),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_86),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_17),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_202),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_80),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_70),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_283),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_257),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_208),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_108),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_9),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_203),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_270),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_117),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_115),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_293),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_39),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_19),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_47),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_70),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_255),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_105),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_290),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_146),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_45),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_54),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_118),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_186),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_213),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_301),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_301),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_350),
.A2(n_428),
.B(n_353),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_302),
.B(n_394),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_353),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_302),
.B(n_394),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_306),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_297),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_461),
.A2(n_127),
.B(n_124),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_461),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_319),
.Y(n_516)
);

BUFx12f_ASAP7_75t_L g517 ( 
.A(n_437),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_323),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_297),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_297),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_390),
.B(n_3),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_297),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_323),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_328),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_337),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_328),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_333),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_333),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_363),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_388),
.A2(n_7),
.B1(n_3),
.B2(n_5),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_409),
.B(n_7),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_328),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_421),
.B(n_8),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_328),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_336),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_336),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_466),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_363),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_437),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_336),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_390),
.B(n_10),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_406),
.B(n_10),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_336),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_309),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_418),
.B(n_427),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_307),
.B(n_11),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_490),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_365),
.B(n_11),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_359),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_468),
.B(n_12),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_309),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_359),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_359),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_365),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_359),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_304),
.B(n_12),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_362),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_366),
.Y(n_561)
);

CKINVDCx6p67_ASAP7_75t_R g562 ( 
.A(n_504),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_366),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_487),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_490),
.B(n_13),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_371),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_320),
.B(n_13),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_371),
.B(n_14),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_487),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_503),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_362),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_382),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_382),
.Y(n_577)
);

CKINVDCx6p67_ASAP7_75t_R g578 ( 
.A(n_391),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_391),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_392),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_417),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_444),
.B(n_459),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_396),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_417),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_438),
.Y(n_585)
);

BUFx8_ASAP7_75t_L g586 ( 
.A(n_351),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_438),
.B(n_132),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_465),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_308),
.A2(n_134),
.B(n_133),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_465),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_459),
.B(n_16),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_327),
.B(n_18),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_498),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_347),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_311),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_298),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_298),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_485),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_322),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_316),
.B(n_318),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_485),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_324),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_329),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_331),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_309),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_334),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_338),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_339),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_521),
.B(n_342),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_524),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_608),
.B(n_356),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_551),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_541),
.B(n_313),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_608),
.B(n_360),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g616 ( 
.A(n_568),
.B(n_335),
.Y(n_616)
);

AND2x6_ASAP7_75t_L g617 ( 
.A(n_521),
.B(n_367),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_551),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_551),
.A2(n_570),
.B1(n_605),
.B2(n_596),
.Y(n_619)
);

AND3x2_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_494),
.C(n_385),
.Y(n_620)
);

AND3x2_ASAP7_75t_L g621 ( 
.A(n_574),
.B(n_473),
.C(n_358),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_575),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_551),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_574),
.Y(n_625)
);

NOR2x1p5_ASAP7_75t_L g626 ( 
.A(n_517),
.B(n_326),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_508),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_516),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_575),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_546),
.B(n_420),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_591),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_521),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_597),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_591),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_550),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_576),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_562),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_521),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_543),
.Y(n_639)
);

BUFx6f_ASAP7_75t_SL g640 ( 
.A(n_543),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_576),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_548),
.B(n_330),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_510),
.B(n_330),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_R g644 ( 
.A(n_562),
.B(n_347),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_543),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_576),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_576),
.Y(n_647)
);

OAI21xp33_ASAP7_75t_SL g648 ( 
.A1(n_603),
.A2(n_303),
.B(n_300),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_594),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_597),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_526),
.B(n_332),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_543),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g653 ( 
.A(n_600),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_577),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_582),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_582),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_577),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_603),
.B(n_332),
.Y(n_660)
);

BUFx10_ASAP7_75t_L g661 ( 
.A(n_512),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_582),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_604),
.B(n_484),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_516),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_564),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_524),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_531),
.A2(n_354),
.B1(n_423),
.B2(n_355),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_524),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_577),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_560),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_564),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_532),
.B(n_474),
.C(n_469),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_517),
.B(n_469),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_608),
.B(n_368),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_604),
.B(n_370),
.Y(n_675)
);

BUFx8_ASAP7_75t_SL g676 ( 
.A(n_549),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_607),
.B(n_377),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_577),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_584),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_607),
.B(n_474),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_584),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_578),
.B(n_477),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_578),
.B(n_378),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_608),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_608),
.B(n_380),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_532),
.B(n_478),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_608),
.B(n_383),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_569),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_549),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_596),
.A2(n_310),
.B1(n_321),
.B2(n_315),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_531),
.A2(n_398),
.B1(n_435),
.B2(n_396),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_569),
.Y(n_692)
);

AO22x2_ASAP7_75t_L g693 ( 
.A1(n_598),
.A2(n_340),
.B1(n_341),
.B2(n_325),
.Y(n_693)
);

OR2x4_ASAP7_75t_L g694 ( 
.A(n_601),
.B(n_344),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_585),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_585),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_586),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_585),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_509),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_583),
.B(n_386),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_509),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_511),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_524),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

AND2x2_ASAP7_75t_SL g705 ( 
.A(n_534),
.B(n_415),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_511),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_507),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_553),
.B(n_478),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_586),
.B(n_489),
.C(n_486),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_553),
.B(n_502),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_609),
.B(n_389),
.Y(n_711)
);

AND3x2_ASAP7_75t_L g712 ( 
.A(n_583),
.B(n_357),
.C(n_349),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_605),
.B(n_393),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_586),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_515),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_605),
.B(n_505),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_581),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_525),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_525),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_538),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_507),
.A2(n_373),
.B1(n_374),
.B2(n_372),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_538),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_540),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_505),
.B(n_395),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_565),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_581),
.Y(n_726)
);

OAI21xp33_ASAP7_75t_SL g727 ( 
.A1(n_514),
.A2(n_404),
.B(n_384),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_609),
.B(n_397),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_593),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_544),
.B(n_592),
.C(n_559),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_593),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_527),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_593),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_507),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_507),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_565),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_609),
.B(n_400),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_589),
.B(n_405),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_609),
.B(n_401),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_506),
.B(n_518),
.Y(n_740)
);

INVx5_ASAP7_75t_L g741 ( 
.A(n_587),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_572),
.Y(n_742)
);

BUFx2_ASAP7_75t_L g743 ( 
.A(n_579),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_579),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_572),
.Y(n_745)
);

CKINVDCx11_ASAP7_75t_R g746 ( 
.A(n_609),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_573),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_527),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_619),
.A2(n_528),
.B1(n_529),
.B2(n_523),
.C(n_518),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_654),
.B(n_296),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_642),
.B(n_296),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_635),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_627),
.B(n_399),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_660),
.B(n_299),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_680),
.B(n_312),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_650),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_628),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_657),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_734),
.A2(n_514),
.B(n_589),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_614),
.B(n_314),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_661),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_644),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_630),
.B(n_317),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_658),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_640),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_630),
.B(n_317),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_653),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_664),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_692),
.B(n_493),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_662),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_651),
.B(n_493),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_631),
.B(n_472),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_653),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_688),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_610),
.A2(n_587),
.B1(n_573),
.B2(n_580),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_634),
.B(n_472),
.Y(n_776)
);

INVx8_ASAP7_75t_L g777 ( 
.A(n_640),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_743),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_663),
.B(n_475),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_670),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_740),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_714),
.B(n_413),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_730),
.B(n_479),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_623),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_623),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_744),
.B(n_482),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_716),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_686),
.B(n_495),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_716),
.Y(n_789)
);

BUFx4_ASAP7_75t_L g790 ( 
.A(n_682),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_643),
.B(n_496),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_699),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_701),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_702),
.Y(n_794)
);

NOR2x1p5_ASAP7_75t_L g795 ( 
.A(n_637),
.B(n_495),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_672),
.B(n_502),
.C(n_501),
.Y(n_796)
);

OAI22x1_ASAP7_75t_SL g797 ( 
.A1(n_649),
.A2(n_453),
.B1(n_450),
.B2(n_447),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_707),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_633),
.B(n_523),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_708),
.B(n_501),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_706),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_715),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_707),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_710),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_610),
.A2(n_588),
.B1(n_590),
.B2(n_580),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_705),
.B(n_588),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_683),
.B(n_528),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_683),
.B(n_529),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_746),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_694),
.B(n_530),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_639),
.A2(n_595),
.B(n_539),
.C(n_557),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_694),
.B(n_613),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_718),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_610),
.A2(n_617),
.B1(n_624),
.B2(n_618),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_617),
.A2(n_557),
.B1(n_561),
.B2(n_539),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_617),
.A2(n_563),
.B1(n_567),
.B2(n_561),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_719),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_673),
.B(n_305),
.Y(n_819)
);

AOI221x1_ASAP7_75t_L g820 ( 
.A1(n_652),
.A2(n_424),
.B1(n_426),
.B2(n_422),
.C(n_416),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_632),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_720),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_722),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_620),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_709),
.B(n_447),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_675),
.B(n_571),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_721),
.A2(n_602),
.B1(n_599),
.B2(n_439),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_675),
.B(n_599),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_697),
.A2(n_457),
.B1(n_470),
.B2(n_450),
.Y(n_829)
);

AND2x6_ASAP7_75t_SL g830 ( 
.A(n_700),
.B(n_419),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_741),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_677),
.B(n_343),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_625),
.B(n_361),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_638),
.B(n_346),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_638),
.B(n_348),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_645),
.B(n_352),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_645),
.B(n_648),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_723),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_676),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_724),
.B(n_431),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_725),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_616),
.A2(n_470),
.B1(n_499),
.B2(n_457),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_713),
.B(n_690),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_724),
.B(n_434),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_736),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_742),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_735),
.A2(n_458),
.B1(n_480),
.B2(n_455),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_735),
.A2(n_492),
.B1(n_497),
.B2(n_481),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_738),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_690),
.B(n_364),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_745),
.B(n_747),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_616),
.B(n_621),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_665),
.Y(n_853)
);

BUFx5_ASAP7_75t_L g854 ( 
.A(n_671),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_616),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_727),
.B(n_412),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_620),
.B(n_414),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_717),
.B(n_425),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_726),
.B(n_429),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_684),
.Y(n_860)
);

OR2x6_ASAP7_75t_L g861 ( 
.A(n_626),
.B(n_500),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_693),
.A2(n_499),
.B1(n_369),
.B2(n_376),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_667),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_612),
.B(n_430),
.Y(n_864)
);

BUFx6f_ASAP7_75t_SL g865 ( 
.A(n_700),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_615),
.B(n_436),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_615),
.B(n_445),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_738),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_674),
.B(n_462),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_685),
.B(n_581),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_687),
.B(n_440),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_693),
.A2(n_375),
.B1(n_381),
.B2(n_379),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_687),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_711),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_728),
.B(n_581),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_693),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_700),
.A2(n_403),
.B1(n_407),
.B2(n_387),
.Y(n_877)
);

INVx8_ASAP7_75t_L g878 ( 
.A(n_611),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_728),
.A2(n_441),
.B(n_443),
.C(n_442),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_737),
.B(n_446),
.Y(n_880)
);

BUFx6f_ASAP7_75t_SL g881 ( 
.A(n_691),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_712),
.B(n_408),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_739),
.A2(n_449),
.B1(n_451),
.B2(n_448),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_712),
.B(n_410),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_691),
.A2(n_432),
.B1(n_433),
.B2(n_411),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_739),
.B(n_581),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_622),
.B(n_345),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_629),
.B(n_452),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_636),
.B(n_454),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_641),
.A2(n_463),
.B(n_456),
.C(n_460),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_641),
.B(n_471),
.Y(n_891)
);

INVx8_ASAP7_75t_L g892 ( 
.A(n_611),
.Y(n_892)
);

OAI221xp5_ASAP7_75t_L g893 ( 
.A1(n_646),
.A2(n_467),
.B1(n_488),
.B2(n_491),
.C(n_476),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_646),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_647),
.B(n_547),
.Y(n_895)
);

OAI22xp33_ASAP7_75t_L g896 ( 
.A1(n_655),
.A2(n_547),
.B1(n_554),
.B2(n_402),
.Y(n_896)
);

NOR3xp33_ASAP7_75t_L g897 ( 
.A(n_655),
.B(n_554),
.C(n_547),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_656),
.B(n_547),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_656),
.B(n_554),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_659),
.B(n_554),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_669),
.B(n_22),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_813),
.B(n_22),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_798),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_853),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_843),
.A2(n_519),
.B1(n_520),
.B2(n_513),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_761),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_805),
.B(n_23),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_765),
.B(n_542),
.Y(n_908)
);

AOI22x1_ASAP7_75t_L g909 ( 
.A1(n_759),
.A2(n_679),
.B1(n_681),
.B2(n_678),
.Y(n_909)
);

CKINVDCx10_ASAP7_75t_R g910 ( 
.A(n_865),
.Y(n_910)
);

CKINVDCx10_ASAP7_75t_R g911 ( 
.A(n_865),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_846),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_853),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_813),
.B(n_24),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_774),
.B(n_24),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_788),
.A2(n_774),
.B1(n_782),
.B2(n_753),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_837),
.A2(n_696),
.B(n_698),
.C(n_695),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_771),
.B(n_25),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_808),
.B(n_809),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_811),
.B(n_25),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_811),
.B(n_26),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_756),
.Y(n_922)
);

OA22x2_ASAP7_75t_L g923 ( 
.A1(n_876),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_837),
.A2(n_731),
.B(n_733),
.C(n_729),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_750),
.B(n_30),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_807),
.B(n_34),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_L g927 ( 
.A1(n_876),
.A2(n_863),
.B1(n_783),
.B2(n_893),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_781),
.B(n_34),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_834),
.A2(n_836),
.B(n_835),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_799),
.Y(n_930)
);

OA22x2_ASAP7_75t_L g931 ( 
.A1(n_862),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_801),
.B(n_38),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_L g933 ( 
.A(n_885),
.B(n_872),
.C(n_877),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_R g934 ( 
.A(n_767),
.B(n_40),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_787),
.B(n_40),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_789),
.B(n_41),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_751),
.B(n_41),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_782),
.A2(n_522),
.B1(n_533),
.B2(n_513),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_784),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_855),
.B(n_42),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_815),
.A2(n_533),
.B1(n_536),
.B2(n_522),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_754),
.B(n_43),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_854),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_749),
.A2(n_533),
.B(n_536),
.C(n_545),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_755),
.B(n_44),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_810),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_749),
.A2(n_536),
.B(n_545),
.C(n_555),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_855),
.B(n_44),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_773),
.B(n_48),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_760),
.B(n_763),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_815),
.A2(n_555),
.B1(n_556),
.B2(n_606),
.Y(n_951)
);

OAI321xp33_ASAP7_75t_L g952 ( 
.A1(n_893),
.A2(n_606),
.A3(n_556),
.B1(n_537),
.B2(n_552),
.C(n_535),
.Y(n_952)
);

AO21x1_ASAP7_75t_L g953 ( 
.A1(n_890),
.A2(n_896),
.B(n_844),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_819),
.B(n_49),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_766),
.B(n_800),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_840),
.B(n_50),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_825),
.A2(n_542),
.B1(n_606),
.B2(n_537),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_840),
.B(n_50),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_765),
.B(n_51),
.Y(n_959)
);

NOR2x1p5_ASAP7_75t_SL g960 ( 
.A(n_854),
.B(n_138),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_844),
.A2(n_785),
.B(n_871),
.C(n_866),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_769),
.B(n_51),
.Y(n_962)
);

XOR2xp5_ASAP7_75t_L g963 ( 
.A(n_797),
.B(n_52),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_778),
.B(n_52),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_839),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_847),
.A2(n_848),
.B1(n_827),
.B2(n_816),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_779),
.B(n_53),
.Y(n_967)
);

BUFx6f_ASAP7_75t_SL g968 ( 
.A(n_824),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_791),
.B(n_54),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_827),
.A2(n_820),
.B(n_812),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_775),
.A2(n_668),
.B(n_666),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_829),
.B(n_55),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_772),
.B(n_57),
.Y(n_973)
);

BUFx12f_ASAP7_75t_L g974 ( 
.A(n_861),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_866),
.A2(n_527),
.B(n_535),
.C(n_537),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_871),
.A2(n_535),
.B(n_537),
.C(n_552),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_804),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_777),
.Y(n_978)
);

NOR2x1_ASAP7_75t_R g979 ( 
.A(n_881),
.B(n_58),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_821),
.Y(n_980)
);

BUFx4f_ASAP7_75t_L g981 ( 
.A(n_777),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_842),
.B(n_833),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_901),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_752),
.Y(n_984)
);

AOI221xp5_ASAP7_75t_L g985 ( 
.A1(n_881),
.A2(n_558),
.B1(n_732),
.B2(n_704),
.C(n_703),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_882),
.A2(n_558),
.B1(n_732),
.B2(n_704),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_776),
.B(n_58),
.Y(n_987)
);

OR2x6_ASAP7_75t_SL g988 ( 
.A(n_777),
.B(n_60),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_848),
.A2(n_558),
.B1(n_748),
.B2(n_732),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_786),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_816),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_758),
.B(n_63),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_796),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_851),
.A2(n_144),
.B(n_140),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_890),
.A2(n_64),
.B(n_66),
.C(n_67),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_764),
.B(n_66),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_873),
.A2(n_148),
.B(n_145),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_770),
.B(n_69),
.Y(n_998)
);

BUFx8_ASAP7_75t_L g999 ( 
.A(n_884),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_874),
.A2(n_154),
.B(n_151),
.Y(n_1000)
);

CKINVDCx10_ASAP7_75t_R g1001 ( 
.A(n_861),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_SL g1002 ( 
.A(n_849),
.B(n_161),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_762),
.B(n_74),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_817),
.B(n_76),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_880),
.A2(n_76),
.B(n_77),
.C(n_79),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_817),
.A2(n_879),
.B(n_806),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_850),
.A2(n_84),
.B(n_86),
.C(n_87),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_832),
.B(n_87),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_861),
.B(n_89),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_792),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_794),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_826),
.B(n_89),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_828),
.B(n_90),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_857),
.B(n_90),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_802),
.Y(n_1015)
);

BUFx2_ASAP7_75t_SL g1016 ( 
.A(n_868),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_852),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_803),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_1018)
);

OR2x6_ASAP7_75t_L g1019 ( 
.A(n_795),
.B(n_96),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_757),
.A2(n_214),
.B(n_287),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_880),
.A2(n_97),
.B(n_98),
.C(n_100),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_877),
.B(n_97),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_793),
.B(n_100),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_814),
.B(n_101),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_822),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_838),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_1026)
);

AO22x1_ASAP7_75t_L g1027 ( 
.A1(n_830),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_841),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_858),
.B(n_109),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_870),
.A2(n_221),
.B(n_281),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_818),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_845),
.B(n_111),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_823),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_875),
.A2(n_220),
.B(n_277),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_883),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_859),
.B(n_113),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_887),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_891),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_790),
.B(n_119),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_864),
.B(n_121),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_867),
.B(n_122),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_891),
.Y(n_1042)
);

AOI221xp5_ASAP7_75t_L g1043 ( 
.A1(n_869),
.A2(n_122),
.B1(n_123),
.B2(n_166),
.C(n_168),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_768),
.A2(n_230),
.B(n_169),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_887),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_780),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_886),
.A2(n_177),
.B(n_180),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_831),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_888),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_895),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_897),
.B(n_196),
.C(n_197),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_878),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_831),
.Y(n_1053)
);

BUFx12f_ASAP7_75t_L g1054 ( 
.A(n_889),
.Y(n_1054)
);

NOR4xp25_ASAP7_75t_L g1055 ( 
.A(n_1018),
.B(n_898),
.C(n_900),
.D(n_894),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_903),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_SL g1057 ( 
.A1(n_916),
.A2(n_897),
.B(n_899),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_922),
.B(n_860),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_SL g1059 ( 
.A1(n_917),
.A2(n_892),
.B(n_212),
.C(n_215),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_927),
.B(n_892),
.Y(n_1060)
);

AOI221xp5_ASAP7_75t_L g1061 ( 
.A1(n_933),
.A2(n_209),
.B1(n_218),
.B2(n_219),
.C(n_222),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_SL g1062 ( 
.A1(n_1003),
.A2(n_225),
.B(n_228),
.C(n_234),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_972),
.B(n_906),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_961),
.A2(n_240),
.B(n_243),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_1009),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_904),
.B(n_913),
.Y(n_1066)
);

AO31x2_ASAP7_75t_L g1067 ( 
.A1(n_924),
.A2(n_245),
.A3(n_247),
.B(n_249),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_1052),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_981),
.Y(n_1069)
);

OA21x2_ASAP7_75t_L g1070 ( 
.A1(n_971),
.A2(n_265),
.B(n_266),
.Y(n_1070)
);

NOR2x1_ASAP7_75t_L g1071 ( 
.A(n_1009),
.B(n_267),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1010),
.Y(n_1072)
);

BUFx4f_ASAP7_75t_L g1073 ( 
.A(n_1009),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_943),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_959),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_974),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_912),
.B(n_273),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_970),
.A2(n_971),
.B(n_1006),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1011),
.B(n_1015),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1025),
.B(n_962),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_907),
.B(n_990),
.Y(n_1081)
);

CKINVDCx11_ASAP7_75t_R g1082 ( 
.A(n_965),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_981),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_946),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_966),
.A2(n_983),
.B1(n_956),
.B2(n_958),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_1001),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_1040),
.A2(n_1038),
.B(n_1042),
.C(n_918),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_954),
.B(n_932),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_982),
.B(n_978),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_910),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1033),
.B(n_964),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_928),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_915),
.B(n_920),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_921),
.B(n_1050),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_1019),
.B(n_1016),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_1019),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_902),
.B(n_914),
.Y(n_1097)
);

NOR4xp25_ASAP7_75t_L g1098 ( 
.A(n_1018),
.B(n_1037),
.C(n_1026),
.D(n_995),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_935),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_939),
.B(n_936),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_940),
.B(n_948),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1012),
.B(n_1013),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_952),
.A2(n_1044),
.B(n_976),
.Y(n_1103)
);

OAI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1019),
.A2(n_988),
.B1(n_931),
.B2(n_923),
.Y(n_1104)
);

INVx1_ASAP7_75t_SL g1105 ( 
.A(n_943),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_953),
.A2(n_905),
.A3(n_989),
.B(n_975),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1022),
.B(n_1031),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1024),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_926),
.B(n_925),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1006),
.A2(n_947),
.B(n_944),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_911),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_934),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_930),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1023),
.B(n_973),
.Y(n_1114)
);

BUFx4f_ASAP7_75t_L g1115 ( 
.A(n_959),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1039),
.B(n_1045),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_1048),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_999),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_987),
.B(n_967),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1032),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_937),
.A2(n_969),
.B(n_942),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_951),
.A2(n_998),
.B(n_992),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_996),
.A2(n_1004),
.B(n_945),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_1005),
.A2(n_1021),
.A3(n_991),
.B(n_941),
.Y(n_1124)
);

AO21x2_ASAP7_75t_L g1125 ( 
.A1(n_1008),
.A2(n_1051),
.B(n_1041),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_994),
.A2(n_997),
.A3(n_1000),
.B(n_1035),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_968),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_949),
.B(n_1014),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1029),
.B(n_1036),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1020),
.A2(n_1030),
.A3(n_1034),
.B(n_1047),
.Y(n_1130)
);

AOI31xp67_ASAP7_75t_L g1131 ( 
.A1(n_1046),
.A2(n_923),
.A3(n_960),
.B(n_986),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_1054),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1007),
.A2(n_1028),
.B(n_993),
.C(n_1043),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_931),
.B(n_1027),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_980),
.B(n_1048),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1049),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_977),
.B(n_1053),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1053),
.B(n_957),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_968),
.B(n_979),
.Y(n_1139)
);

CKINVDCx16_ASAP7_75t_R g1140 ( 
.A(n_963),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_SL g1141 ( 
.A1(n_1017),
.A2(n_938),
.B(n_985),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_999),
.B(n_908),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_933),
.A2(n_919),
.B1(n_966),
.B2(n_927),
.Y(n_1143)
);

AOI221x1_ASAP7_75t_L g1144 ( 
.A1(n_971),
.A2(n_1037),
.B1(n_970),
.B2(n_917),
.C(n_924),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_922),
.B(n_761),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_906),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_906),
.B(n_904),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_984),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_933),
.A2(n_919),
.B1(n_966),
.B2(n_927),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_919),
.B(n_927),
.Y(n_1150)
);

INVxp67_ASAP7_75t_SL g1151 ( 
.A(n_903),
.Y(n_1151)
);

AO221x2_ASAP7_75t_L g1152 ( 
.A1(n_963),
.A2(n_583),
.B1(n_1018),
.B2(n_1037),
.C(n_1027),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_906),
.B(n_904),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_919),
.B(n_927),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1052),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_950),
.A2(n_837),
.B(n_929),
.C(n_961),
.Y(n_1156)
);

NOR3xp33_ASAP7_75t_L g1157 ( 
.A(n_979),
.B(n_1027),
.C(n_933),
.Y(n_1157)
);

NAND2xp33_ASAP7_75t_L g1158 ( 
.A(n_943),
.B(n_799),
.Y(n_1158)
);

AOI21xp33_ASAP7_75t_SL g1159 ( 
.A1(n_963),
.A2(n_797),
.B(n_691),
.Y(n_1159)
);

NOR4xp25_ASAP7_75t_L g1160 ( 
.A(n_1018),
.B(n_1037),
.C(n_1026),
.D(n_995),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_961),
.A2(n_727),
.B(n_759),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_950),
.A2(n_837),
.B(n_929),
.C(n_961),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_903),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_903),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_933),
.B(n_1043),
.C(n_1007),
.Y(n_1165)
);

AO221x2_ASAP7_75t_L g1166 ( 
.A1(n_963),
.A2(n_583),
.B1(n_1018),
.B2(n_1037),
.C(n_1027),
.Y(n_1166)
);

BUFx4_ASAP7_75t_SL g1167 ( 
.A(n_1009),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_950),
.A2(n_837),
.B(n_929),
.C(n_961),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_984),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_961),
.A2(n_727),
.B(n_759),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_906),
.Y(n_1171)
);

AO21x1_ASAP7_75t_L g1172 ( 
.A1(n_1002),
.A2(n_1044),
.B(n_856),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_919),
.A2(n_966),
.B1(n_983),
.B2(n_619),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_903),
.Y(n_1174)
);

BUFx10_ASAP7_75t_L g1175 ( 
.A(n_1009),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_950),
.A2(n_837),
.B(n_929),
.C(n_961),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_971),
.A2(n_759),
.B(n_909),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_919),
.A2(n_955),
.B(n_950),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_961),
.A2(n_727),
.B(n_759),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_917),
.A2(n_924),
.A3(n_953),
.B(n_905),
.Y(n_1180)
);

NOR4xp25_ASAP7_75t_L g1181 ( 
.A(n_1018),
.B(n_1037),
.C(n_1026),
.D(n_995),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_984),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_922),
.B(n_761),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_922),
.B(n_761),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_917),
.A2(n_924),
.A3(n_953),
.B(n_905),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_984),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_919),
.B(n_927),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_933),
.A2(n_881),
.B1(n_863),
.B2(n_876),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_SL g1189 ( 
.A(n_965),
.Y(n_1189)
);

NAND3x1_ASAP7_75t_L g1190 ( 
.A(n_933),
.B(n_842),
.C(n_531),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_984),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_919),
.A2(n_966),
.B1(n_983),
.B2(n_782),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_903),
.B(n_689),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_919),
.B(n_927),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_903),
.B(n_689),
.Y(n_1195)
);

AOI221x1_ASAP7_75t_L g1196 ( 
.A1(n_971),
.A2(n_1037),
.B1(n_970),
.B2(n_917),
.C(n_924),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_917),
.A2(n_924),
.A3(n_953),
.B(n_905),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_984),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_974),
.B(n_767),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_982),
.B(n_863),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_919),
.B(n_927),
.Y(n_1201)
);

BUFx10_ASAP7_75t_L g1202 ( 
.A(n_1009),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_917),
.A2(n_924),
.A3(n_953),
.B(n_905),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1156),
.A2(n_1168),
.B(n_1162),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1095),
.B(n_1167),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1066),
.Y(n_1206)
);

CKINVDCx8_ASAP7_75t_R g1207 ( 
.A(n_1090),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1200),
.B(n_1193),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1095),
.B(n_1096),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1195),
.B(n_1073),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1078),
.A2(n_1170),
.B(n_1161),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_1068),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1182),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1144),
.A2(n_1196),
.A3(n_1172),
.B(n_1085),
.Y(n_1215)
);

BUFx8_ASAP7_75t_L g1216 ( 
.A(n_1086),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1073),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1186),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1178),
.B(n_1089),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1189),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1115),
.B(n_1155),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1072),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1069),
.B(n_1199),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1148),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1150),
.B(n_1154),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1083),
.B(n_1065),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1121),
.A2(n_1176),
.B(n_1179),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1063),
.B(n_1152),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_SL g1229 ( 
.A1(n_1192),
.A2(n_1071),
.B(n_1064),
.Y(n_1229)
);

BUFx2_ASAP7_75t_R g1230 ( 
.A(n_1118),
.Y(n_1230)
);

AOI221xp5_ASAP7_75t_L g1231 ( 
.A1(n_1159),
.A2(n_1104),
.B1(n_1173),
.B2(n_1201),
.C(n_1187),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1147),
.B(n_1153),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1097),
.A2(n_1177),
.B(n_1087),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1194),
.B(n_1143),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1143),
.B(n_1149),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1102),
.A2(n_1109),
.B(n_1119),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1188),
.B(n_1081),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1149),
.A2(n_1085),
.B(n_1110),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1191),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1173),
.B(n_1198),
.Y(n_1240)
);

BUFx12f_ASAP7_75t_L g1241 ( 
.A(n_1082),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1084),
.B(n_1132),
.Y(n_1242)
);

OR2x2_ASAP7_75t_L g1243 ( 
.A(n_1056),
.B(n_1163),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1079),
.B(n_1099),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1105),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1136),
.Y(n_1246)
);

OAI21xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1074),
.A2(n_1105),
.B(n_1134),
.Y(n_1247)
);

AOI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1103),
.A2(n_1070),
.B(n_1093),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1152),
.B(n_1166),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1174),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1113),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1146),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1166),
.B(n_1151),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1165),
.A2(n_1190),
.B1(n_1080),
.B2(n_1088),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1165),
.A2(n_1133),
.B(n_1110),
.C(n_1123),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1129),
.B(n_1101),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1137),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1122),
.A2(n_1125),
.B(n_1059),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1108),
.B(n_1120),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1125),
.A2(n_1114),
.B(n_1100),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1058),
.Y(n_1261)
);

AOI21xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1111),
.A2(n_1157),
.B(n_1140),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1077),
.B(n_1171),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1077),
.B(n_1092),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1117),
.A2(n_1141),
.B(n_1060),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1061),
.A2(n_1057),
.B(n_1107),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1055),
.A2(n_1131),
.B(n_1094),
.Y(n_1267)
);

AO21x2_ASAP7_75t_L g1268 ( 
.A1(n_1062),
.A2(n_1098),
.B(n_1181),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1057),
.A2(n_1138),
.B(n_1091),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1128),
.A2(n_1130),
.B(n_1158),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1124),
.B(n_1181),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1138),
.A2(n_1203),
.B(n_1197),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1175),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1112),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1202),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1098),
.A2(n_1160),
.B(n_1135),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1106),
.A2(n_1203),
.B(n_1197),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1164),
.B(n_1075),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1160),
.A2(n_1142),
.B1(n_1202),
.B2(n_1145),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1183),
.A2(n_1184),
.B(n_1116),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1124),
.B(n_1197),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1106),
.A2(n_1203),
.B(n_1185),
.Y(n_1282)
);

CKINVDCx14_ASAP7_75t_R g1283 ( 
.A(n_1076),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1075),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1180),
.A2(n_1067),
.B(n_1126),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1127),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1067),
.B(n_1139),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1082),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1169),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1144),
.A2(n_1196),
.A3(n_1172),
.B(n_1085),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1073),
.B(n_1115),
.Y(n_1291)
);

OR2x6_ASAP7_75t_L g1292 ( 
.A(n_1095),
.B(n_1009),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1193),
.B(n_903),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1156),
.A2(n_1168),
.B(n_1162),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1105),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1240),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1289),
.B(n_1276),
.Y(n_1297)
);

BUFx8_ASAP7_75t_L g1298 ( 
.A(n_1241),
.Y(n_1298)
);

BUFx2_ASAP7_75t_SL g1299 ( 
.A(n_1213),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1213),
.Y(n_1300)
);

AO21x2_ASAP7_75t_L g1301 ( 
.A1(n_1258),
.A2(n_1267),
.B(n_1204),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1235),
.B(n_1271),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1256),
.B(n_1206),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1221),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1231),
.A2(n_1249),
.B1(n_1237),
.B2(n_1254),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1221),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1204),
.A2(n_1294),
.B(n_1227),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1260),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1222),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1250),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1250),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1244),
.B(n_1228),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1235),
.B(n_1271),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1224),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1293),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1251),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1247),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1234),
.B(n_1244),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1216),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1234),
.B(n_1238),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1219),
.B(n_1214),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1256),
.B(n_1231),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1219),
.B(n_1218),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1265),
.B(n_1238),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1239),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1212),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1269),
.B(n_1225),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1213),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1246),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1213),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1243),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1255),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_SL g1333 ( 
.A(n_1207),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1245),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1294),
.A2(n_1227),
.B(n_1233),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1236),
.A2(n_1255),
.B(n_1237),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1220),
.Y(n_1337)
);

AO21x1_ASAP7_75t_SL g1338 ( 
.A1(n_1257),
.A2(n_1295),
.B(n_1245),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1295),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1257),
.B(n_1209),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1269),
.B(n_1225),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1292),
.A2(n_1253),
.B1(n_1279),
.B2(n_1208),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_1264),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1248),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1303),
.B(n_1262),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1304),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1327),
.Y(n_1347)
);

OAI211xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1322),
.A2(n_1280),
.B(n_1273),
.C(n_1275),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1319),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1297),
.B(n_1336),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_1327),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1310),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1311),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1302),
.B(n_1272),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1297),
.B(n_1272),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1344),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1312),
.B(n_1277),
.Y(n_1357)
);

OAI211xp5_ASAP7_75t_L g1358 ( 
.A1(n_1305),
.A2(n_1342),
.B(n_1287),
.C(n_1283),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1312),
.B(n_1282),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1331),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1324),
.B(n_1281),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1332),
.B(n_1279),
.C(n_1287),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_SL g1363 ( 
.A(n_1338),
.B(n_1292),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1318),
.A2(n_1292),
.B1(n_1205),
.B2(n_1264),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1334),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1321),
.B(n_1268),
.Y(n_1366)
);

BUFx12f_ASAP7_75t_L g1367 ( 
.A(n_1319),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1324),
.B(n_1270),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1324),
.B(n_1215),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1321),
.B(n_1268),
.Y(n_1370)
);

INVx4_ASAP7_75t_L g1371 ( 
.A(n_1304),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1339),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1323),
.B(n_1307),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1304),
.Y(n_1374)
);

INVx5_ASAP7_75t_L g1375 ( 
.A(n_1316),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1323),
.B(n_1285),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1307),
.B(n_1215),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1313),
.B(n_1215),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1306),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1296),
.Y(n_1380)
);

INVxp33_ASAP7_75t_L g1381 ( 
.A(n_1333),
.Y(n_1381)
);

AND2x4_ASAP7_75t_SL g1382 ( 
.A(n_1340),
.B(n_1205),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1332),
.B(n_1290),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_SL g1384 ( 
.A(n_1337),
.B(n_1220),
.C(n_1291),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1347),
.B(n_1341),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1373),
.B(n_1301),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1347),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1380),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1380),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1351),
.B(n_1341),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1371),
.B(n_1308),
.Y(n_1391)
);

NOR2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1371),
.B(n_1319),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1373),
.B(n_1301),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1357),
.B(n_1301),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1375),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1357),
.B(n_1301),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1368),
.B(n_1324),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1352),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1359),
.B(n_1335),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1359),
.B(n_1335),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1378),
.B(n_1335),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1376),
.B(n_1326),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1365),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1356),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1371),
.B(n_1209),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1346),
.B(n_1210),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1376),
.B(n_1326),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1360),
.B(n_1309),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1345),
.A2(n_1320),
.B1(n_1266),
.B2(n_1229),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1404),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1385),
.B(n_1350),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1388),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1394),
.B(n_1366),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1394),
.B(n_1370),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1396),
.B(n_1370),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1386),
.B(n_1383),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1388),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1389),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1399),
.B(n_1369),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1386),
.B(n_1383),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1399),
.B(n_1369),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1385),
.B(n_1354),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1391),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1400),
.B(n_1369),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1400),
.B(n_1355),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1389),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1390),
.B(n_1354),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1393),
.B(n_1355),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1393),
.B(n_1377),
.Y(n_1429)
);

AND2x4_ASAP7_75t_SL g1430 ( 
.A(n_1397),
.B(n_1361),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1428),
.B(n_1390),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1429),
.B(n_1413),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1412),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1412),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1429),
.B(n_1398),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1410),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1423),
.A2(n_1392),
.B(n_1382),
.C(n_1391),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1428),
.B(n_1401),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1417),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1425),
.B(n_1402),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1417),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1414),
.B(n_1403),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1425),
.B(n_1402),
.Y(n_1444)
);

NOR2xp33_ASAP7_75t_L g1445 ( 
.A(n_1411),
.B(n_1349),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1418),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1415),
.B(n_1407),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1415),
.B(n_1408),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1426),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1449),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1431),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1436),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1437),
.A2(n_1423),
.B(n_1381),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_SL g1454 ( 
.A1(n_1437),
.A2(n_1405),
.B(n_1384),
.C(n_1392),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_L g1455 ( 
.A(n_1445),
.B(n_1409),
.C(n_1353),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1435),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1436),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1440),
.B(n_1419),
.Y(n_1458)
);

O2A1O1Ixp5_ASAP7_75t_L g1459 ( 
.A1(n_1443),
.A2(n_1358),
.B(n_1406),
.C(n_1416),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1449),
.Y(n_1460)
);

NAND2x1_ASAP7_75t_L g1461 ( 
.A(n_1440),
.B(n_1387),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1438),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1448),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1431),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1438),
.Y(n_1465)
);

OAI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1433),
.A2(n_1364),
.B1(n_1411),
.B2(n_1205),
.C(n_1317),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1444),
.A2(n_1283),
.B(n_1387),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1444),
.B(n_1419),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1434),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1439),
.Y(n_1470)
);

OAI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1461),
.A2(n_1432),
.B(n_1441),
.Y(n_1471)
);

AOI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1459),
.A2(n_1456),
.B1(n_1463),
.B2(n_1454),
.C(n_1465),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_L g1473 ( 
.A(n_1453),
.B(n_1455),
.C(n_1461),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1469),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1458),
.B(n_1447),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1467),
.A2(n_1363),
.B(n_1395),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1469),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1466),
.A2(n_1422),
.B1(n_1427),
.B2(n_1317),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1462),
.B(n_1447),
.Y(n_1479)
);

AOI21xp33_ASAP7_75t_L g1480 ( 
.A1(n_1470),
.A2(n_1367),
.B(n_1298),
.Y(n_1480)
);

AOI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1462),
.A2(n_1465),
.B1(n_1451),
.B2(n_1464),
.C(n_1470),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1473),
.Y(n_1482)
);

NAND4xp25_ASAP7_75t_L g1483 ( 
.A(n_1472),
.B(n_1217),
.C(n_1348),
.D(n_1210),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1471),
.A2(n_1363),
.B(n_1458),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1481),
.B(n_1468),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1480),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1480),
.B(n_1367),
.Y(n_1487)
);

INVxp67_ASAP7_75t_SL g1488 ( 
.A(n_1474),
.Y(n_1488)
);

O2A1O1Ixp5_ASAP7_75t_L g1489 ( 
.A1(n_1478),
.A2(n_1450),
.B(n_1460),
.C(n_1457),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1476),
.A2(n_1382),
.B(n_1291),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1477),
.A2(n_1450),
.B1(n_1468),
.B2(n_1460),
.C(n_1372),
.Y(n_1491)
);

NOR2x1_ASAP7_75t_L g1492 ( 
.A(n_1475),
.B(n_1242),
.Y(n_1492)
);

OAI221xp5_ASAP7_75t_SL g1493 ( 
.A1(n_1479),
.A2(n_1422),
.B1(n_1427),
.B2(n_1420),
.C(n_1416),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1472),
.A2(n_1430),
.B(n_1452),
.Y(n_1494)
);

NOR2x1p5_ASAP7_75t_SL g1495 ( 
.A(n_1482),
.B(n_1452),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1486),
.A2(n_1242),
.B(n_1457),
.Y(n_1496)
);

OAI211xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1487),
.A2(n_1286),
.B(n_1298),
.C(n_1280),
.Y(n_1497)
);

NOR3xp33_ASAP7_75t_L g1498 ( 
.A(n_1483),
.B(n_1286),
.C(n_1252),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_SL g1499 ( 
.A(n_1492),
.B(n_1298),
.Y(n_1499)
);

NAND4xp25_ASAP7_75t_SL g1500 ( 
.A(n_1484),
.B(n_1298),
.C(n_1274),
.D(n_1288),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1494),
.B(n_1216),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1491),
.B(n_1485),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1490),
.A2(n_1419),
.B1(n_1421),
.B2(n_1424),
.Y(n_1503)
);

NOR2xp67_ASAP7_75t_L g1504 ( 
.A(n_1489),
.B(n_1395),
.Y(n_1504)
);

AOI31xp33_ASAP7_75t_L g1505 ( 
.A1(n_1499),
.A2(n_1230),
.A3(n_1488),
.B(n_1223),
.Y(n_1505)
);

AND3x4_ASAP7_75t_L g1506 ( 
.A(n_1498),
.B(n_1230),
.C(n_1223),
.Y(n_1506)
);

NAND4xp25_ASAP7_75t_L g1507 ( 
.A(n_1502),
.B(n_1493),
.C(n_1252),
.D(n_1211),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1500),
.B(n_1242),
.Y(n_1508)
);

AOI211xp5_ASAP7_75t_L g1509 ( 
.A1(n_1497),
.A2(n_1263),
.B(n_1343),
.C(n_1362),
.Y(n_1509)
);

NOR3xp33_ASAP7_75t_SL g1510 ( 
.A(n_1501),
.B(n_1274),
.C(n_1284),
.Y(n_1510)
);

NAND3xp33_ASAP7_75t_L g1511 ( 
.A(n_1496),
.B(n_1315),
.C(n_1233),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1504),
.Y(n_1512)
);

NOR3xp33_ASAP7_75t_L g1513 ( 
.A(n_1495),
.B(n_1278),
.C(n_1259),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1508),
.B(n_1503),
.Y(n_1514)
);

NAND2x1p5_ASAP7_75t_SL g1515 ( 
.A(n_1506),
.B(n_1300),
.Y(n_1515)
);

NOR2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1512),
.B(n_1306),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1507),
.B(n_1420),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1511),
.B(n_1442),
.Y(n_1518)
);

NOR2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1505),
.B(n_1374),
.Y(n_1519)
);

NAND4xp75_ASAP7_75t_L g1520 ( 
.A(n_1510),
.B(n_1300),
.C(n_1328),
.D(n_1330),
.Y(n_1520)
);

XNOR2xp5_ASAP7_75t_L g1521 ( 
.A(n_1513),
.B(n_1232),
.Y(n_1521)
);

NOR3xp33_ASAP7_75t_L g1522 ( 
.A(n_1509),
.B(n_1263),
.C(n_1259),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1518),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1521),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_SL g1525 ( 
.A(n_1520),
.B(n_1299),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1517),
.B(n_1446),
.Y(n_1526)
);

XOR2xp5_ASAP7_75t_L g1527 ( 
.A(n_1514),
.B(n_1232),
.Y(n_1527)
);

AND2x2_ASAP7_75t_SL g1528 ( 
.A(n_1524),
.B(n_1522),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1523),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1527),
.A2(n_1516),
.B1(n_1519),
.B2(n_1515),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1529),
.Y(n_1531)
);

AO22x2_ASAP7_75t_L g1532 ( 
.A1(n_1531),
.A2(n_1530),
.B1(n_1528),
.B2(n_1526),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1531),
.B(n_1526),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1533),
.A2(n_1525),
.B(n_1516),
.C(n_1532),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_SL g1535 ( 
.A(n_1534),
.B(n_1226),
.Y(n_1535)
);

AO221x2_ASAP7_75t_L g1536 ( 
.A1(n_1535),
.A2(n_1261),
.B1(n_1329),
.B2(n_1325),
.C(n_1314),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1536),
.A2(n_1379),
.B1(n_1374),
.B2(n_1299),
.Y(n_1537)
);


endmodule