module fake_netlist_6_1429_n_2106 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2106);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2106;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1052;
wire n_1033;
wire n_462;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_160),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_75),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_95),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_136),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_30),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_81),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_40),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_36),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_123),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_188),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_51),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_150),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_158),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_24),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_102),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_114),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_42),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_80),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_118),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_169),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_22),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_194),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_39),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_101),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_113),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_181),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_124),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_171),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_157),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_65),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_141),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_15),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_110),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_142),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_49),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_154),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_109),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_116),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_129),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_24),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_164),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_62),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_215),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_53),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_148),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_202),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_60),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_79),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_29),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_107),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_46),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_163),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_108),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_1),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_43),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_134),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_40),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_140),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_63),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_179),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_195),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_9),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_26),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_27),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_61),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_198),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_37),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_153),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_212),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_137),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_204),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_26),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_145),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_182),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_183),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_165),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_59),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_17),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_126),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_192),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_191),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_18),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_55),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_1),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_203),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_111),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_57),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_51),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_120),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_201),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_200),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_151),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_146),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_197),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_175),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_176),
.Y(n_320)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_173),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_76),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_93),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_190),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_49),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_55),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_147),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_33),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_91),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_83),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_106),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_29),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_4),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_135),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_43),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_2),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_3),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_78),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_75),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_25),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_39),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_70),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_44),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_94),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_18),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_143),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_34),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_104),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_189),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_67),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_207),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_174),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_122),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_167),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_28),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_132),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_64),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_178),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_46),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_64),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_155),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_82),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_168),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_10),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_209),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_97),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_21),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_144),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_130),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_21),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_66),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_86),
.Y(n_372)
);

BUFx5_ASAP7_75t_L g373 ( 
.A(n_196),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_32),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_7),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_180),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_205),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_4),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_35),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_159),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_50),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_206),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_92),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_41),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_131),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_25),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_2),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_44),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_177),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_138),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_36),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_33),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_99),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_70),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_119),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_216),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_186),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_68),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_84),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_47),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_28),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_17),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_59),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_16),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_9),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_125),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_185),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_3),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_32),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_10),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_103),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_53),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_90),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_19),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_8),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_37),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_117),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_5),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_199),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_112),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_71),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_50),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_214),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_71),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_208),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_73),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_6),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_54),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_213),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_7),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_23),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_8),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_272),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_217),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_225),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g440 ( 
.A(n_271),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_396),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_217),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_219),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_355),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_336),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_235),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_220),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_222),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_357),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_319),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_246),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_246),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_265),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_227),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_405),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_231),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_305),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_265),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_302),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_239),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_239),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_302),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_233),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_306),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_306),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_243),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_277),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_218),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_431),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_234),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_257),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_260),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_305),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g483 ( 
.A(n_254),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_277),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_243),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_255),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_259),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_262),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_257),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_266),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_323),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_278),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_281),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_283),
.Y(n_494)
);

INVxp33_ASAP7_75t_SL g495 ( 
.A(n_245),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_288),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_296),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_301),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_307),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_329),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_308),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_267),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_311),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_332),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_339),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_341),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_343),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_370),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_379),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_386),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_257),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_257),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_388),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_323),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_391),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_392),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_245),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_394),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_270),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_421),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_403),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_299),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_313),
.Y(n_526)
);

INVxp33_ASAP7_75t_SL g527 ( 
.A(n_426),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_414),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_414),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_426),
.Y(n_530)
);

INVxp33_ASAP7_75t_SL g531 ( 
.A(n_427),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_295),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_295),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_300),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_300),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_315),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_304),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_304),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_257),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_427),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_303),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_235),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_428),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_316),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_303),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_324),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_309),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_344),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_344),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_309),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_334),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_399),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_436),
.B(n_298),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_445),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_435),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_532),
.A2(n_389),
.B(n_322),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_437),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_480),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_474),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_451),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_453),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_SL g564 ( 
.A(n_440),
.B(n_287),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_437),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_438),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_R g568 ( 
.A(n_433),
.B(n_399),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_441),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_442),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_461),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_439),
.A2(n_342),
.B1(n_364),
.B2(n_287),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_459),
.B(n_298),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_442),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_436),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_450),
.A2(n_364),
.B1(n_374),
.B2(n_342),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_532),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_464),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_446),
.B(n_447),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_480),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_533),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_471),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_446),
.B(n_318),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_489),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_443),
.A2(n_430),
.B1(n_374),
.B2(n_456),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_489),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_511),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_511),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_512),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_533),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_512),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_479),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_534),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_539),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_535),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_482),
.B(n_491),
.Y(n_599)
);

OA21x2_ASAP7_75t_L g600 ( 
.A1(n_535),
.A2(n_389),
.B(n_322),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_537),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_537),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_538),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_468),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_538),
.Y(n_605)
);

CKINVDCx6p67_ASAP7_75t_R g606 ( 
.A(n_500),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_547),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_469),
.B(n_321),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_547),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_447),
.B(n_318),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_485),
.B(n_261),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_444),
.B(n_430),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_514),
.B(n_327),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_R g614 ( 
.A(n_481),
.B(n_338),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_550),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_550),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_476),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_476),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_474),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_448),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_448),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_477),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_L g623 ( 
.A(n_488),
.B(n_428),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_477),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_542),
.A2(n_268),
.B1(n_286),
.B2(n_252),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_502),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_460),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_519),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_478),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_449),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_R g631 ( 
.A(n_495),
.B(n_238),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_452),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_523),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_517),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_478),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_458),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_452),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_454),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_454),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_486),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_486),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_455),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_487),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_520),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_455),
.Y(n_645)
);

AO22x2_ASAP7_75t_L g646 ( 
.A1(n_577),
.A2(n_327),
.B1(n_354),
.B2(n_348),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_599),
.B(n_473),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_599),
.B(n_526),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_585),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_584),
.B(n_228),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_574),
.A2(n_530),
.B1(n_520),
.B2(n_348),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_555),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_636),
.Y(n_653)
);

AOI21x1_ASAP7_75t_L g654 ( 
.A1(n_558),
.A2(n_229),
.B(n_223),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_555),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_588),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_R g657 ( 
.A(n_568),
.B(n_527),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_SL g658 ( 
.A1(n_611),
.A2(n_470),
.B(n_467),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_585),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_585),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_555),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_587),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_577),
.B(n_549),
.C(n_545),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_587),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_559),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_588),
.Y(n_666)
);

AOI21x1_ASAP7_75t_L g667 ( 
.A1(n_558),
.A2(n_237),
.B(n_236),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_559),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_588),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_587),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_580),
.B(n_458),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_636),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_567),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_574),
.B(n_536),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_589),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_589),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_567),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_589),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_613),
.B(n_544),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_592),
.Y(n_682)
);

AO21x2_ASAP7_75t_L g683 ( 
.A1(n_613),
.A2(n_274),
.B(n_263),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_636),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_608),
.B(n_546),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_567),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_569),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_604),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_608),
.B(n_551),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_569),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_588),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_569),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_584),
.A2(n_530),
.B1(n_354),
.B2(n_531),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_596),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_588),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_584),
.A2(n_610),
.B1(n_580),
.B2(n_554),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_596),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_575),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_584),
.B(n_465),
.Y(n_699)
);

BUFx6f_ASAP7_75t_SL g700 ( 
.A(n_554),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_596),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_560),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_614),
.B(n_540),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_588),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_560),
.Y(n_705)
);

BUFx4f_ASAP7_75t_L g706 ( 
.A(n_558),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_575),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_604),
.Y(n_708)
);

AO21x2_ASAP7_75t_L g709 ( 
.A1(n_623),
.A2(n_280),
.B(n_276),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_561),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_586),
.A2(n_321),
.B1(n_224),
.B2(n_226),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_575),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_556),
.B(n_261),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_L g714 ( 
.A1(n_586),
.A2(n_398),
.B1(n_402),
.B2(n_326),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_632),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_625),
.A2(n_416),
.B1(n_408),
.B2(n_230),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_562),
.B(n_521),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_631),
.A2(n_543),
.B1(n_240),
.B2(n_241),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_634),
.Y(n_719)
);

INVx4_ASAP7_75t_L g720 ( 
.A(n_565),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_610),
.B(n_465),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_632),
.Y(n_722)
);

INVx5_ASAP7_75t_L g723 ( 
.A(n_560),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_563),
.B(n_483),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_560),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_572),
.B(n_509),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_581),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_632),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_610),
.B(n_249),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_579),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_561),
.A2(n_475),
.B1(n_484),
.B2(n_466),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_580),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_576),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_634),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_565),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_632),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_610),
.B(n_290),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_581),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_581),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_581),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_583),
.B(n_238),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_632),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_632),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_593),
.B(n_473),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_590),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_642),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_554),
.B(n_349),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_580),
.B(n_467),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_590),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_642),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_642),
.Y(n_751)
);

INVx8_ASAP7_75t_L g752 ( 
.A(n_626),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_554),
.B(n_351),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_576),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_590),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_590),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_642),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_597),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_642),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_619),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_597),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_553),
.B(n_353),
.Y(n_762)
);

CKINVDCx11_ASAP7_75t_R g763 ( 
.A(n_557),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_597),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_628),
.B(n_240),
.Y(n_765)
);

BUFx10_ASAP7_75t_L g766 ( 
.A(n_633),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_565),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_553),
.B(n_358),
.Y(n_768)
);

AND2x4_ASAP7_75t_SL g769 ( 
.A(n_606),
.B(n_627),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_642),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_566),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_625),
.A2(n_232),
.B1(n_264),
.B2(n_221),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_619),
.B(n_241),
.Y(n_773)
);

AND2x6_ASAP7_75t_L g774 ( 
.A(n_576),
.B(n_228),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_644),
.B(n_242),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_644),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_606),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_566),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_558),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_617),
.B(n_472),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_565),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_578),
.B(n_472),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_558),
.A2(n_490),
.B1(n_269),
.B2(n_293),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_570),
.B(n_361),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_564),
.A2(n_242),
.B1(n_244),
.B2(n_247),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_570),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_597),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_576),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_576),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_571),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_573),
.B(n_244),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_571),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_606),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_598),
.B(n_362),
.Y(n_794)
);

AND3x2_ASAP7_75t_L g795 ( 
.A(n_617),
.B(n_256),
.C(n_429),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_576),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_601),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_600),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_600),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_578),
.B(n_457),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_573),
.B(n_247),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_565),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_600),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_565),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_648),
.B(n_228),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_760),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_771),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_724),
.B(n_618),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_732),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_675),
.B(n_598),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_732),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_672),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_688),
.B(n_612),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_727),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_681),
.B(n_248),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_706),
.B(n_228),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_696),
.B(n_598),
.Y(n_817)
);

INVxp33_ASAP7_75t_L g818 ( 
.A(n_726),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_647),
.B(n_248),
.Y(n_819)
);

NOR2xp67_ASAP7_75t_L g820 ( 
.A(n_717),
.B(n_618),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_672),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_706),
.B(n_228),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_727),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_SL g824 ( 
.A1(n_798),
.A2(n_598),
.B(n_282),
.C(n_285),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_800),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_800),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_647),
.B(n_250),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_647),
.B(n_250),
.Y(n_828)
);

O2A1O1Ixp5_ASAP7_75t_L g829 ( 
.A1(n_706),
.A2(n_284),
.B(n_294),
.C(n_292),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_714),
.B(n_624),
.C(n_622),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_748),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_748),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_727),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_798),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_688),
.B(n_541),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_792),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_646),
.A2(n_269),
.B1(n_320),
.B2(n_293),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_779),
.B(n_620),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_673),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_779),
.B(n_620),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_646),
.A2(n_269),
.B1(n_320),
.B2(n_293),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_792),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_783),
.B(n_620),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_658),
.B(n_269),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_771),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_647),
.B(n_251),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_L g847 ( 
.A(n_731),
.B(n_716),
.C(n_791),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_708),
.B(n_548),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_685),
.B(n_251),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_673),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_745),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_689),
.B(n_253),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_778),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_801),
.B(n_624),
.C(n_622),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_744),
.B(n_253),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_760),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_745),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_729),
.A2(n_635),
.B(n_640),
.C(n_629),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_745),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_718),
.B(n_629),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_778),
.Y(n_861)
);

BUFx5_ASAP7_75t_L g862 ( 
.A(n_799),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_755),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_653),
.B(n_635),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_658),
.A2(n_709),
.B1(n_737),
.B2(n_684),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_755),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_803),
.B(n_653),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_755),
.B(n_293),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_787),
.B(n_320),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_786),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_786),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_646),
.A2(n_397),
.B1(n_352),
.B2(n_320),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_699),
.B(n_258),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_787),
.B(n_330),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_752),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_794),
.B(n_638),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_721),
.B(n_638),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_708),
.B(n_612),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_709),
.B(n_638),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_709),
.B(n_638),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_790),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_656),
.Y(n_882)
);

OAI21xp33_ASAP7_75t_L g883 ( 
.A1(n_651),
.A2(n_529),
.B(n_528),
.Y(n_883)
);

NOR2x1p5_ASAP7_75t_L g884 ( 
.A(n_777),
.B(n_273),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_790),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_747),
.A2(n_552),
.B1(n_376),
.B2(n_372),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_654),
.A2(n_310),
.B(n_297),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_L g888 ( 
.A(n_711),
.B(n_641),
.C(n_640),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_797),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_787),
.B(n_602),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_702),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_762),
.B(n_602),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_719),
.B(n_641),
.Y(n_893)
);

O2A1O1Ixp5_ASAP7_75t_L g894 ( 
.A1(n_654),
.A2(n_417),
.B(n_317),
.C(n_413),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_702),
.Y(n_895)
);

INVx5_ASAP7_75t_L g896 ( 
.A(n_774),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_768),
.B(n_602),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_705),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_784),
.B(n_602),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_741),
.B(n_258),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_652),
.Y(n_901)
);

OAI22xp33_ASAP7_75t_L g902 ( 
.A1(n_780),
.A2(n_346),
.B1(n_411),
.B2(n_331),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_683),
.B(n_602),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_782),
.A2(n_643),
.B(n_582),
.C(n_591),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_683),
.B(n_695),
.Y(n_905)
);

NAND2xp33_ASAP7_75t_L g906 ( 
.A(n_650),
.B(n_257),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_705),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_753),
.A2(n_395),
.B1(n_366),
.B2(n_368),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_652),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_765),
.B(n_419),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_655),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_655),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_725),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_715),
.B(n_330),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_650),
.B(n_373),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_725),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_L g917 ( 
.A(n_693),
.B(n_279),
.C(n_275),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_738),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_703),
.B(n_419),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_666),
.B(n_601),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_661),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_752),
.B(n_528),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_646),
.A2(n_397),
.B1(n_352),
.B2(n_330),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_763),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_661),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_715),
.B(n_330),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_722),
.B(n_330),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_719),
.B(n_643),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_776),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_666),
.B(n_603),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_670),
.B(n_603),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_L g932 ( 
.A(n_650),
.B(n_373),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_734),
.B(n_529),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_738),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_657),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_722),
.B(n_352),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_739),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_754),
.B(n_314),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_670),
.B(n_603),
.Y(n_939)
);

NOR3xp33_ASAP7_75t_L g940 ( 
.A(n_773),
.B(n_493),
.C(n_492),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_420),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_734),
.B(n_582),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_665),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_796),
.A2(n_616),
.B(n_607),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_L g945 ( 
.A(n_663),
.B(n_493),
.C(n_492),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_728),
.B(n_352),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_728),
.B(n_352),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_710),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_739),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_736),
.B(n_397),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_740),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_700),
.A2(n_780),
.B1(n_713),
.B2(n_785),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_736),
.B(n_397),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_742),
.B(n_373),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_776),
.B(n_710),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_795),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_740),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_665),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_700),
.A2(n_406),
.B1(n_382),
.B2(n_383),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_749),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_780),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_668),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_749),
.B(n_607),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_742),
.B(n_373),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_780),
.B(n_420),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_756),
.B(n_616),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_818),
.B(n_730),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_834),
.B(n_752),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_807),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_807),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_837),
.A2(n_772),
.B1(n_793),
.B2(n_777),
.Y(n_971)
);

AND2x6_ASAP7_75t_SL g972 ( 
.A(n_835),
.B(n_494),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_955),
.B(n_730),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_871),
.Y(n_974)
);

NOR2x2_ASAP7_75t_L g975 ( 
.A(n_922),
.B(n_769),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_871),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_834),
.B(n_756),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_891),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_839),
.B(n_769),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_935),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_808),
.B(n_730),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_875),
.B(n_754),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_924),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_895),
.Y(n_984)
);

O2A1O1Ixp5_ASAP7_75t_L g985 ( 
.A1(n_805),
.A2(n_667),
.B(n_796),
.C(n_746),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_SL g986 ( 
.A1(n_813),
.A2(n_878),
.B1(n_793),
.B2(n_948),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_847),
.A2(n_700),
.B1(n_650),
.B2(n_758),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_892),
.A2(n_691),
.B(n_656),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_875),
.B(n_752),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_839),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_848),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_834),
.B(n_758),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_850),
.B(n_494),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_834),
.B(n_862),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_898),
.Y(n_995)
);

AND3x1_ASAP7_75t_SL g996 ( 
.A(n_884),
.B(n_497),
.C(n_496),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_864),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_907),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_815),
.B(n_761),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_806),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_913),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_889),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_856),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_815),
.B(n_761),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_855),
.B(n_764),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_831),
.A2(n_764),
.B1(n_746),
.B2(n_750),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_834),
.B(n_649),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_834),
.B(n_649),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_929),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_855),
.B(n_788),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_933),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_864),
.B(n_862),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_850),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_862),
.B(n_659),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_814),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_832),
.A2(n_660),
.B1(n_662),
.B2(n_659),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_862),
.B(n_660),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_862),
.B(n_662),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_862),
.B(n_664),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_889),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_823),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_810),
.B(n_664),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_922),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_836),
.B(n_671),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_893),
.B(n_766),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_849),
.B(n_766),
.Y(n_1026)
);

OR2x6_ASAP7_75t_L g1027 ( 
.A(n_922),
.B(n_766),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_842),
.B(n_671),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_867),
.B(n_676),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_825),
.B(n_676),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_805),
.A2(n_677),
.B1(n_679),
.B2(n_680),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_916),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_918),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_820),
.B(n_788),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_826),
.B(n_677),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_934),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_849),
.B(n_656),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_928),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_888),
.A2(n_679),
.B1(n_680),
.B2(n_682),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_956),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_937),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_852),
.B(n_425),
.C(n_423),
.Y(n_1042)
);

AND2x6_ASAP7_75t_SL g1043 ( 
.A(n_852),
.B(n_496),
.Y(n_1043)
);

INVx5_ASAP7_75t_L g1044 ( 
.A(n_882),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_949),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_833),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_882),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_873),
.B(n_788),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_812),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_941),
.B(n_910),
.C(n_900),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_821),
.B(n_497),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_901),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_909),
.Y(n_1053)
);

AND2x6_ASAP7_75t_SL g1054 ( 
.A(n_941),
.B(n_498),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_942),
.B(n_423),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_865),
.A2(n_743),
.B1(n_750),
.B2(n_751),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_900),
.B(n_425),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_851),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_951),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_957),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_960),
.Y(n_1061)
);

OR2x2_ASAP7_75t_SL g1062 ( 
.A(n_917),
.B(n_356),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_896),
.B(n_804),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_838),
.B(n_694),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_882),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_882),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_830),
.A2(n_701),
.B1(n_697),
.B2(n_377),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_840),
.B(n_877),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_961),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_809),
.A2(n_751),
.B1(n_770),
.B2(n_757),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_811),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_845),
.B(n_853),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_861),
.B(n_697),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_870),
.B(n_701),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_844),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_860),
.B(n_498),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_881),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_910),
.B(n_919),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_854),
.B(n_499),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_885),
.B(n_757),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_873),
.A2(n_759),
.B1(n_770),
.B2(n_804),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_844),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_819),
.A2(n_827),
.B1(n_846),
.B2(n_828),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_962),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_962),
.Y(n_1085)
);

AND2x6_ASAP7_75t_SL g1086 ( 
.A(n_819),
.B(n_499),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_896),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_827),
.B(n_656),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_886),
.B(n_952),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_945),
.B(n_501),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_857),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_816),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_859),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_817),
.B(n_759),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_828),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_846),
.B(n_656),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_816),
.B(n_668),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_965),
.B(n_691),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_965),
.B(n_691),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_822),
.B(n_669),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_858),
.A2(n_669),
.B(n_712),
.C(n_707),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_863),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_SL g1103 ( 
.A1(n_837),
.A2(n_347),
.B1(n_289),
.B2(n_291),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_822),
.A2(n_804),
.B1(n_365),
.B2(n_369),
.Y(n_1104)
);

NAND2x1_ASAP7_75t_L g1105 ( 
.A(n_866),
.B(n_720),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_896),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_897),
.A2(n_899),
.B(n_876),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_959),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_911),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_908),
.B(n_691),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_896),
.B(n_691),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_938),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_912),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_879),
.B(n_674),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_902),
.B(n_704),
.Y(n_1115)
);

AO22x1_ASAP7_75t_L g1116 ( 
.A1(n_940),
.A2(n_345),
.B1(n_325),
.B2(n_312),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_905),
.A2(n_380),
.B1(n_385),
.B2(n_704),
.Y(n_1117)
);

AND2x6_ASAP7_75t_L g1118 ( 
.A(n_903),
.B(n_704),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_938),
.Y(n_1119)
);

AND2x4_ASAP7_75t_SL g1120 ( 
.A(n_921),
.B(n_704),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_925),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_880),
.B(n_674),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_883),
.B(n_704),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_894),
.A2(n_667),
.B(n_678),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_954),
.B(n_501),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_943),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_SL g1127 ( 
.A(n_904),
.B(n_333),
.C(n_328),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_954),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_841),
.B(n_503),
.Y(n_1129)
);

AND3x1_ASAP7_75t_L g1130 ( 
.A(n_841),
.B(n_504),
.C(n_503),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_872),
.B(n_733),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_843),
.B(n_678),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_958),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_963),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_966),
.Y(n_1135)
);

BUFx8_ASAP7_75t_L g1136 ( 
.A(n_923),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_964),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_964),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_923),
.B(n_733),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_868),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_890),
.B(n_504),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_920),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_887),
.A2(n_690),
.B1(n_698),
.B2(n_707),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_930),
.B(n_335),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_931),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_939),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_1003),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1025),
.Y(n_1148)
);

INVx6_ASAP7_75t_L g1149 ( 
.A(n_990),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_988),
.A2(n_829),
.B(n_944),
.Y(n_1150)
);

BUFx8_ASAP7_75t_SL g1151 ( 
.A(n_983),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_1009),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1134),
.B(n_868),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1066),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1050),
.A2(n_824),
.B(n_869),
.C(n_874),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_994),
.A2(n_735),
.B(n_720),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_994),
.A2(n_767),
.B(n_720),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1087),
.A2(n_781),
.B(n_733),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1083),
.B(n_363),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1057),
.A2(n_824),
.B(n_950),
.C(n_947),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_997),
.B(n_393),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_997),
.B(n_407),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1026),
.B(n_789),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_980),
.B(n_337),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1135),
.B(n_686),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_990),
.Y(n_1166)
);

AO21x1_ASAP7_75t_L g1167 ( 
.A1(n_1037),
.A2(n_926),
.B(n_914),
.Y(n_1167)
);

NOR2xp67_ASAP7_75t_L g1168 ( 
.A(n_967),
.B(n_914),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_R g1169 ( 
.A(n_1095),
.B(n_906),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1136),
.B(n_789),
.Y(n_1170)
);

OAI21xp33_ASAP7_75t_SL g1171 ( 
.A1(n_1131),
.A2(n_927),
.B(n_926),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1072),
.Y(n_1172)
);

OR2x6_ASAP7_75t_SL g1173 ( 
.A(n_971),
.B(n_340),
.Y(n_1173)
);

BUFx8_ASAP7_75t_L g1174 ( 
.A(n_1040),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1005),
.B(n_686),
.Y(n_1175)
);

O2A1O1Ixp5_ASAP7_75t_L g1176 ( 
.A1(n_1110),
.A2(n_953),
.B(n_950),
.C(n_947),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1011),
.B(n_350),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1072),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1145),
.B(n_687),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_979),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1146),
.B(n_1136),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1038),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_990),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1049),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1012),
.B(n_687),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_991),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1087),
.A2(n_789),
.B(n_915),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1068),
.B(n_690),
.Y(n_1188)
);

NOR3xp33_ASAP7_75t_SL g1189 ( 
.A(n_986),
.B(n_359),
.C(n_360),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1002),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1087),
.A2(n_789),
.B(n_932),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1068),
.B(n_692),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1013),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_973),
.B(n_367),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1020),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1129),
.B(n_692),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1000),
.Y(n_1197)
);

OAI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_1090),
.A2(n_375),
.B(n_378),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_999),
.B(n_1004),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_SL g1200 ( 
.A1(n_1088),
.A2(n_712),
.B(n_698),
.C(n_595),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1087),
.A2(n_1107),
.B(n_1114),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_970),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_979),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1089),
.A2(n_373),
.B1(n_390),
.B2(n_936),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1042),
.A2(n_953),
.B(n_946),
.C(n_515),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1114),
.A2(n_789),
.B(n_802),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1122),
.A2(n_802),
.B(n_946),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1092),
.A2(n_1075),
.B1(n_1082),
.B2(n_1096),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1013),
.B(n_971),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1122),
.A2(n_802),
.B(n_723),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1103),
.A2(n_373),
.B1(n_390),
.B2(n_595),
.Y(n_1211)
);

O2A1O1Ixp5_ASAP7_75t_L g1212 ( 
.A1(n_1098),
.A2(n_591),
.B(n_594),
.C(n_609),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1141),
.B(n_616),
.Y(n_1213)
);

NOR3xp33_ASAP7_75t_SL g1214 ( 
.A(n_981),
.B(n_381),
.C(n_384),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_989),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_1027),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1076),
.B(n_802),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1044),
.A2(n_1065),
.B(n_1047),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1044),
.A2(n_723),
.B(n_594),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1076),
.B(n_605),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1112),
.B(n_605),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_SL g1222 ( 
.A(n_1119),
.B(n_387),
.Y(n_1222)
);

O2A1O1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1055),
.A2(n_510),
.B(n_513),
.C(n_516),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_993),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1086),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1137),
.A2(n_404),
.B1(n_418),
.B2(n_415),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_SL g1227 ( 
.A1(n_1108),
.A2(n_401),
.B1(n_409),
.B2(n_410),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1069),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1141),
.B(n_615),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_993),
.Y(n_1230)
);

OAI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1023),
.A2(n_412),
.B1(n_510),
.B2(n_513),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1079),
.B(n_505),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1071),
.B(n_505),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_996),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1144),
.A2(n_774),
.B1(n_621),
.B2(n_645),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1142),
.B(n_621),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1010),
.A2(n_723),
.B1(n_621),
.B2(n_645),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_987),
.A2(n_723),
.B1(n_630),
.B2(n_645),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_SL g1239 ( 
.A1(n_1099),
.A2(n_516),
.B(n_506),
.C(n_507),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_SL g1240 ( 
.A1(n_1139),
.A2(n_515),
.B(n_506),
.C(n_507),
.Y(n_1240)
);

NAND2xp33_ASAP7_75t_R g1241 ( 
.A(n_1127),
.B(n_77),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1051),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1079),
.B(n_1125),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1044),
.B(n_723),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1047),
.A2(n_639),
.B(n_637),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1047),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1047),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1052),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1030),
.B(n_630),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1043),
.B(n_5),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_R g1251 ( 
.A(n_1054),
.B(n_85),
.Y(n_1251)
);

NOR3xp33_ASAP7_75t_SL g1252 ( 
.A(n_978),
.B(n_995),
.C(n_984),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1027),
.B(n_508),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_998),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1062),
.B(n_6),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1053),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1065),
.Y(n_1257)
);

BUFx4f_ASAP7_75t_L g1258 ( 
.A(n_1027),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1001),
.B(n_11),
.Y(n_1259)
);

AOI221xp5_ASAP7_75t_L g1260 ( 
.A1(n_1116),
.A2(n_522),
.B1(n_525),
.B2(n_524),
.C(n_508),
.Y(n_1260)
);

NOR3xp33_ASAP7_75t_SL g1261 ( 
.A(n_1032),
.B(n_518),
.C(n_522),
.Y(n_1261)
);

OAI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1033),
.A2(n_524),
.B(n_525),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1030),
.B(n_630),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1035),
.B(n_637),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1035),
.B(n_774),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_974),
.Y(n_1266)
);

AOI221xp5_ASAP7_75t_L g1267 ( 
.A1(n_1130),
.A2(n_518),
.B1(n_463),
.B2(n_462),
.C(n_457),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_982),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1022),
.B(n_1029),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1123),
.A2(n_463),
.B1(n_462),
.B2(n_390),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1007),
.A2(n_774),
.B(n_133),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1036),
.B(n_390),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1007),
.A2(n_774),
.B(n_139),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1041),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1274)
);

OR2x6_ASAP7_75t_L g1275 ( 
.A(n_982),
.B(n_210),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1008),
.A2(n_1017),
.B(n_1014),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1045),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1085),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1022),
.B(n_390),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1059),
.B(n_12),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1060),
.A2(n_390),
.B1(n_14),
.B2(n_15),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1061),
.B(n_13),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1077),
.B(n_193),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1084),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1106),
.B(n_1138),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1029),
.B(n_187),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_SL g1287 ( 
.A1(n_1117),
.A2(n_172),
.B(n_170),
.C(n_162),
.Y(n_1287)
);

OR2x6_ASAP7_75t_SL g1288 ( 
.A(n_975),
.B(n_14),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1008),
.A2(n_161),
.B1(n_156),
.B2(n_149),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_969),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_976),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1128),
.A2(n_16),
.B(n_19),
.C(n_20),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1113),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1018),
.A2(n_128),
.B(n_121),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1066),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1015),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1015),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1019),
.A2(n_105),
.B(n_100),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1201),
.A2(n_968),
.B(n_1048),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1182),
.Y(n_1300)
);

O2A1O1Ixp5_ASAP7_75t_L g1301 ( 
.A1(n_1167),
.A2(n_1115),
.B(n_985),
.C(n_1094),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1171),
.A2(n_1094),
.B(n_1097),
.Y(n_1302)
);

AOI221x1_ASAP7_75t_L g1303 ( 
.A1(n_1231),
.A2(n_1208),
.B1(n_1292),
.B2(n_1270),
.C(n_1255),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1183),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1172),
.B(n_1024),
.Y(n_1305)
);

NOR3xp33_ASAP7_75t_L g1306 ( 
.A(n_1194),
.B(n_1034),
.C(n_1024),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1199),
.B(n_1028),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1237),
.A2(n_1100),
.A3(n_1097),
.B(n_992),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1148),
.B(n_1138),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1279),
.A2(n_1100),
.A3(n_992),
.B(n_977),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1279),
.A2(n_1206),
.A3(n_1207),
.B(n_1286),
.Y(n_1311)
);

NAND2xp33_ASAP7_75t_R g1312 ( 
.A(n_1214),
.B(n_1021),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1243),
.B(n_1133),
.Y(n_1313)
);

INVx4_ASAP7_75t_L g1314 ( 
.A(n_1246),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1150),
.A2(n_1157),
.B(n_1156),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1232),
.B(n_1109),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1249),
.A2(n_1073),
.B(n_1074),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1210),
.A2(n_1124),
.B(n_1185),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1228),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1242),
.B(n_1233),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1184),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1151),
.Y(n_1322)
);

AO21x1_ASAP7_75t_L g1323 ( 
.A1(n_1209),
.A2(n_1028),
.B(n_1056),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1181),
.B(n_1173),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1202),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_L g1326 ( 
.A(n_1147),
.B(n_1091),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1246),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1176),
.A2(n_1080),
.B(n_1101),
.Y(n_1328)
);

OAI22x1_ASAP7_75t_L g1329 ( 
.A1(n_1181),
.A2(n_972),
.B1(n_1140),
.B2(n_1102),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1230),
.B(n_1021),
.Y(n_1330)
);

NAND4xp25_ASAP7_75t_SL g1331 ( 
.A(n_1274),
.B(n_1104),
.C(n_1067),
.D(n_1039),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1252),
.A2(n_1093),
.B(n_1006),
.C(n_1081),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1158),
.A2(n_1191),
.B(n_1187),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1266),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1233),
.B(n_1126),
.Y(n_1335)
);

AOI21xp33_ASAP7_75t_L g1336 ( 
.A1(n_1159),
.A2(n_1073),
.B(n_1074),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1188),
.A2(n_1132),
.B(n_977),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1192),
.A2(n_1179),
.B(n_1245),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1288),
.Y(n_1339)
);

NOR2x1_ASAP7_75t_SL g1340 ( 
.A(n_1257),
.B(n_1064),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1238),
.A2(n_1121),
.A3(n_1118),
.B(n_1031),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1249),
.A2(n_1143),
.B(n_1070),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_L g1343 ( 
.A1(n_1272),
.A2(n_1105),
.B(n_1111),
.C(n_1046),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1179),
.A2(n_1046),
.B(n_1058),
.Y(n_1344)
);

NOR4xp25_ASAP7_75t_L g1345 ( 
.A(n_1281),
.B(n_1016),
.C(n_1058),
.D(n_23),
.Y(n_1345)
);

OAI21xp33_ASAP7_75t_L g1346 ( 
.A1(n_1177),
.A2(n_1120),
.B(n_1063),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1178),
.B(n_1118),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1183),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1215),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1175),
.B(n_1118),
.Y(n_1350)
);

NOR2x1_ASAP7_75t_L g1351 ( 
.A(n_1166),
.B(n_1257),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1284),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_SL g1353 ( 
.A(n_1164),
.B(n_1118),
.Y(n_1353)
);

AO21x2_ASAP7_75t_L g1354 ( 
.A1(n_1200),
.A2(n_98),
.B(n_96),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1155),
.A2(n_89),
.B(n_88),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1254),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1197),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1196),
.A2(n_87),
.B(n_27),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1224),
.B(n_22),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1160),
.A2(n_30),
.B(n_31),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1277),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1291),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1196),
.A2(n_31),
.B(n_34),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1229),
.B(n_35),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1263),
.A2(n_38),
.B(n_42),
.Y(n_1365)
);

OA21x2_ASAP7_75t_L g1366 ( 
.A1(n_1263),
.A2(n_38),
.B(n_45),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1264),
.B(n_45),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1264),
.A2(n_47),
.B(n_48),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1190),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1170),
.A2(n_48),
.B1(n_52),
.B2(n_54),
.Y(n_1370)
);

NOR2x1_ASAP7_75t_L g1371 ( 
.A(n_1166),
.B(n_52),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1153),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1153),
.A2(n_56),
.B(n_58),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1229),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_1374)
);

BUFx10_ASAP7_75t_L g1375 ( 
.A(n_1253),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1186),
.B(n_65),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1183),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1285),
.A2(n_66),
.B(n_67),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1165),
.B(n_68),
.Y(n_1379)
);

AO32x2_ASAP7_75t_L g1380 ( 
.A1(n_1289),
.A2(n_1227),
.A3(n_1226),
.B1(n_1261),
.B2(n_1240),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1195),
.Y(n_1381)
);

AO22x1_ASAP7_75t_L g1382 ( 
.A1(n_1225),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1265),
.A2(n_1218),
.B(n_1236),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1265),
.A2(n_74),
.B(n_1212),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1250),
.A2(n_1198),
.B(n_1259),
.Y(n_1385)
);

AO31x2_ASAP7_75t_L g1386 ( 
.A1(n_1271),
.A2(n_1273),
.A3(n_1213),
.B(n_1298),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1219),
.A2(n_1213),
.B(n_1294),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1152),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1248),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_SL g1390 ( 
.A(n_1258),
.B(n_1216),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1149),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1221),
.B(n_1220),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1168),
.A2(n_1161),
.B(n_1162),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1235),
.A2(n_1204),
.B(n_1205),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1193),
.Y(n_1395)
);

AOI22x1_ASAP7_75t_L g1396 ( 
.A1(n_1256),
.A2(n_1290),
.B1(n_1278),
.B2(n_1293),
.Y(n_1396)
);

O2A1O1Ixp5_ASAP7_75t_L g1397 ( 
.A1(n_1283),
.A2(n_1217),
.B(n_1287),
.C(n_1258),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1211),
.B(n_1280),
.C(n_1282),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1262),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1296),
.B(n_1297),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1246),
.A2(n_1247),
.B(n_1244),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1203),
.B(n_1234),
.Y(n_1402)
);

AND2x6_ASAP7_75t_L g1403 ( 
.A(n_1154),
.B(n_1247),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1247),
.Y(n_1404)
);

NOR4xp25_ASAP7_75t_L g1405 ( 
.A(n_1239),
.B(n_1223),
.C(n_1260),
.D(n_1267),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1180),
.B(n_1189),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1268),
.A2(n_1297),
.B(n_1296),
.C(n_1222),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1296),
.B(n_1297),
.Y(n_1408)
);

AOI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1275),
.A2(n_1169),
.B(n_1241),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1295),
.B(n_1275),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1295),
.B(n_1275),
.Y(n_1411)
);

INVx6_ASAP7_75t_SL g1412 ( 
.A(n_1174),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1295),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1251),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_1174),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1243),
.B(n_1011),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1150),
.A2(n_1201),
.B(n_1206),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1172),
.B(n_1178),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1257),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1202),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1199),
.A2(n_1050),
.B(n_1078),
.C(n_1026),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1167),
.A2(n_1201),
.A3(n_1270),
.B(n_1237),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1202),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1186),
.Y(n_1424)
);

AOI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1163),
.A2(n_1201),
.B(n_1279),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1167),
.A2(n_1201),
.A3(n_1270),
.B(n_1237),
.Y(n_1426)
);

AO31x2_ASAP7_75t_L g1427 ( 
.A1(n_1167),
.A2(n_1201),
.A3(n_1270),
.B(n_1237),
.Y(n_1427)
);

NAND3x1_ASAP7_75t_L g1428 ( 
.A(n_1250),
.B(n_847),
.C(n_573),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_SL g1429 ( 
.A1(n_1269),
.A2(n_994),
.B(n_875),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_L g1430 ( 
.A(n_1255),
.B(n_1026),
.C(n_1078),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1171),
.A2(n_1050),
.B(n_1276),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1181),
.B(n_818),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1171),
.A2(n_1050),
.B(n_1276),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1199),
.A2(n_1050),
.B(n_1078),
.C(n_1026),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1202),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1243),
.B(n_1011),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1202),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1183),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1199),
.B(n_1172),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1167),
.A2(n_1201),
.B(n_1176),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1151),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1171),
.A2(n_1050),
.B(n_1276),
.Y(n_1442)
);

AOI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1163),
.A2(n_1201),
.B(n_1279),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_SL g1444 ( 
.A(n_1148),
.B(n_1025),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1172),
.B(n_1178),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1183),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1201),
.A2(n_968),
.B(n_1269),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1202),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1150),
.A2(n_1201),
.B(n_1206),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1181),
.B(n_818),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1430),
.B(n_1385),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1325),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1357),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1299),
.A2(n_1447),
.B(n_1433),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1430),
.A2(n_1439),
.B1(n_1398),
.B2(n_1307),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1456)
);

OR2x6_ASAP7_75t_SL g1457 ( 
.A(n_1349),
.B(n_1414),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1421),
.A2(n_1434),
.B(n_1306),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1334),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1416),
.B(n_1436),
.Y(n_1460)
);

AO32x2_ASAP7_75t_L g1461 ( 
.A1(n_1372),
.A2(n_1374),
.A3(n_1370),
.B1(n_1360),
.B2(n_1345),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1319),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1352),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1449),
.A2(n_1383),
.B(n_1344),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1403),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1313),
.B(n_1316),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1387),
.A2(n_1328),
.B(n_1425),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1360),
.A2(n_1355),
.B(n_1385),
.C(n_1433),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1318),
.A2(n_1338),
.B(n_1443),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1418),
.A2(n_1445),
.B1(n_1305),
.B2(n_1432),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1420),
.Y(n_1471)
);

OAI221xp5_ASAP7_75t_L g1472 ( 
.A1(n_1345),
.A2(n_1355),
.B1(n_1450),
.B2(n_1324),
.C(n_1444),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1423),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1431),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1424),
.B(n_1357),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1320),
.B(n_1300),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1435),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1437),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1428),
.A2(n_1392),
.B1(n_1326),
.B2(n_1361),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1302),
.A2(n_1301),
.B(n_1337),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1364),
.B(n_1335),
.Y(n_1481)
);

INVx5_ASAP7_75t_L g1482 ( 
.A(n_1403),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1372),
.A2(n_1374),
.B1(n_1370),
.B2(n_1331),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1302),
.A2(n_1317),
.B(n_1442),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1356),
.B(n_1388),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1448),
.Y(n_1487)
);

A2O1A1Ixp33_ASAP7_75t_SL g1488 ( 
.A1(n_1442),
.A2(n_1384),
.B(n_1429),
.C(n_1394),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1396),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1440),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1402),
.A2(n_1329),
.B1(n_1376),
.B2(n_1441),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1390),
.A2(n_1366),
.B1(n_1373),
.B2(n_1363),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1336),
.A2(n_1303),
.B(n_1397),
.Y(n_1493)
);

INVx6_ASAP7_75t_L g1494 ( 
.A(n_1375),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1336),
.A2(n_1332),
.B(n_1405),
.Y(n_1495)
);

INVx8_ASAP7_75t_L g1496 ( 
.A(n_1403),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1440),
.A2(n_1350),
.B(n_1343),
.Y(n_1497)
);

OAI222xp33_ASAP7_75t_L g1498 ( 
.A1(n_1378),
.A2(n_1371),
.B1(n_1353),
.B2(n_1379),
.C1(n_1367),
.C2(n_1399),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1350),
.A2(n_1409),
.B(n_1393),
.Y(n_1499)
);

OA21x2_ASAP7_75t_L g1500 ( 
.A1(n_1323),
.A2(n_1394),
.B(n_1367),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1340),
.A2(n_1346),
.B(n_1347),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1347),
.A2(n_1358),
.B(n_1342),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1342),
.A2(n_1401),
.B(n_1379),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1405),
.A2(n_1330),
.B(n_1309),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1362),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1321),
.B(n_1369),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1381),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1389),
.Y(n_1508)
);

NAND2xp33_ASAP7_75t_SL g1509 ( 
.A(n_1406),
.B(n_1312),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1366),
.A2(n_1419),
.B(n_1351),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1348),
.Y(n_1511)
);

BUFx2_ASAP7_75t_SL g1512 ( 
.A(n_1322),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1412),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1390),
.A2(n_1359),
.B1(n_1382),
.B2(n_1391),
.Y(n_1514)
);

BUFx12f_ASAP7_75t_L g1515 ( 
.A(n_1415),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1407),
.A2(n_1391),
.B1(n_1400),
.B2(n_1408),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1419),
.A2(n_1408),
.B(n_1413),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1311),
.A2(n_1422),
.B(n_1426),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1311),
.A2(n_1386),
.B(n_1427),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1310),
.Y(n_1520)
);

OAI222xp33_ASAP7_75t_L g1521 ( 
.A1(n_1380),
.A2(n_1404),
.B1(n_1327),
.B2(n_1314),
.C1(n_1339),
.C2(n_1412),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1354),
.A2(n_1386),
.B(n_1310),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1310),
.Y(n_1523)
);

AO31x2_ASAP7_75t_L g1524 ( 
.A1(n_1422),
.A2(n_1426),
.A3(n_1308),
.B(n_1354),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1308),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1341),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1341),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1327),
.A2(n_1404),
.B(n_1380),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1304),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1377),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1415),
.A2(n_1395),
.B1(n_1438),
.B2(n_1446),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1438),
.A2(n_1433),
.B(n_1431),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1415),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1438),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1441),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1403),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1409),
.B(n_1275),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1325),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1325),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1409),
.B(n_1275),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1325),
.Y(n_1541)
);

AOI21xp33_ASAP7_75t_L g1542 ( 
.A1(n_1398),
.A2(n_1026),
.B(n_1078),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1441),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1544)
);

NOR2xp67_ASAP7_75t_L g1545 ( 
.A(n_1424),
.B(n_980),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1325),
.Y(n_1546)
);

AOI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1409),
.A2(n_1317),
.B(n_1201),
.Y(n_1547)
);

OAI22x1_ASAP7_75t_L g1548 ( 
.A1(n_1430),
.A2(n_1083),
.B1(n_1026),
.B2(n_1398),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1431),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1300),
.Y(n_1550)
);

CKINVDCx14_ASAP7_75t_R g1551 ( 
.A(n_1441),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1431),
.A2(n_1442),
.B(n_1433),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1398),
.A2(n_1050),
.B1(n_847),
.B2(n_1078),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_SL g1555 ( 
.A(n_1441),
.B(n_1151),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1325),
.Y(n_1556)
);

AOI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1409),
.A2(n_1317),
.B(n_1201),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1398),
.B(n_1026),
.C(n_1078),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1319),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1409),
.B(n_1275),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1325),
.Y(n_1563)
);

BUFx12f_ASAP7_75t_L g1564 ( 
.A(n_1415),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1428),
.A2(n_1050),
.B1(n_1026),
.B2(n_627),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1325),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1385),
.A2(n_1050),
.B(n_1078),
.C(n_1421),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1431),
.A2(n_1442),
.B(n_1433),
.Y(n_1568)
);

NAND3xp33_ASAP7_75t_L g1569 ( 
.A(n_1398),
.B(n_1026),
.C(n_1078),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1319),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1300),
.B(n_1364),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1325),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1418),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1439),
.B(n_1418),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1325),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1325),
.Y(n_1577)
);

OR3x4_ASAP7_75t_SL g1578 ( 
.A(n_1428),
.B(n_456),
.C(n_443),
.Y(n_1578)
);

AOI22x1_ASAP7_75t_L g1579 ( 
.A1(n_1360),
.A2(n_1329),
.B1(n_1355),
.B2(n_1431),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1398),
.A2(n_1050),
.B(n_1078),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1431),
.A2(n_1442),
.B(n_1433),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1319),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1300),
.B(n_1364),
.Y(n_1583)
);

NOR2xp67_ASAP7_75t_L g1584 ( 
.A(n_1424),
.B(n_980),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1325),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1398),
.A2(n_1050),
.B1(n_847),
.B2(n_1078),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1300),
.B(n_1364),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1360),
.A2(n_1136),
.B1(n_444),
.B2(n_460),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1325),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1431),
.A2(n_1442),
.B(n_1433),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1439),
.B(n_1418),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1410),
.B(n_1411),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1325),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1598)
);

BUFx8_ASAP7_75t_L g1599 ( 
.A(n_1415),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1325),
.Y(n_1600)
);

BUFx12f_ASAP7_75t_L g1601 ( 
.A(n_1415),
.Y(n_1601)
);

NAND2x1p5_ASAP7_75t_L g1602 ( 
.A(n_1309),
.B(n_1257),
.Y(n_1602)
);

AOI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1409),
.A2(n_1317),
.B(n_1201),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1325),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1325),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1385),
.A2(n_1050),
.B(n_1078),
.C(n_1421),
.Y(n_1606)
);

OA21x2_ASAP7_75t_L g1607 ( 
.A1(n_1431),
.A2(n_1442),
.B(n_1433),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1416),
.B(n_1436),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1333),
.A2(n_1315),
.B(n_1417),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1325),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1532),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1466),
.B(n_1460),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1470),
.B(n_1575),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1594),
.B(n_1574),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1522),
.A2(n_1493),
.B(n_1484),
.Y(n_1615)
);

O2A1O1Ixp5_ASAP7_75t_L g1616 ( 
.A1(n_1468),
.A2(n_1458),
.B(n_1495),
.C(n_1488),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1574),
.B(n_1455),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1481),
.B(n_1553),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1481),
.B(n_1553),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1608),
.B(n_1451),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1590),
.A2(n_1472),
.B1(n_1565),
.B2(n_1483),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1488),
.A2(n_1468),
.B(n_1454),
.Y(n_1622)
);

O2A1O1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1542),
.A2(n_1606),
.B(n_1567),
.C(n_1580),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1590),
.A2(n_1483),
.B1(n_1588),
.B2(n_1451),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1491),
.A2(n_1588),
.B1(n_1533),
.B2(n_1578),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1459),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1558),
.A2(n_1569),
.B1(n_1579),
.B2(n_1479),
.Y(n_1627)
);

AND2x6_ASAP7_75t_L g1628 ( 
.A(n_1465),
.B(n_1526),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1459),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1572),
.B(n_1583),
.Y(n_1630)
);

CKINVDCx11_ASAP7_75t_R g1631 ( 
.A(n_1515),
.Y(n_1631)
);

O2A1O1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1498),
.A2(n_1514),
.B(n_1521),
.C(n_1504),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1463),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1548),
.A2(n_1536),
.B(n_1537),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1471),
.Y(n_1635)
);

OA21x2_ASAP7_75t_L g1636 ( 
.A1(n_1480),
.A2(n_1490),
.B(n_1519),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1471),
.Y(n_1637)
);

NOR2xp67_ASAP7_75t_L g1638 ( 
.A(n_1545),
.B(n_1584),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1582),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1599),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1478),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1478),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1514),
.A2(n_1498),
.B1(n_1474),
.B2(n_1549),
.C(n_1521),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1462),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1544),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1537),
.A2(n_1562),
.B(n_1540),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1596),
.B(n_1476),
.Y(n_1647)
);

O2A1O1Ixp5_ASAP7_75t_L g1648 ( 
.A1(n_1547),
.A2(n_1603),
.B(n_1557),
.C(n_1528),
.Y(n_1648)
);

AOI21x1_ASAP7_75t_SL g1649 ( 
.A1(n_1461),
.A2(n_1596),
.B(n_1578),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1589),
.A2(n_1453),
.B1(n_1550),
.B2(n_1531),
.Y(n_1650)
);

O2A1O1Ixp5_ASAP7_75t_L g1651 ( 
.A1(n_1501),
.A2(n_1525),
.B(n_1509),
.C(n_1520),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1537),
.B(n_1540),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1506),
.B(n_1485),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1487),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1540),
.A2(n_1562),
.B(n_1552),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1485),
.B(n_1507),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1562),
.A2(n_1552),
.B(n_1568),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1538),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1568),
.A2(n_1593),
.B(n_1581),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1568),
.A2(n_1593),
.B(n_1581),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1507),
.B(n_1475),
.Y(n_1661)
);

OA21x2_ASAP7_75t_L g1662 ( 
.A1(n_1467),
.A2(n_1469),
.B(n_1502),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1551),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1546),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1492),
.A2(n_1550),
.B1(n_1607),
.B2(n_1500),
.C(n_1516),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_SL g1666 ( 
.A(n_1482),
.B(n_1520),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1482),
.B(n_1465),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1502),
.A2(n_1497),
.B(n_1503),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1563),
.B(n_1586),
.Y(n_1669)
);

OA21x2_ASAP7_75t_L g1670 ( 
.A1(n_1497),
.A2(n_1503),
.B(n_1464),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1482),
.B(n_1586),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1532),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1505),
.B(n_1508),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1505),
.B(n_1452),
.Y(n_1674)
);

BUFx10_ASAP7_75t_L g1675 ( 
.A(n_1513),
.Y(n_1675)
);

NOR2x1_ASAP7_75t_SL g1676 ( 
.A(n_1482),
.B(n_1523),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1473),
.B(n_1610),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1477),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1539),
.B(n_1541),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1556),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1531),
.A2(n_1457),
.B1(n_1494),
.B2(n_1570),
.Y(n_1681)
);

OA21x2_ASAP7_75t_L g1682 ( 
.A1(n_1554),
.A2(n_1587),
.B(n_1585),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1566),
.B(n_1573),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1576),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1577),
.B(n_1591),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1597),
.A2(n_1604),
.B(n_1605),
.C(n_1600),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1607),
.A2(n_1532),
.B(n_1602),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1517),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1511),
.B(n_1534),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1529),
.B(n_1530),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1499),
.B(n_1527),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1494),
.A2(n_1559),
.B1(n_1602),
.B2(n_1533),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1512),
.B(n_1551),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1496),
.A2(n_1513),
.B1(n_1564),
.B2(n_1515),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1510),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1564),
.A2(n_1601),
.B1(n_1543),
.B2(n_1535),
.Y(n_1696)
);

OAI31xp33_ASAP7_75t_L g1697 ( 
.A1(n_1555),
.A2(n_1489),
.A3(n_1599),
.B(n_1601),
.Y(n_1697)
);

O2A1O1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1489),
.A2(n_1518),
.B(n_1524),
.C(n_1599),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1535),
.B(n_1543),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1560),
.A2(n_1571),
.B(n_1561),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1592),
.A2(n_1595),
.B1(n_1598),
.B2(n_1609),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1572),
.B(n_1583),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1532),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1468),
.A2(n_1050),
.B(n_1078),
.C(n_1385),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1590),
.A2(n_1173),
.B1(n_1472),
.B2(n_1026),
.Y(n_1705)
);

NOR2x1_ASAP7_75t_SL g1706 ( 
.A(n_1537),
.B(n_1540),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1468),
.A2(n_1026),
.B(n_875),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1468),
.A2(n_1050),
.B(n_1078),
.C(n_1385),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1466),
.B(n_1460),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1522),
.A2(n_1493),
.B(n_1484),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1466),
.B(n_1460),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1453),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1572),
.B(n_1583),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1459),
.Y(n_1714)
);

OA21x2_ASAP7_75t_L g1715 ( 
.A1(n_1522),
.A2(n_1493),
.B(n_1484),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1590),
.A2(n_1173),
.B1(n_1472),
.B2(n_1026),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_SL g1717 ( 
.A1(n_1458),
.A2(n_1026),
.B(n_1360),
.C(n_1493),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1470),
.B(n_1575),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1456),
.B(n_1486),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1590),
.A2(n_1173),
.B1(n_1472),
.B2(n_1026),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1453),
.Y(n_1721)
);

AOI21xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1468),
.A2(n_1026),
.B(n_875),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1590),
.A2(n_1173),
.B1(n_1472),
.B2(n_1026),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1532),
.Y(n_1724)
);

CKINVDCx11_ASAP7_75t_R g1725 ( 
.A(n_1515),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1582),
.Y(n_1726)
);

CKINVDCx16_ASAP7_75t_R g1727 ( 
.A(n_1555),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1535),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1470),
.B(n_1575),
.Y(n_1729)
);

O2A1O1Ixp33_ASAP7_75t_L g1730 ( 
.A1(n_1468),
.A2(n_1050),
.B(n_1078),
.C(n_1385),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1551),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1466),
.B(n_1460),
.Y(n_1732)
);

AND2x6_ASAP7_75t_L g1733 ( 
.A(n_1465),
.B(n_1526),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1459),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1572),
.B(n_1583),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1646),
.B(n_1655),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1626),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1611),
.B(n_1672),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1611),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1652),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1621),
.A2(n_1723),
.B1(n_1720),
.B2(n_1716),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1672),
.B(n_1703),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1724),
.B(n_1615),
.Y(n_1743)
);

AOI21x1_ASAP7_75t_L g1744 ( 
.A1(n_1622),
.A2(n_1627),
.B(n_1701),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1652),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1691),
.Y(n_1746)
);

NOR2xp67_ASAP7_75t_L g1747 ( 
.A(n_1688),
.B(n_1665),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1620),
.B(n_1669),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1633),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1624),
.A2(n_1705),
.B1(n_1616),
.B2(n_1623),
.C(n_1704),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1668),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1678),
.B(n_1680),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1617),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1656),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1695),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1642),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1658),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1664),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1613),
.B(n_1718),
.Y(n_1759)
);

INVx5_ASAP7_75t_L g1760 ( 
.A(n_1628),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1683),
.Y(n_1761)
);

NOR2x1_ASAP7_75t_R g1762 ( 
.A(n_1631),
.B(n_1725),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1685),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1647),
.B(n_1673),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1625),
.A2(n_1619),
.B1(n_1618),
.B2(n_1643),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1714),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1659),
.B(n_1660),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1686),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1684),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1706),
.B(n_1719),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1684),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1636),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1636),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1670),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1670),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1677),
.B(n_1679),
.Y(n_1776)
);

OAI21xp33_ASAP7_75t_L g1777 ( 
.A1(n_1704),
.A2(n_1708),
.B(n_1730),
.Y(n_1777)
);

AO21x2_ASAP7_75t_L g1778 ( 
.A1(n_1717),
.A2(n_1657),
.B(n_1698),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1661),
.B(n_1719),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1729),
.B(n_1614),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1682),
.Y(n_1781)
);

OA21x2_ASAP7_75t_L g1782 ( 
.A1(n_1616),
.A2(n_1648),
.B(n_1651),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1686),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1629),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1645),
.B(n_1635),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1637),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1641),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1671),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1654),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1630),
.B(n_1702),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1662),
.Y(n_1791)
);

OR2x6_ASAP7_75t_L g1792 ( 
.A(n_1687),
.B(n_1634),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1665),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1734),
.B(n_1710),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1674),
.Y(n_1795)
);

OA21x2_ASAP7_75t_L g1796 ( 
.A1(n_1648),
.A2(n_1651),
.B(n_1643),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1710),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1698),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1715),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1713),
.B(n_1735),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1628),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1733),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1666),
.Y(n_1803)
);

OR2x6_ASAP7_75t_L g1804 ( 
.A(n_1707),
.B(n_1722),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1676),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1781),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1794),
.B(n_1743),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1739),
.Y(n_1808)
);

INVx4_ASAP7_75t_L g1809 ( 
.A(n_1760),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1770),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1753),
.B(n_1623),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1791),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1743),
.B(n_1700),
.Y(n_1813)
);

A2O1A1Ixp33_ASAP7_75t_L g1814 ( 
.A1(n_1750),
.A2(n_1632),
.B(n_1730),
.C(n_1708),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1769),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1738),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1753),
.B(n_1653),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1776),
.B(n_1612),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1741),
.A2(n_1765),
.B1(n_1793),
.B2(n_1804),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1750),
.A2(n_1632),
.B(n_1681),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1776),
.B(n_1711),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1771),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1771),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1748),
.B(n_1764),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1760),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1746),
.B(n_1721),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1748),
.B(n_1732),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1746),
.B(n_1712),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1764),
.B(n_1709),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1765),
.A2(n_1697),
.B(n_1696),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1760),
.Y(n_1831)
);

NOR2x1p5_ASAP7_75t_L g1832 ( 
.A(n_1759),
.B(n_1640),
.Y(n_1832)
);

BUFx2_ASAP7_75t_SL g1833 ( 
.A(n_1760),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1770),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1780),
.B(n_1650),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1737),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1793),
.A2(n_1649),
.B1(n_1727),
.B2(n_1663),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1737),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1742),
.B(n_1690),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1742),
.B(n_1689),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1780),
.B(n_1692),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1749),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1768),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1749),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1768),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1761),
.B(n_1726),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1783),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1759),
.B(n_1639),
.Y(n_1848)
);

BUFx3_ASAP7_75t_L g1849 ( 
.A(n_1760),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1814),
.A2(n_1777),
.B(n_1804),
.Y(n_1850)
);

OAI222xp33_ASAP7_75t_L g1851 ( 
.A1(n_1837),
.A2(n_1804),
.B1(n_1736),
.B2(n_1754),
.C1(n_1745),
.C2(n_1800),
.Y(n_1851)
);

AOI211xp5_ASAP7_75t_L g1852 ( 
.A1(n_1819),
.A2(n_1777),
.B(n_1747),
.C(n_1762),
.Y(n_1852)
);

OA21x2_ASAP7_75t_L g1853 ( 
.A1(n_1806),
.A2(n_1751),
.B(n_1773),
.Y(n_1853)
);

AOI33xp33_ASAP7_75t_L g1854 ( 
.A1(n_1837),
.A2(n_1783),
.A3(n_1798),
.B1(n_1795),
.B2(n_1644),
.B3(n_1754),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1819),
.A2(n_1804),
.B1(n_1796),
.B2(n_1747),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1836),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1812),
.Y(n_1857)
);

OR2x6_ASAP7_75t_L g1858 ( 
.A(n_1833),
.B(n_1736),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1836),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1820),
.A2(n_1804),
.B1(n_1796),
.B2(n_1800),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_R g1861 ( 
.A(n_1811),
.B(n_1804),
.Y(n_1861)
);

AOI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1820),
.A2(n_1795),
.B1(n_1798),
.B2(n_1763),
.C(n_1761),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1808),
.Y(n_1863)
);

OAI211xp5_ASAP7_75t_L g1864 ( 
.A1(n_1830),
.A2(n_1744),
.B(n_1796),
.C(n_1782),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1838),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1825),
.B(n_1770),
.Y(n_1866)
);

OAI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1830),
.A2(n_1736),
.B1(n_1792),
.B2(n_1790),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1817),
.B(n_1790),
.Y(n_1868)
);

INVxp67_ASAP7_75t_L g1869 ( 
.A(n_1846),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1817),
.B(n_1763),
.Y(n_1870)
);

AOI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1835),
.A2(n_1752),
.B1(n_1779),
.B2(n_1778),
.C(n_1785),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1842),
.Y(n_1872)
);

INVxp33_ASAP7_75t_L g1873 ( 
.A(n_1835),
.Y(n_1873)
);

AOI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1841),
.A2(n_1752),
.B1(n_1779),
.B2(n_1778),
.C(n_1756),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1844),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1839),
.B(n_1740),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1816),
.B(n_1840),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1841),
.A2(n_1778),
.B1(n_1757),
.B2(n_1758),
.C(n_1766),
.Y(n_1878)
);

INVx2_ASAP7_75t_SL g1879 ( 
.A(n_1810),
.Y(n_1879)
);

NAND4xp25_ASAP7_75t_SL g1880 ( 
.A(n_1813),
.B(n_1731),
.C(n_1693),
.D(n_1699),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1844),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_R g1882 ( 
.A(n_1848),
.B(n_1728),
.Y(n_1882)
);

OAI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1845),
.A2(n_1638),
.B(n_1736),
.Y(n_1883)
);

NOR4xp25_ASAP7_75t_SL g1884 ( 
.A(n_1843),
.B(n_1802),
.C(n_1762),
.D(n_1801),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1826),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1847),
.A2(n_1787),
.B1(n_1786),
.B2(n_1784),
.C(n_1789),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1816),
.B(n_1755),
.Y(n_1887)
);

OAI31xp33_ASAP7_75t_L g1888 ( 
.A1(n_1832),
.A2(n_1694),
.A3(n_1770),
.B(n_1802),
.Y(n_1888)
);

OAI221xp5_ASAP7_75t_L g1889 ( 
.A1(n_1848),
.A2(n_1736),
.B1(n_1792),
.B2(n_1803),
.C(n_1805),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1832),
.A2(n_1792),
.B1(n_1667),
.B2(n_1788),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1808),
.Y(n_1891)
);

AOI211xp5_ASAP7_75t_L g1892 ( 
.A1(n_1813),
.A2(n_1767),
.B(n_1799),
.C(n_1797),
.Y(n_1892)
);

NOR2x1_ASAP7_75t_SL g1893 ( 
.A(n_1833),
.B(n_1792),
.Y(n_1893)
);

NAND2xp33_ASAP7_75t_R g1894 ( 
.A(n_1884),
.B(n_1810),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1863),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1853),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1856),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1863),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1866),
.B(n_1834),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1882),
.B(n_1675),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1859),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1865),
.Y(n_1902)
);

BUFx8_ASAP7_75t_L g1903 ( 
.A(n_1864),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1872),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1875),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1881),
.Y(n_1906)
);

OR2x6_ASAP7_75t_L g1907 ( 
.A(n_1858),
.B(n_1809),
.Y(n_1907)
);

OR2x6_ASAP7_75t_L g1908 ( 
.A(n_1858),
.B(n_1809),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1891),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1873),
.B(n_1824),
.Y(n_1910)
);

CKINVDCx14_ASAP7_75t_R g1911 ( 
.A(n_1885),
.Y(n_1911)
);

NAND3xp33_ASAP7_75t_L g1912 ( 
.A(n_1852),
.B(n_1796),
.C(n_1826),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1879),
.B(n_1807),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1887),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1869),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1888),
.B(n_1828),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1877),
.B(n_1828),
.Y(n_1917)
);

BUFx2_ASAP7_75t_L g1918 ( 
.A(n_1858),
.Y(n_1918)
);

NOR2x1p5_ASAP7_75t_L g1919 ( 
.A(n_1885),
.B(n_1849),
.Y(n_1919)
);

OA21x2_ASAP7_75t_L g1920 ( 
.A1(n_1878),
.A2(n_1775),
.B(n_1774),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1868),
.B(n_1824),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1862),
.B(n_1870),
.Y(n_1922)
);

OA21x2_ASAP7_75t_L g1923 ( 
.A1(n_1874),
.A2(n_1775),
.B(n_1772),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1912),
.A2(n_1850),
.B1(n_1860),
.B2(n_1855),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1896),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1919),
.B(n_1892),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1919),
.B(n_1893),
.Y(n_1927)
);

INVx5_ASAP7_75t_L g1928 ( 
.A(n_1907),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1922),
.B(n_1871),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1912),
.A2(n_1860),
.B1(n_1855),
.B2(n_1867),
.Y(n_1930)
);

OAI31xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1916),
.A2(n_1867),
.A3(n_1880),
.B(n_1883),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1897),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1901),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1911),
.B(n_1675),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1902),
.Y(n_1935)
);

OAI211xp5_ASAP7_75t_SL g1936 ( 
.A1(n_1900),
.A2(n_1854),
.B(n_1909),
.C(n_1889),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1909),
.B(n_1886),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1902),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1915),
.B(n_1818),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1899),
.B(n_1918),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1918),
.B(n_1907),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1907),
.B(n_1825),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1921),
.B(n_1827),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1904),
.B(n_1818),
.Y(n_1944)
);

NOR2xp33_ASAP7_75t_L g1945 ( 
.A(n_1910),
.B(n_1827),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1907),
.B(n_1908),
.Y(n_1946)
);

NAND2xp33_ASAP7_75t_R g1947 ( 
.A(n_1908),
.B(n_1846),
.Y(n_1947)
);

AOI221xp5_ASAP7_75t_L g1948 ( 
.A1(n_1895),
.A2(n_1851),
.B1(n_1823),
.B2(n_1822),
.C(n_1815),
.Y(n_1948)
);

NAND2x1_ASAP7_75t_L g1949 ( 
.A(n_1908),
.B(n_1857),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1908),
.B(n_1876),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_1898),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1951),
.B(n_1917),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1929),
.B(n_1914),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1951),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1929),
.B(n_1917),
.Y(n_1955)
);

INVx4_ASAP7_75t_L g1956 ( 
.A(n_1928),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1937),
.B(n_1923),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1927),
.B(n_1913),
.Y(n_1958)
);

INVxp67_ASAP7_75t_SL g1959 ( 
.A(n_1947),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1932),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1940),
.Y(n_1961)
);

OAI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1948),
.A2(n_1861),
.B1(n_1894),
.B2(n_1890),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1933),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1925),
.Y(n_1964)
);

NOR2x1p5_ASAP7_75t_L g1965 ( 
.A(n_1926),
.B(n_1831),
.Y(n_1965)
);

NOR2xp67_ASAP7_75t_L g1966 ( 
.A(n_1928),
.B(n_1905),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1934),
.B(n_1829),
.Y(n_1967)
);

INVx2_ASAP7_75t_SL g1968 ( 
.A(n_1928),
.Y(n_1968)
);

NAND2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1926),
.B(n_1854),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1945),
.B(n_1943),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1928),
.B(n_1923),
.Y(n_1971)
);

NAND3xp33_ASAP7_75t_L g1972 ( 
.A(n_1931),
.B(n_1903),
.C(n_1923),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1936),
.B(n_1829),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1939),
.B(n_1821),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1933),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1939),
.B(n_1937),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1928),
.B(n_1950),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1931),
.B(n_1944),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1928),
.B(n_1906),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1935),
.Y(n_1980)
);

INVx4_ASAP7_75t_L g1981 ( 
.A(n_1956),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1959),
.B(n_1928),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1956),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1961),
.B(n_1946),
.Y(n_1984)
);

AND2x4_ASAP7_75t_SL g1985 ( 
.A(n_1954),
.B(n_1941),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1957),
.B(n_1938),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1961),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1977),
.B(n_1946),
.Y(n_1988)
);

NAND3xp33_ASAP7_75t_L g1989 ( 
.A(n_1969),
.B(n_1924),
.C(n_1948),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1960),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1971),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1971),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1952),
.Y(n_1993)
);

NOR2xp33_ASAP7_75t_L g1994 ( 
.A(n_1967),
.B(n_1936),
.Y(n_1994)
);

NOR2x1_ASAP7_75t_L g1995 ( 
.A(n_1972),
.B(n_1949),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1960),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1964),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1963),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1969),
.A2(n_1924),
.B1(n_1930),
.B2(n_1903),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1963),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1975),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1977),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1958),
.B(n_1941),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1978),
.A2(n_1930),
.B1(n_1903),
.B2(n_1920),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1966),
.B(n_1942),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1975),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1952),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1973),
.B(n_1938),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1958),
.B(n_1942),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1987),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1987),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1987),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1985),
.Y(n_2013)
);

NAND2x1_ASAP7_75t_L g2014 ( 
.A(n_2005),
.B(n_1956),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1989),
.A2(n_1962),
.B1(n_1965),
.B2(n_1903),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1993),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1993),
.Y(n_2017)
);

INVxp67_ASAP7_75t_L g2018 ( 
.A(n_2002),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1989),
.B(n_1953),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1986),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1986),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1985),
.Y(n_2022)
);

OAI22xp33_ASAP7_75t_SL g2023 ( 
.A1(n_1995),
.A2(n_1968),
.B1(n_1976),
.B2(n_1955),
.Y(n_2023)
);

AOI21xp5_ASAP7_75t_L g2024 ( 
.A1(n_1999),
.A2(n_1968),
.B(n_1970),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1986),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1990),
.Y(n_2026)
);

OAI22xp5_ASAP7_75t_SL g2027 ( 
.A1(n_1999),
.A2(n_1942),
.B1(n_1920),
.B2(n_1980),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1990),
.Y(n_2028)
);

AOI21xp33_ASAP7_75t_SL g2029 ( 
.A1(n_1994),
.A2(n_1942),
.B(n_1979),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1996),
.Y(n_2030)
);

INVxp67_ASAP7_75t_L g2031 ( 
.A(n_1984),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_2007),
.B(n_1974),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2013),
.B(n_1985),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_2019),
.B(n_2007),
.Y(n_2034)
);

NOR2x1p5_ASAP7_75t_SL g2035 ( 
.A(n_2022),
.B(n_1991),
.Y(n_2035)
);

INVxp67_ASAP7_75t_L g2036 ( 
.A(n_2016),
.Y(n_2036)
);

INVx2_ASAP7_75t_SL g2037 ( 
.A(n_2014),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2017),
.Y(n_2038)
);

INVx3_ASAP7_75t_SL g2039 ( 
.A(n_2010),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_2032),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2018),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_2018),
.B(n_2002),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2031),
.B(n_1984),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_2029),
.B(n_1988),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2024),
.B(n_1984),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2011),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2012),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2020),
.Y(n_2048)
);

OAI211xp5_ASAP7_75t_L g2049 ( 
.A1(n_2045),
.A2(n_2019),
.B(n_2015),
.C(n_2004),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2034),
.B(n_2024),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_2043),
.B(n_2008),
.Y(n_2051)
);

NAND4xp25_ASAP7_75t_L g2052 ( 
.A(n_2034),
.B(n_2004),
.C(n_1995),
.D(n_1982),
.Y(n_2052)
);

OAI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_2040),
.A2(n_2023),
.B(n_1982),
.Y(n_2053)
);

NAND3xp33_ASAP7_75t_L g2054 ( 
.A(n_2033),
.B(n_1982),
.C(n_2002),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_R g2055 ( 
.A(n_2037),
.B(n_1983),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_SL g2056 ( 
.A(n_2033),
.B(n_2037),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2044),
.A2(n_2027),
.B1(n_1988),
.B2(n_2003),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2042),
.B(n_2041),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_2039),
.A2(n_1988),
.B1(n_2003),
.B2(n_2009),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_2036),
.A2(n_2008),
.B(n_1983),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_2042),
.A2(n_2025),
.B(n_2021),
.Y(n_2061)
);

AOI211xp5_ASAP7_75t_L g2062 ( 
.A1(n_2039),
.A2(n_2026),
.B(n_2030),
.C(n_2028),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_2042),
.A2(n_2003),
.B1(n_2009),
.B2(n_2041),
.Y(n_2063)
);

INVx2_ASAP7_75t_SL g2064 ( 
.A(n_2038),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2058),
.Y(n_2065)
);

INVx2_ASAP7_75t_SL g2066 ( 
.A(n_2055),
.Y(n_2066)
);

XOR2xp5_ASAP7_75t_L g2067 ( 
.A(n_2052),
.B(n_2048),
.Y(n_2067)
);

INVxp33_ASAP7_75t_SL g2068 ( 
.A(n_2056),
.Y(n_2068)
);

INVx1_ASAP7_75t_SL g2069 ( 
.A(n_2063),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2054),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2061),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2064),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_2050),
.A2(n_1983),
.B(n_1981),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2066),
.Y(n_2074)
);

NOR3xp33_ASAP7_75t_L g2075 ( 
.A(n_2065),
.B(n_2049),
.C(n_2053),
.Y(n_2075)
);

NAND2x1_ASAP7_75t_SL g2076 ( 
.A(n_2071),
.B(n_1983),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2068),
.B(n_2059),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2069),
.B(n_2051),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2072),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2068),
.B(n_2035),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_2070),
.B(n_2057),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2075),
.A2(n_2067),
.B1(n_2070),
.B2(n_2005),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2078),
.B(n_2080),
.Y(n_2083)
);

INVx1_ASAP7_75t_SL g2084 ( 
.A(n_2076),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_R g2085 ( 
.A(n_2077),
.B(n_2046),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_2074),
.Y(n_2086)
);

NAND3x2_ASAP7_75t_L g2087 ( 
.A(n_2079),
.B(n_2047),
.C(n_2005),
.Y(n_2087)
);

NOR4xp75_ASAP7_75t_L g2088 ( 
.A(n_2081),
.B(n_2060),
.C(n_2062),
.D(n_2073),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2086),
.B(n_1991),
.Y(n_2089)
);

INVxp67_ASAP7_75t_SL g2090 ( 
.A(n_2087),
.Y(n_2090)
);

OAI211xp5_ASAP7_75t_L g2091 ( 
.A1(n_2082),
.A2(n_1981),
.B(n_1998),
.C(n_1996),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_2084),
.Y(n_2092)
);

BUFx2_ASAP7_75t_L g2093 ( 
.A(n_2089),
.Y(n_2093)
);

NOR3xp33_ASAP7_75t_L g2094 ( 
.A(n_2093),
.B(n_2090),
.C(n_2083),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_2094),
.Y(n_2095)
);

NAND2x1_ASAP7_75t_SL g2096 ( 
.A(n_2094),
.B(n_2092),
.Y(n_2096)
);

OAI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2095),
.A2(n_1981),
.B1(n_2091),
.B2(n_1992),
.Y(n_2097)
);

OAI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_2096),
.A2(n_1981),
.B1(n_2088),
.B2(n_2085),
.C(n_1991),
.Y(n_2098)
);

CKINVDCx20_ASAP7_75t_R g2099 ( 
.A(n_2097),
.Y(n_2099)
);

OAI21xp5_ASAP7_75t_SL g2100 ( 
.A1(n_2098),
.A2(n_1992),
.B(n_1998),
.Y(n_2100)
);

CKINVDCx20_ASAP7_75t_R g2101 ( 
.A(n_2099),
.Y(n_2101)
);

AOI21xp5_ASAP7_75t_L g2102 ( 
.A1(n_2101),
.A2(n_2100),
.B(n_1981),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2102),
.B(n_2000),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2103),
.A2(n_1992),
.B1(n_1997),
.B2(n_2000),
.Y(n_2104)
);

AOI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_2104),
.A2(n_2005),
.B1(n_1997),
.B2(n_2001),
.Y(n_2105)
);

AOI211xp5_ASAP7_75t_L g2106 ( 
.A1(n_2105),
.A2(n_2006),
.B(n_2001),
.C(n_1997),
.Y(n_2106)
);


endmodule