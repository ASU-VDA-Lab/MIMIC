module fake_jpeg_397_n_454 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_454);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_454;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_442;
wire n_299;
wire n_300;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_48),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_61),
.Y(n_95)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_54),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_23),
.B(n_0),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_63),
.Y(n_96)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_0),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_25),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_77),
.Y(n_98)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_25),
.B(n_1),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

CKINVDCx9p33_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_21),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_57),
.A2(n_26),
.B1(n_44),
.B2(n_21),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_84),
.A2(n_107),
.B1(n_124),
.B2(n_2),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_83),
.B1(n_81),
.B2(n_76),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_91),
.A2(n_102),
.B1(n_108),
.B2(n_123),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_43),
.B1(n_38),
.B2(n_31),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_43),
.B1(n_38),
.B2(n_31),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_126),
.B1(n_134),
.B2(n_135),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_26),
.B1(n_44),
.B2(n_21),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_43),
.B1(n_38),
.B2(n_31),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_125),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_116),
.B(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_45),
.B(n_20),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_117),
.B(n_118),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_48),
.B(n_29),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_34),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_42),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_20),
.B1(n_24),
.B2(n_29),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_26),
.B1(n_42),
.B2(n_44),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_48),
.B(n_24),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_46),
.A2(n_47),
.B1(n_62),
.B2(n_51),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_50),
.B(n_36),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_130),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_70),
.B(n_36),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_79),
.A2(n_33),
.B1(n_32),
.B2(n_18),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_27),
.B1(n_42),
.B2(n_44),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_32),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_53),
.B(n_33),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_49),
.A2(n_38),
.B1(n_31),
.B2(n_40),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_54),
.A2(n_44),
.B1(n_42),
.B2(n_40),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_53),
.B(n_34),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_53),
.B(n_27),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_142),
.B(n_149),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_143),
.A2(n_110),
.B1(n_94),
.B2(n_137),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_88),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g214 ( 
.A(n_144),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_146),
.B(n_194),
.Y(n_211)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_96),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g150 ( 
.A(n_135),
.B(n_2),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_150),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_151),
.Y(n_237)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_42),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_153),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_95),
.B(n_2),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_161),
.Y(n_218)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_163),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_102),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_139),
.B1(n_128),
.B2(n_115),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_92),
.Y(n_165)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_90),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_110),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_95),
.B(n_4),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_90),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_86),
.B(n_5),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_187),
.Y(n_223)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_176),
.B(n_179),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_126),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_177)
);

OAI22x1_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_139),
.B1(n_115),
.B2(n_128),
.Y(n_199)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_181),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_89),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_189),
.Y(n_234)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_185),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_106),
.B(n_14),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g243 ( 
.A(n_184),
.B(n_13),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_87),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_98),
.B(n_7),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_106),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_136),
.B(n_121),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_112),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_113),
.A2(n_8),
.B(n_9),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_190),
.B(n_184),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_108),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_127),
.B1(n_93),
.B2(n_114),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_100),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_195),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_122),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_87),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_122),
.B(n_10),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_197),
.B(n_13),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_198),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_199),
.A2(n_232),
.B1(n_214),
.B2(n_198),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_113),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_217),
.Y(n_247)
);

AO21x2_ASAP7_75t_L g204 ( 
.A1(n_145),
.A2(n_104),
.B(n_137),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_204),
.A2(n_161),
.B1(n_158),
.B2(n_147),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_205),
.A2(n_227),
.B1(n_235),
.B2(n_165),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_142),
.A2(n_162),
.B(n_194),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_209),
.A2(n_225),
.B(n_244),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_151),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_224),
.B1(n_232),
.B2(n_238),
.Y(n_249)
);

AO22x1_ASAP7_75t_SL g221 ( 
.A1(n_186),
.A2(n_121),
.B1(n_112),
.B2(n_127),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_241),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_93),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_156),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_145),
.A2(n_100),
.B1(n_136),
.B2(n_105),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_146),
.A2(n_105),
.B1(n_88),
.B2(n_138),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_167),
.A2(n_88),
.B1(n_11),
.B2(n_13),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_164),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_197),
.A2(n_154),
.B1(n_168),
.B2(n_153),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_166),
.B1(n_172),
.B2(n_148),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_144),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_188),
.A2(n_184),
.B(n_178),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_175),
.B(n_187),
.Y(n_257)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_250),
.Y(n_293)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_251),
.Y(n_294)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_203),
.B(n_223),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_253),
.B(n_258),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_204),
.A2(n_153),
.B1(n_143),
.B2(n_179),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_263),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_255),
.A2(n_276),
.B1(n_284),
.B2(n_217),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_236),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_SL g316 ( 
.A1(n_257),
.A2(n_242),
.B(n_237),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_148),
.Y(n_258)
);

BUFx4f_ASAP7_75t_SL g260 ( 
.A(n_228),
.Y(n_260)
);

INVx13_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_262),
.B(n_266),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_204),
.A2(n_172),
.B1(n_166),
.B2(n_192),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_264),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_223),
.B(n_206),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_265),
.B(n_277),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_211),
.A2(n_157),
.B(n_180),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_272),
.B(n_236),
.Y(n_292)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_204),
.A2(n_176),
.B1(n_163),
.B2(n_152),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_270),
.A2(n_273),
.B1(n_275),
.B2(n_279),
.Y(n_323)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_230),
.Y(n_271)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_211),
.A2(n_181),
.B(n_185),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_204),
.A2(n_185),
.B1(n_171),
.B2(n_183),
.Y(n_273)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_282),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_227),
.A2(n_195),
.B1(n_174),
.B2(n_173),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_222),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_206),
.B(n_193),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_287),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_209),
.A2(n_159),
.B1(n_196),
.B2(n_229),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_218),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_289),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_231),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_214),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_285),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_229),
.A2(n_208),
.B1(n_221),
.B2(n_220),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_201),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_286),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_208),
.A2(n_221),
.B1(n_216),
.B2(n_205),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_202),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_290),
.Y(n_324)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_248),
.A2(n_216),
.B1(n_225),
.B2(n_246),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_291),
.A2(n_298),
.B1(n_299),
.B2(n_263),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_292),
.A2(n_283),
.B(n_260),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_226),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_296),
.A2(n_266),
.A3(n_283),
.B1(n_287),
.B2(n_269),
.C1(n_250),
.C2(n_251),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_248),
.A2(n_243),
.B1(n_200),
.B2(n_199),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_243),
.B1(n_200),
.B2(n_236),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_301),
.B(n_324),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_242),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_303),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_259),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_307),
.B(n_326),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_233),
.C(n_239),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_317),
.C(n_301),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_245),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_316),
.Y(n_357)
);

NAND2x1p5_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_233),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_314),
.A2(n_261),
.B(n_252),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_247),
.B(n_219),
.C(n_242),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_219),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_228),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_237),
.Y(n_326)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_307),
.A2(n_272),
.B(n_268),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_329),
.A2(n_334),
.B(n_340),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_295),
.A2(n_284),
.B1(n_249),
.B2(n_255),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_330),
.A2(n_337),
.B1(n_338),
.B2(n_358),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_331),
.B(n_336),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_343),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_307),
.A2(n_273),
.B(n_254),
.Y(n_334)
);

AOI221xp5_ASAP7_75t_L g336 ( 
.A1(n_292),
.A2(n_321),
.B1(n_304),
.B2(n_309),
.C(n_297),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_249),
.B1(n_270),
.B2(n_275),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_290),
.B1(n_281),
.B2(n_264),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_345),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_304),
.A2(n_271),
.B(n_212),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_341),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_212),
.C(n_215),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_344),
.C(n_317),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_215),
.C(n_286),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_274),
.B(n_267),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_L g374 ( 
.A1(n_348),
.A2(n_340),
.B(n_354),
.Y(n_374)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_349),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_319),
.B(n_260),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_351),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_302),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_355),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_291),
.B(n_283),
.Y(n_354)
);

AO22x1_ASAP7_75t_L g383 ( 
.A1(n_354),
.A2(n_298),
.B1(n_323),
.B2(n_313),
.Y(n_383)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_323),
.A2(n_260),
.B1(n_267),
.B2(n_238),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_328),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_353),
.A2(n_304),
.B(n_314),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_365),
.A2(n_374),
.B(n_353),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_321),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_368),
.C(n_373),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_296),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_319),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_369),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_350),
.B(n_309),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_SL g391 ( 
.A(n_372),
.B(n_352),
.C(n_355),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_305),
.C(n_299),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_303),
.C(n_312),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_379),
.C(n_380),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_347),
.B(n_303),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_376),
.A2(n_382),
.B1(n_306),
.B2(n_357),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_312),
.C(n_322),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_322),
.C(n_320),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_335),
.B(n_320),
.C(n_313),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_349),
.C(n_341),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_356),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_331),
.B(n_337),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_384),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_400),
.C(n_360),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_378),
.A2(n_330),
.B1(n_334),
.B2(n_335),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_389),
.Y(n_420)
);

NAND4xp25_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_391),
.C(n_404),
.D(n_384),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_371),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_363),
.A2(n_354),
.B1(n_357),
.B2(n_333),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_393),
.A2(n_383),
.B1(n_378),
.B2(n_377),
.Y(n_419)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_394),
.Y(n_414)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_398),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_366),
.B(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_381),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_401),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_348),
.C(n_345),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_333),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_402),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_403),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_417),
.C(n_412),
.Y(n_425)
);

AOI31xp33_ASAP7_75t_L g430 ( 
.A1(n_409),
.A2(n_404),
.A3(n_400),
.B(n_361),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_390),
.B(n_364),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_412),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_373),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_368),
.C(n_380),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_418),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_359),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_419),
.A2(n_383),
.B1(n_420),
.B2(n_389),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_377),
.C(n_361),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_421),
.B(n_386),
.C(n_399),
.Y(n_424)
);

AO221x1_ASAP7_75t_L g422 ( 
.A1(n_407),
.A2(n_397),
.B1(n_387),
.B2(n_363),
.C(n_391),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_425),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_SL g423 ( 
.A1(n_420),
.A2(n_377),
.B(n_393),
.C(n_388),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_423),
.A2(n_408),
.B(n_365),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_431),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_413),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_427),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_401),
.C(n_396),
.Y(n_427)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_430),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_402),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_419),
.Y(n_433)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_433),
.A2(n_438),
.B(n_394),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_421),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_437),
.A2(n_429),
.B(n_428),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_423),
.A2(n_416),
.B1(n_398),
.B2(n_411),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_440),
.A2(n_423),
.B(n_411),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_442),
.Y(n_448)
);

AO22x1_ASAP7_75t_L g442 ( 
.A1(n_436),
.A2(n_416),
.B1(n_423),
.B2(n_414),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_443),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_444),
.B(n_445),
.Y(n_446)
);

A2O1A1Ixp33_ASAP7_75t_SL g445 ( 
.A1(n_439),
.A2(n_427),
.B(n_415),
.C(n_395),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_435),
.C(n_434),
.Y(n_449)
);

OAI311xp33_ASAP7_75t_L g451 ( 
.A1(n_449),
.A2(n_450),
.A3(n_447),
.B1(n_418),
.C1(n_315),
.Y(n_451)
);

O2A1O1Ixp33_ASAP7_75t_SL g450 ( 
.A1(n_446),
.A2(n_438),
.B(n_440),
.C(n_433),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_451),
.A2(n_358),
.B(n_300),
.Y(n_452)
);

AO21x1_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_300),
.B(n_311),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_315),
.Y(n_454)
);


endmodule