module fake_netlist_1_9468_n_26 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_26);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_6), .Y(n_11) );
AND2x4_ASAP7_75t_L g12 ( .A(n_3), .B(n_0), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
BUFx3_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_14), .B(n_0), .Y(n_18) );
AOI211xp5_ASAP7_75t_L g19 ( .A1(n_18), .A2(n_13), .B(n_12), .C(n_14), .Y(n_19) );
OAI221xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_17), .B1(n_15), .B2(n_16), .C(n_11), .Y(n_20) );
INVxp67_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_17), .B1(n_12), .B2(n_4), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_22), .B(n_5), .Y(n_23) );
NAND4xp25_ASAP7_75t_L g24 ( .A(n_23), .B(n_8), .C(n_9), .D(n_10), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
endmodule