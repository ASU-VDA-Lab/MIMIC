module real_jpeg_21590_n_17 (n_8, n_0, n_2, n_338, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_338;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_1),
.A2(n_39),
.B1(n_71),
.B2(n_72),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_1),
.A2(n_39),
.B1(n_49),
.B2(n_50),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_2),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_71),
.B1(n_72),
.B2(n_118),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_118),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_118),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_3),
.A2(n_53),
.B1(n_71),
.B2(n_72),
.Y(n_250)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_50),
.B(n_67),
.C(n_103),
.D(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_4),
.B(n_48),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_4),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_4),
.A2(n_124),
.B(n_126),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_4),
.A2(n_36),
.B(n_43),
.C(n_160),
.D(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_4),
.B(n_36),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_40),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_4),
.A2(n_35),
.B(n_37),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_141),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_71),
.B1(n_72),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_5),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_123),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_123),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_123),
.Y(n_261)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_7),
.B(n_72),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_7),
.B(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_7),
.Y(n_135)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_7),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_7),
.A2(n_125),
.B1(n_171),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_8),
.A2(n_64),
.B1(n_71),
.B2(n_72),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_8),
.A2(n_36),
.B1(n_37),
.B2(n_64),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_10),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_10),
.A2(n_71),
.B1(n_72),
.B2(n_85),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_85),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_85),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_11),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_11),
.A2(n_71),
.B1(n_72),
.B2(n_106),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_106),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_106),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_13),
.A2(n_29),
.B1(n_71),
.B2(n_72),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_13),
.A2(n_29),
.B1(n_49),
.B2(n_50),
.Y(n_252)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_91),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_77),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_77),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_54),
.B1(n_55),
.B2(n_76),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_21),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_41),
.B2(n_42),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_25),
.A2(n_31),
.B1(n_34),
.B2(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_32),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_27),
.A2(n_32),
.B(n_141),
.C(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_30),
.A2(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_30),
.B(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_31),
.A2(n_34),
.B1(n_63),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_31),
.A2(n_34),
.B1(n_230),
.B2(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_31),
.A2(n_221),
.B(n_261),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_34),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_34),
.A2(n_84),
.B(n_231),
.Y(n_303)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_44),
.B(n_47),
.C(n_48),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_40),
.B(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_48),
.B(n_51),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_43),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_43),
.A2(n_48),
.B1(n_258),
.B2(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_43),
.A2(n_48),
.B1(n_90),
.B2(n_277),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_44),
.B(n_50),
.Y(n_168)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_47),
.A2(n_49),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_68),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.C(n_65),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_57),
.B1(n_65),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_58),
.A2(n_60),
.B1(n_180),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_58),
.A2(n_216),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_60),
.B(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_60),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_60),
.A2(n_181),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_62),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_65),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_74),
.B(n_75),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_66),
.A2(n_74),
.B1(n_117),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_66),
.A2(n_158),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_66),
.A2(n_74),
.B1(n_213),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_66),
.A2(n_74),
.B1(n_243),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_66),
.A2(n_74),
.B1(n_252),
.B2(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_67),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_67),
.A2(n_70),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_72),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_71),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_117),
.B(n_119),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_74),
.B(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_74),
.A2(n_119),
.B(n_213),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_75),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.C(n_86),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_322),
.Y(n_328)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.C(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_83),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_83),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_86),
.B(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI321xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_319),
.A3(n_329),
.B1(n_334),
.B2(n_335),
.C(n_337),
.Y(n_93)
);

AOI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_269),
.A3(n_307),
.B1(n_313),
.B2(n_318),
.C(n_338),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_224),
.C(n_265),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_195),
.B(n_223),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_174),
.B(n_194),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_152),
.B(n_173),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_128),
.B(n_151),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_101),
.B(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_107),
.B1(n_108),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_104),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_121),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_116),
.C(n_121),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_124),
.B(n_126),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_124),
.A2(n_135),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_124),
.A2(n_206),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_124),
.A2(n_135),
.B1(n_241),
.B2(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_124),
.A2(n_143),
.B(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_127),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_138),
.B(n_150),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_136),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_141),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_145),
.B(n_149),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_142),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_144),
.B(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_143),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_153),
.B(n_154),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_165),
.B2(n_172),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_163),
.B2(n_164),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_164),
.C(n_172),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_160),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_161),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_169),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_188),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_190),
.C(n_192),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_183),
.B2(n_187),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_184),
.C(n_185),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_183),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_189),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_196),
.B(n_197),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_210),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_199),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_199),
.B(n_209),
.C(n_210),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_204),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_207),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_225),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_245),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_226),
.B(n_245),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_237),
.C(n_244),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_236),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_242),
.Y(n_254)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_263),
.B2(n_264),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_253),
.C(n_264),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_251),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_259),
.C(n_262),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_256),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_267),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_287),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_270),
.B(n_287),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_280),
.C(n_286),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_271),
.A2(n_272),
.B1(n_280),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_285),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_281),
.A2(n_282),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_299),
.B(n_303),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_283),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_283),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_284),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_305),
.B2(n_306),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_297),
.B2(n_298),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_298),
.C(n_306),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_295),
.B(n_296),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_295),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_296),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_296),
.A2(n_321),
.B1(n_325),
.B2(n_333),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_310),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_327),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.C(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_321),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);


endmodule