module fake_jpeg_12848_n_139 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_20),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_29),
.A2(n_31),
.B1(n_37),
.B2(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_30),
.B(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_18),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_34),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_5),
.C(n_7),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_35),
.C(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_12),
.B(n_8),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_41),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_18),
.A2(n_22),
.B1(n_12),
.B2(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_18),
.A2(n_22),
.B1(n_26),
.B2(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_24),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g47 ( 
.A(n_12),
.B(n_19),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_19),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_19),
.A2(n_26),
.B1(n_15),
.B2(n_24),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_26),
.B1(n_15),
.B2(n_27),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_54),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_40),
.C(n_51),
.Y(n_79)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_50),
.B1(n_57),
.B2(n_73),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_72),
.Y(n_93)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_35),
.B(n_48),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_29),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_31),
.B(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_91),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_90),
.B1(n_89),
.B2(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_94),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_71),
.C(n_64),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_60),
.B1(n_65),
.B2(n_69),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_60),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_69),
.B1(n_58),
.B2(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_98),
.B1(n_86),
.B2(n_88),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_92),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_73),
.B1(n_29),
.B2(n_77),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_106),
.Y(n_115)
);

XOR2x2_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_115),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_93),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_118),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_85),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_126),
.B1(n_117),
.B2(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_105),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_119),
.A2(n_110),
.B1(n_101),
.B2(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_104),
.B1(n_100),
.B2(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_129),
.B(n_96),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_124),
.C(n_123),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_100),
.B(n_127),
.C(n_121),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_136),
.B(n_133),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_126),
.C(n_130),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_124),
.Y(n_139)
);


endmodule