module fake_jpeg_24487_n_323 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_6),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_8),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_49),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_37),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_63),
.B(n_65),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_29),
.B1(n_25),
.B2(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_56),
.B1(n_70),
.B2(n_71),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_54),
.A2(n_57),
.B1(n_85),
.B2(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_43),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_66),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_25),
.B1(n_29),
.B2(n_37),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_26),
.B1(n_36),
.B2(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_58),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_32),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_75),
.B1(n_77),
.B2(n_81),
.Y(n_90)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_27),
.B1(n_36),
.B2(n_26),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_27),
.B1(n_36),
.B2(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_76),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_30),
.B1(n_19),
.B2(n_21),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_24),
.B1(n_19),
.B2(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_0),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_33),
.B1(n_28),
.B2(n_22),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_0),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_20),
.B1(n_38),
.B2(n_2),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_20),
.B1(n_11),
.B2(n_17),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_20),
.B1(n_38),
.B2(n_11),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_38),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_93),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_95),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_50),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_103),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_1),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_86),
.B1(n_56),
.B2(n_53),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_116),
.B1(n_69),
.B2(n_80),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_119),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_112),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_118),
.B1(n_50),
.B2(n_59),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

CKINVDCx10_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_7),
.C(n_16),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_0),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_63),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_120),
.Y(n_143)
);

CKINVDCx9p33_ASAP7_75t_R g117 ( 
.A(n_62),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_71),
.B1(n_82),
.B2(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_61),
.B(n_10),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_52),
.B(n_1),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_13),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_122),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_123),
.B(n_131),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_128),
.B1(n_107),
.B2(n_89),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_74),
.B1(n_60),
.B2(n_79),
.Y(n_128)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_16),
.Y(n_131)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_60),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_150),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_69),
.C(n_80),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_105),
.C(n_109),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_144),
.A2(n_108),
.B1(n_96),
.B2(n_119),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_80),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_149),
.Y(n_165)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_113),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_96),
.B(n_13),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_95),
.B(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_50),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_152),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_59),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_153),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_121),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_156),
.A2(n_160),
.B1(n_174),
.B2(n_148),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_89),
.B1(n_118),
.B2(n_90),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_104),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_171),
.B(n_123),
.Y(n_199)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_173),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_115),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_166),
.A2(n_185),
.B(n_134),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_167),
.A2(n_175),
.B1(n_185),
.B2(n_171),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_176),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_144),
.B1(n_90),
.B2(n_132),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_125),
.A2(n_117),
.B1(n_98),
.B2(n_88),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_183),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_114),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_186),
.C(n_134),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_110),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_184),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_149),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_122),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g185 ( 
.A1(n_129),
.A2(n_113),
.B1(n_91),
.B2(n_154),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_135),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_124),
.B(n_78),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_200),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_206),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_124),
.B(n_131),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_213),
.B(n_185),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_211),
.C(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_170),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_203),
.Y(n_242)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_210),
.Y(n_225)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_161),
.B(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_215),
.B(n_174),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_212),
.C(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_175),
.A2(n_129),
.B(n_141),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_129),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_141),
.B(n_127),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_91),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_91),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_167),
.B1(n_210),
.B2(n_156),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_161),
.B(n_130),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_227),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_208),
.B(n_193),
.Y(n_246)
);

BUFx12f_ASAP7_75t_SL g226 ( 
.A(n_213),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_228),
.B1(n_193),
.B2(n_200),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_166),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_233),
.B1(n_235),
.B2(n_226),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_239),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_235),
.B1(n_219),
.B2(n_197),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_215),
.A2(n_160),
.B1(n_173),
.B2(n_166),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_168),
.B1(n_164),
.B2(n_169),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_196),
.B1(n_190),
.B2(n_195),
.Y(n_256)
);

OAI22x1_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_182),
.B1(n_172),
.B2(n_176),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_182),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_164),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_256),
.B(n_234),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_209),
.C(n_212),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_238),
.C(n_236),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_198),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_241),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_216),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_251),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_223),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_191),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_242),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_192),
.B1(n_195),
.B2(n_199),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_225),
.B1(n_228),
.B2(n_231),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_192),
.B1(n_187),
.B2(n_188),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_220),
.A2(n_172),
.B1(n_180),
.B2(n_105),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_260),
.A2(n_243),
.B1(n_147),
.B2(n_109),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_225),
.A2(n_172),
.B1(n_206),
.B2(n_162),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_279),
.B1(n_253),
.B2(n_246),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_276),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_272),
.C(n_275),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_230),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_273),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_221),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_227),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_232),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_257),
.B(n_262),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_165),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_277),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_258),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_289),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_266),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_265),
.A2(n_261),
.B(n_248),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_287),
.B(n_12),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_250),
.C(n_256),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_270),
.C(n_275),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_239),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_153),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_294),
.B(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_270),
.C(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_286),
.B(n_269),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_297),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_292),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_276),
.C(n_153),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_301),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_282),
.B(n_288),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_147),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_281),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_4),
.C(n_5),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_285),
.Y(n_307)
);

NOR4xp25_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_310),
.C(n_299),
.D(n_7),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_299),
.C(n_293),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_303),
.B(n_17),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_313),
.A2(n_304),
.A3(n_305),
.B1(n_4),
.B2(n_5),
.C1(n_13),
.C2(n_17),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_15),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_314),
.C(n_312),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_318),
.B(n_2),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_320),
.B(n_2),
.C(n_3),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_3),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_322),
.Y(n_323)
);


endmodule