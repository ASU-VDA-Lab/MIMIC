module fake_jpeg_10324_n_59 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_21),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_32),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_31),
.B(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_22),
.B1(n_15),
.B2(n_16),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_29),
.B1(n_26),
.B2(n_6),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_26),
.B1(n_5),
.B2(n_6),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_4),
.B(n_5),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_13),
.C(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_39),
.B1(n_50),
.B2(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_49),
.Y(n_57)
);

AOI21x1_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_52),
.B(n_43),
.Y(n_58)
);

AOI321xp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_48),
.A3(n_40),
.B1(n_54),
.B2(n_51),
.C(n_46),
.Y(n_59)
);


endmodule