module fake_jpeg_20508_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx16_ASAP7_75t_R g6 ( 
.A(n_0),
.Y(n_6)
);

INVx6_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_10),
.B(n_4),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_14),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g13 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_15),
.B1(n_6),
.B2(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

OA22x2_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_7),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_18),
.A2(n_20),
.B1(n_15),
.B2(n_9),
.Y(n_23)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_20),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_23),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_29),
.B(n_25),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_22),
.B1(n_21),
.B2(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_31),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_27),
.B(n_21),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_29),
.B(n_15),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_9),
.Y(n_34)
);


endmodule