module real_jpeg_1274_n_29 (n_17, n_8, n_0, n_157, n_21, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_24, n_6, n_159, n_28, n_153, n_151, n_161, n_23, n_11, n_14, n_160, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_158, n_16, n_15, n_13, n_155, n_29);

input n_17;
input n_8;
input n_0;
input n_157;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_24;
input n_6;
input n_159;
input n_28;
input n_153;
input n_151;
input n_161;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_158;
input n_16;
input n_15;
input n_13;
input n_155;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_0),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_2),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_50),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_5),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_7),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_8),
.Y(n_145)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_68),
.B1(n_100),
.B2(n_103),
.Y(n_67)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_12),
.B(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_13),
.B(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_13),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_14),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_15),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_72),
.C(n_87),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_17),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_19),
.A2(n_78),
.B(n_82),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_20),
.A2(n_31),
.B1(n_141),
.B2(n_144),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_33),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_20),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_20),
.A2(n_142),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

AO22x1_ASAP7_75t_L g72 ( 
.A1(n_21),
.A2(n_73),
.B1(n_76),
.B2(n_86),
.Y(n_72)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_22),
.B(n_70),
.C(n_94),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_23),
.B(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_23),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_24),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_146),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_40),
.B(n_140),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_35),
.B(n_145),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_36),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_36),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_36),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_36),
.B(n_139),
.Y(n_138)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g93 ( 
.A(n_39),
.Y(n_93)
);

MAJx2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_136),
.C(n_137),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_135),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_43),
.B(n_46),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B(n_53),
.C(n_134),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_52),
.B(n_149),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_130),
.C(n_131),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_129),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_56),
.B(n_60),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_99),
.Y(n_98)
);

OAI221xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_66),
.B1(n_67),
.B2(n_105),
.C(n_119),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_96),
.C(n_97),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_89),
.C(n_90),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_83),
.Y(n_82)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_84),
.C(n_85),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_82),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_114),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_120),
.A3(n_121),
.B1(n_124),
.B2(n_125),
.C1(n_128),
.C2(n_161),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.C(n_111),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_151),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_152),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_153),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_154),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_155),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_156),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_157),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_158),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_159),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_160),
.Y(n_118)
);


endmodule