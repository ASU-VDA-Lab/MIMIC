module real_aes_2988_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_792;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g530 ( .A(n_0), .B(n_227), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_1), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g161 ( .A(n_2), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_3), .B(n_533), .Y(n_552) );
NAND2xp33_ASAP7_75t_SL g523 ( .A(n_4), .B(n_182), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_5), .B(n_195), .Y(n_218) );
INVx1_ASAP7_75t_L g515 ( .A(n_6), .Y(n_515) );
INVx1_ASAP7_75t_L g252 ( .A(n_7), .Y(n_252) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_9), .Y(n_269) );
AND2x2_ASAP7_75t_L g550 ( .A(n_10), .B(n_151), .Y(n_550) );
INVx2_ASAP7_75t_L g152 ( .A(n_11), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_12), .Y(n_114) );
INVx1_ASAP7_75t_L g228 ( .A(n_13), .Y(n_228) );
AOI221x1_ASAP7_75t_L g518 ( .A1(n_14), .A2(n_184), .B1(n_519), .B2(n_521), .C(n_522), .Y(n_518) );
OAI22xp5_ASAP7_75t_SL g804 ( .A1(n_14), .A2(n_58), .B1(n_805), .B2(n_806), .Y(n_804) );
INVxp67_ASAP7_75t_L g806 ( .A(n_14), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_15), .B(n_533), .Y(n_586) );
NOR2xp33_ASAP7_75t_SL g109 ( .A(n_16), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g127 ( .A(n_16), .Y(n_127) );
INVx1_ASAP7_75t_L g225 ( .A(n_17), .Y(n_225) );
INVx1_ASAP7_75t_SL g173 ( .A(n_18), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_19), .B(n_176), .Y(n_198) );
AOI33xp33_ASAP7_75t_L g243 ( .A1(n_20), .A2(n_48), .A3(n_158), .B1(n_169), .B2(n_244), .B3(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_21), .A2(n_521), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_22), .B(n_227), .Y(n_555) );
AOI221xp5_ASAP7_75t_SL g595 ( .A1(n_23), .A2(n_39), .B1(n_521), .B2(n_533), .C(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g262 ( .A(n_24), .Y(n_262) );
OR2x2_ASAP7_75t_L g153 ( .A(n_25), .B(n_93), .Y(n_153) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_25), .A2(n_93), .B(n_152), .Y(n_186) );
INVxp67_ASAP7_75t_L g517 ( .A(n_26), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_27), .B(n_230), .Y(n_590) );
AND2x2_ASAP7_75t_L g544 ( .A(n_28), .B(n_150), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_29), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_30), .B(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_31), .A2(n_521), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_32), .B(n_230), .Y(n_597) );
AND2x2_ASAP7_75t_L g163 ( .A(n_33), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g168 ( .A(n_33), .Y(n_168) );
AND2x2_ASAP7_75t_L g182 ( .A(n_33), .B(n_161), .Y(n_182) );
NOR3xp33_ASAP7_75t_L g111 ( .A(n_34), .B(n_112), .C(n_114), .Y(n_111) );
OR2x6_ASAP7_75t_L g125 ( .A(n_34), .B(n_126), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_35), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_36), .B(n_156), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_37), .A2(n_185), .B1(n_191), .B2(n_195), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_38), .B(n_200), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_40), .A2(n_85), .B1(n_166), .B2(n_521), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_41), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_42), .B(n_227), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_43), .B(n_202), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_44), .B(n_176), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_45), .Y(n_194) );
AND2x2_ASAP7_75t_L g534 ( .A(n_46), .B(n_150), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_47), .B(n_150), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_49), .B(n_176), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_50), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_50), .A2(n_63), .B1(n_441), .B2(n_817), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_51), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g159 ( .A(n_52), .Y(n_159) );
INVx1_ASAP7_75t_L g178 ( .A(n_52), .Y(n_178) );
AOI22x1_ASAP7_75t_L g131 ( .A1(n_53), .A2(n_132), .B1(n_133), .B2(n_134), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_53), .Y(n_132) );
AND2x2_ASAP7_75t_L g294 ( .A(n_54), .B(n_150), .Y(n_294) );
AOI221xp5_ASAP7_75t_L g250 ( .A1(n_55), .A2(n_78), .B1(n_156), .B2(n_166), .C(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_56), .B(n_156), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_57), .B(n_533), .Y(n_543) );
INVx1_ASAP7_75t_L g805 ( .A(n_58), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_59), .B(n_185), .Y(n_271) );
AOI21xp5_ASAP7_75t_SL g207 ( .A1(n_60), .A2(n_166), .B(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g571 ( .A(n_61), .B(n_150), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_62), .B(n_230), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_63), .Y(n_817) );
INVx1_ASAP7_75t_L g221 ( .A(n_64), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_65), .B(n_227), .Y(n_569) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_66), .B(n_151), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_67), .A2(n_521), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g292 ( .A(n_68), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_69), .B(n_230), .Y(n_556) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_70), .B(n_202), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_71), .A2(n_106), .B1(n_115), .B2(n_827), .Y(n_105) );
XOR2xp5_ASAP7_75t_L g130 ( .A(n_72), .B(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_73), .A2(n_104), .B1(n_135), .B2(n_136), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_73), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_74), .A2(n_166), .B(n_291), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_75), .A2(n_815), .B1(n_816), .B2(n_818), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_75), .Y(n_815) );
INVx1_ASAP7_75t_L g164 ( .A(n_76), .Y(n_164) );
INVx1_ASAP7_75t_L g180 ( .A(n_76), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_77), .B(n_156), .Y(n_246) );
AND2x2_ASAP7_75t_L g183 ( .A(n_79), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g222 ( .A(n_80), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_81), .A2(n_166), .B(n_172), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_82), .A2(n_166), .B(n_197), .C(n_201), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_83), .A2(n_88), .B1(n_156), .B2(n_533), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_84), .B(n_533), .Y(n_570) );
INVx1_ASAP7_75t_L g110 ( .A(n_86), .Y(n_110) );
AND2x2_ASAP7_75t_SL g205 ( .A(n_87), .B(n_184), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_89), .A2(n_166), .B1(n_241), .B2(n_242), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_90), .B(n_227), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_91), .B(n_227), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_92), .A2(n_521), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g209 ( .A(n_94), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_95), .B(n_230), .Y(n_568) );
AND2x2_ASAP7_75t_L g247 ( .A(n_96), .B(n_184), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_97), .A2(n_260), .B(n_261), .C(n_263), .Y(n_259) );
INVxp67_ASAP7_75t_L g520 ( .A(n_98), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_99), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_100), .B(n_230), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_101), .A2(n_521), .B(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g120 ( .A(n_102), .Y(n_120) );
INVx1_ASAP7_75t_SL g802 ( .A(n_102), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_103), .B(n_176), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_104), .Y(n_136) );
INVx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g828 ( .A(n_107), .Y(n_828) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_111), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_110), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g124 ( .A(n_114), .B(n_125), .Y(n_124) );
AND2x6_ASAP7_75t_SL g505 ( .A(n_114), .B(n_125), .Y(n_505) );
OR2x6_ASAP7_75t_SL g796 ( .A(n_114), .B(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_114), .B(n_797), .Y(n_823) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_800), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_128), .Y(n_121) );
INVx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g797 ( .A(n_125), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B1(n_137), .B2(n_798), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_504), .B1(n_506), .B2(n_794), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_139), .A2(n_504), .B1(n_507), .B2(n_799), .Y(n_798) );
AND3x1_ASAP7_75t_L g139 ( .A(n_140), .B(n_498), .C(n_501), .Y(n_139) );
NAND5xp2_ASAP7_75t_L g140 ( .A(n_141), .B(n_398), .C(n_428), .D(n_442), .E(n_468), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI21xp33_ASAP7_75t_L g498 ( .A1(n_142), .A2(n_441), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g811 ( .A(n_142), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_347), .Y(n_142) );
NOR3xp33_ASAP7_75t_SL g143 ( .A(n_144), .B(n_295), .C(n_329), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_212), .B(n_234), .C(n_273), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_187), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_147), .B(n_285), .Y(n_350) );
AND2x2_ASAP7_75t_L g437 ( .A(n_147), .B(n_215), .Y(n_437) );
HB1xp67_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OR2x2_ASAP7_75t_L g233 ( .A(n_148), .B(n_204), .Y(n_233) );
INVx1_ASAP7_75t_L g275 ( .A(n_148), .Y(n_275) );
INVx2_ASAP7_75t_L g280 ( .A(n_148), .Y(n_280) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_148), .Y(n_308) );
INVx1_ASAP7_75t_L g322 ( .A(n_148), .Y(n_322) );
AND2x2_ASAP7_75t_L g326 ( .A(n_148), .B(n_217), .Y(n_326) );
AND2x2_ASAP7_75t_L g407 ( .A(n_148), .B(n_216), .Y(n_407) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_154), .B(n_183), .Y(n_148) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_149), .A2(n_538), .B(n_544), .Y(n_537) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_149), .A2(n_565), .B(n_571), .Y(n_564) );
AO21x2_ASAP7_75t_L g602 ( .A1(n_149), .A2(n_538), .B(n_544), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_150), .Y(n_149) );
OA21x2_ASAP7_75t_L g594 ( .A1(n_150), .A2(n_595), .B(n_599), .Y(n_594) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x4_ASAP7_75t_L g195 ( .A(n_152), .B(n_153), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_165), .Y(n_154) );
INVx1_ASAP7_75t_L g272 ( .A(n_156), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_156), .A2(n_166), .B1(n_514), .B2(n_516), .Y(n_513) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_162), .Y(n_156) );
INVx1_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_160), .Y(n_157) );
OR2x6_ASAP7_75t_L g174 ( .A(n_158), .B(n_170), .Y(n_174) );
INVxp33_ASAP7_75t_L g244 ( .A(n_158), .Y(n_244) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g171 ( .A(n_159), .B(n_161), .Y(n_171) );
AND2x4_ASAP7_75t_L g230 ( .A(n_159), .B(n_179), .Y(n_230) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
BUFx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x6_ASAP7_75t_L g521 ( .A(n_163), .B(n_171), .Y(n_521) );
INVx2_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
AND2x6_ASAP7_75t_L g227 ( .A(n_164), .B(n_177), .Y(n_227) );
INVxp67_ASAP7_75t_L g270 ( .A(n_166), .Y(n_270) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_171), .Y(n_166) );
NOR2x1p5_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
INVx1_ASAP7_75t_L g245 ( .A(n_169), .Y(n_245) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_181), .Y(n_172) );
INVx2_ASAP7_75t_L g200 ( .A(n_174), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_174), .A2(n_181), .B(n_209), .C(n_210), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_174), .A2(n_221), .B1(n_222), .B2(n_223), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_SL g251 ( .A1(n_174), .A2(n_181), .B(n_252), .C(n_253), .Y(n_251) );
INVxp67_ASAP7_75t_L g260 ( .A(n_174), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_174), .A2(n_181), .B(n_292), .C(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
AND2x4_ASAP7_75t_L g533 ( .A(n_176), .B(n_182), .Y(n_533) );
AND2x4_ASAP7_75t_L g176 ( .A(n_177), .B(n_179), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_181), .A2(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_181), .B(n_195), .Y(n_231) );
INVx1_ASAP7_75t_L g241 ( .A(n_181), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_181), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_181), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_181), .A2(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_181), .A2(n_568), .B(n_569), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_181), .A2(n_589), .B(n_590), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_181), .A2(n_597), .B(n_598), .Y(n_596) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_182), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_184), .A2(n_259), .B1(n_264), .B2(n_265), .Y(n_258) );
INVx3_ASAP7_75t_L g265 ( .A(n_184), .Y(n_265) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_185), .B(n_268), .Y(n_267) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_185), .A2(n_527), .B(n_534), .Y(n_526) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx4f_ASAP7_75t_L g202 ( .A(n_186), .Y(n_202) );
AND2x4_ASAP7_75t_SL g187 ( .A(n_188), .B(n_203), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
AND2x2_ASAP7_75t_L g276 ( .A(n_189), .B(n_217), .Y(n_276) );
AND2x2_ASAP7_75t_L g297 ( .A(n_189), .B(n_204), .Y(n_297) );
INVx1_ASAP7_75t_L g320 ( .A(n_189), .Y(n_320) );
AND2x4_ASAP7_75t_L g387 ( .A(n_189), .B(n_216), .Y(n_387) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_196), .Y(n_189) );
NOR3xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .C(n_194), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_195), .A2(n_207), .B(n_211), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_195), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_195), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_195), .B(n_520), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_195), .B(n_223), .C(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_195), .A2(n_552), .B(n_553), .Y(n_551) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_201), .A2(n_239), .B(n_247), .Y(n_238) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_201), .A2(n_239), .B(n_247), .Y(n_302) );
AOI21x1_ASAP7_75t_L g559 ( .A1(n_201), .A2(n_560), .B(n_563), .Y(n_559) );
INVx2_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_202), .A2(n_250), .B(n_254), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_202), .A2(n_586), .B(n_587), .Y(n_585) );
AND2x4_ASAP7_75t_L g403 ( .A(n_203), .B(n_320), .Y(n_403) );
OR2x2_ASAP7_75t_L g444 ( .A(n_203), .B(n_445), .Y(n_444) );
NOR2xp67_ASAP7_75t_SL g463 ( .A(n_203), .B(n_336), .Y(n_463) );
NOR2x1_ASAP7_75t_L g481 ( .A(n_203), .B(n_395), .Y(n_481) );
INVx4_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2x1_ASAP7_75t_SL g281 ( .A(n_204), .B(n_217), .Y(n_281) );
AND2x4_ASAP7_75t_L g319 ( .A(n_204), .B(n_320), .Y(n_319) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_204), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_204), .B(n_279), .Y(n_357) );
INVx2_ASAP7_75t_L g371 ( .A(n_204), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_204), .B(n_323), .Y(n_393) );
AND2x2_ASAP7_75t_L g485 ( .A(n_204), .B(n_343), .Y(n_485) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2x1_ASAP7_75t_L g213 ( .A(n_214), .B(n_233), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_215), .B(n_322), .Y(n_336) );
AND2x2_ASAP7_75t_SL g345 ( .A(n_215), .B(n_325), .Y(n_345) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_232), .Y(n_215) );
INVx1_ASAP7_75t_L g323 ( .A(n_216), .Y(n_323) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g343 ( .A(n_217), .Y(n_343) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_224), .B(n_231), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_223), .B(n_262), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B1(n_228), .B2(n_229), .Y(n_224) );
INVxp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVxp67_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g376 ( .A(n_232), .Y(n_376) );
INVx2_ASAP7_75t_SL g421 ( .A(n_233), .Y(n_421) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_255), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_236), .B(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g367 ( .A(n_236), .Y(n_367) );
AND2x2_ASAP7_75t_L g491 ( .A(n_236), .B(n_316), .Y(n_491) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_248), .Y(n_236) );
AND2x4_ASAP7_75t_L g304 ( .A(n_237), .B(n_286), .Y(n_304) );
INVx1_ASAP7_75t_L g315 ( .A(n_237), .Y(n_315) );
AND2x2_ASAP7_75t_L g346 ( .A(n_237), .B(n_301), .Y(n_346) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_238), .B(n_249), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_238), .B(n_287), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_240), .B(n_246), .Y(n_239) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g284 ( .A(n_249), .Y(n_284) );
AND2x4_ASAP7_75t_L g352 ( .A(n_249), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g364 ( .A(n_249), .Y(n_364) );
INVx1_ASAP7_75t_L g406 ( .A(n_249), .Y(n_406) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_249), .Y(n_418) );
AND2x2_ASAP7_75t_L g434 ( .A(n_249), .B(n_257), .Y(n_434) );
BUFx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g381 ( .A(n_256), .B(n_339), .Y(n_381) );
INVx1_ASAP7_75t_SL g383 ( .A(n_256), .Y(n_383) );
AND2x2_ASAP7_75t_L g404 ( .A(n_256), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x4_ASAP7_75t_L g283 ( .A(n_257), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g311 ( .A(n_257), .Y(n_311) );
INVx2_ASAP7_75t_L g317 ( .A(n_257), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_257), .B(n_287), .Y(n_332) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_266), .Y(n_257) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_265), .A2(n_288), .B(n_294), .Y(n_287) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_265), .A2(n_288), .B(n_294), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B1(n_271), .B2(n_272), .Y(n_266) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B(n_282), .Y(n_273) );
INVx1_ASAP7_75t_L g413 ( .A(n_274), .Y(n_413) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g333 ( .A(n_276), .Y(n_333) );
AND2x2_ASAP7_75t_L g389 ( .A(n_276), .B(n_325), .Y(n_389) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx1_ASAP7_75t_L g303 ( .A(n_278), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_278), .B(n_319), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_278), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g410 ( .A(n_278), .B(n_403), .Y(n_410) );
AND2x2_ASAP7_75t_L g484 ( .A(n_278), .B(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_279), .Y(n_472) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_280), .Y(n_392) );
AND2x2_ASAP7_75t_L g305 ( .A(n_281), .B(n_306), .Y(n_305) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_281), .A2(n_494), .B(n_496), .Y(n_493) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx3_ASAP7_75t_L g379 ( .A(n_283), .Y(n_379) );
NAND2x1_ASAP7_75t_SL g423 ( .A(n_283), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g426 ( .A(n_283), .B(n_304), .Y(n_426) );
AND2x2_ASAP7_75t_L g338 ( .A(n_285), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g475 ( .A(n_285), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g486 ( .A(n_285), .B(n_434), .Y(n_486) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_286), .B(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g417 ( .A(n_287), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
OAI21xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_309), .B(n_312), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_304), .B2(n_305), .Y(n_296) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_297), .Y(n_354) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .Y(n_298) );
AND2x2_ASAP7_75t_L g327 ( .A(n_299), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g433 ( .A(n_299), .B(n_434), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_299), .A2(n_452), .B1(n_453), .B2(n_454), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_299), .B(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g316 ( .A(n_301), .B(n_317), .Y(n_316) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_301), .B(n_317), .Y(n_397) );
NOR2x1_ASAP7_75t_L g405 ( .A(n_301), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g353 ( .A(n_302), .Y(n_353) );
AND2x2_ASAP7_75t_L g361 ( .A(n_302), .B(n_317), .Y(n_361) );
INVx1_ASAP7_75t_L g424 ( .A(n_302), .Y(n_424) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2x1_ASAP7_75t_L g342 ( .A(n_307), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g454 ( .A(n_310), .B(n_339), .Y(n_454) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g328 ( .A(n_311), .Y(n_328) );
AND2x2_ASAP7_75t_L g351 ( .A(n_311), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g439 ( .A(n_311), .B(n_346), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_318), .B1(n_324), .B2(n_327), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g447 ( .A(n_314), .B(n_448), .Y(n_447) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g477 ( .A(n_317), .B(n_364), .Y(n_477) );
AND2x2_ASAP7_75t_SL g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx2_ASAP7_75t_L g344 ( .A(n_319), .Y(n_344) );
OAI21xp33_ASAP7_75t_SL g490 ( .A1(n_319), .A2(n_491), .B(n_492), .Y(n_490) );
AND2x4_ASAP7_75t_SL g321 ( .A(n_322), .B(n_323), .Y(n_321) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_322), .Y(n_480) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
O2A1O1Ixp33_ASAP7_75t_SL g422 ( .A1(n_325), .A2(n_423), .B(n_425), .C(n_427), .Y(n_422) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_326), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g427 ( .A(n_326), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_326), .B(n_403), .Y(n_467) );
INVx1_ASAP7_75t_SL g334 ( .A(n_327), .Y(n_334) );
AND2x2_ASAP7_75t_L g415 ( .A(n_328), .B(n_352), .Y(n_415) );
INVx1_ASAP7_75t_L g460 ( .A(n_328), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B1(n_334), .B2(n_335), .C(n_337), .Y(n_329) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_330), .Y(n_449) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g497 ( .A(n_332), .B(n_340), .Y(n_497) );
OR2x2_ASAP7_75t_L g356 ( .A(n_333), .B(n_357), .Y(n_356) );
NOR2x1_ASAP7_75t_L g369 ( .A(n_333), .B(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_333), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g495 ( .A(n_333), .B(n_392), .Y(n_495) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI32xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .A3(n_344), .B1(n_345), .B2(n_346), .Y(n_337) );
INVx1_ASAP7_75t_L g358 ( .A(n_339), .Y(n_358) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_341), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g453 ( .A(n_342), .Y(n_453) );
OAI22xp33_ASAP7_75t_SL g435 ( .A1(n_344), .A2(n_436), .B1(n_438), .B2(n_440), .Y(n_435) );
INVx1_ASAP7_75t_L g466 ( .A(n_345), .Y(n_466) );
AOI211x1_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_354), .B(n_355), .C(n_372), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_349), .B(n_434), .Y(n_440) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g396 ( .A(n_352), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g462 ( .A(n_352), .Y(n_462) );
OAI222xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B1(n_359), .B2(n_365), .C1(n_366), .C2(n_368), .Y(n_355) );
INVxp67_ASAP7_75t_L g452 ( .A(n_356), .Y(n_452) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_360), .B(n_445), .Y(n_492) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g408 ( .A(n_361), .B(n_405), .Y(n_408) );
INVx3_ASAP7_75t_L g448 ( .A(n_363), .Y(n_448) );
BUFx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g386 ( .A(n_371), .B(n_387), .Y(n_386) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_377), .B1(n_380), .B2(n_385), .C(n_388), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_374), .A2(n_431), .B(n_433), .Y(n_430) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g384 ( .A(n_378), .Y(n_384) );
OR2x2_ASAP7_75t_L g488 ( .A(n_379), .B(n_424), .Y(n_488) );
NOR2xp67_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_382), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_385), .A2(n_414), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_386), .A2(n_458), .B(n_465), .Y(n_464) );
INVx4_ASAP7_75t_L g395 ( .A(n_387), .Y(n_395) );
OAI31xp33_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_390), .A3(n_394), .B(n_396), .Y(n_388) );
INVx1_ASAP7_75t_L g446 ( .A(n_390), .Y(n_446) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_411), .Y(n_398) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_399), .B(n_411), .C(n_430), .D(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_409), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_404), .B1(n_407), .B2(n_408), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g471 ( .A(n_403), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_404), .B(n_424), .Y(n_432) );
INVx1_ASAP7_75t_SL g445 ( .A(n_407), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_422), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_416), .B2(n_419), .Y(n_412) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2x1_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_421), .A2(n_484), .B1(n_486), .B2(n_487), .Y(n_483) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_435), .C(n_441), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g500 ( .A(n_435), .Y(n_500) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI21xp33_ASAP7_75t_L g501 ( .A1(n_441), .A2(n_502), .B(n_503), .Y(n_501) );
INVxp33_ASAP7_75t_L g502 ( .A(n_442), .Y(n_502) );
AND2x2_ASAP7_75t_L g810 ( .A(n_442), .B(n_468), .Y(n_810) );
NOR2xp67_ASAP7_75t_L g442 ( .A(n_443), .B(n_450), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .B1(n_447), .B2(n_449), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_447), .A2(n_470), .B(n_473), .Y(n_469) );
INVx2_ASAP7_75t_L g457 ( .A(n_448), .Y(n_457) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_455), .C(n_464), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_458), .B1(n_461), .B2(n_463), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVxp33_ASAP7_75t_SL g503 ( .A(n_468), .Y(n_503) );
NOR3x1_ASAP7_75t_L g468 ( .A(n_469), .B(n_482), .C(n_489), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_490), .B(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g812 ( .A(n_499), .Y(n_812) );
CKINVDCx11_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_671), .Y(n_507) );
NOR4xp25_ASAP7_75t_L g508 ( .A(n_509), .B(n_614), .C(n_653), .D(n_660), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_535), .B1(n_572), .B2(n_581), .C(n_600), .Y(n_509) );
OR2x2_ASAP7_75t_L g744 ( .A(n_510), .B(n_606), .Y(n_744) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g659 ( .A(n_511), .B(n_584), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_511), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_SL g724 ( .A(n_511), .B(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_524), .Y(n_511) );
AND2x4_ASAP7_75t_SL g583 ( .A(n_512), .B(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g605 ( .A(n_512), .Y(n_605) );
AND2x2_ASAP7_75t_L g640 ( .A(n_512), .B(n_613), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_512), .B(n_525), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_512), .B(n_607), .Y(n_692) );
OR2x2_ASAP7_75t_L g770 ( .A(n_512), .B(n_584), .Y(n_770) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_518), .Y(n_512) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g592 ( .A(n_525), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_525), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g618 ( .A(n_525), .Y(n_618) );
OR2x2_ASAP7_75t_L g623 ( .A(n_525), .B(n_607), .Y(n_623) );
AND2x2_ASAP7_75t_L g636 ( .A(n_525), .B(n_594), .Y(n_636) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_525), .Y(n_639) );
INVx1_ASAP7_75t_L g651 ( .A(n_525), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_525), .B(n_605), .Y(n_716) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_532), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_536), .B(n_545), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g580 ( .A(n_537), .B(n_564), .Y(n_580) );
AND2x4_ASAP7_75t_L g610 ( .A(n_537), .B(n_549), .Y(n_610) );
INVx2_ASAP7_75t_L g644 ( .A(n_537), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_537), .B(n_564), .Y(n_702) );
AND2x2_ASAP7_75t_L g749 ( .A(n_537), .B(n_578), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
AOI222xp33_ASAP7_75t_L g737 ( .A1(n_545), .A2(n_609), .B1(n_652), .B2(n_712), .C1(n_738), .C2(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_557), .Y(n_546) );
AND2x2_ASAP7_75t_L g656 ( .A(n_547), .B(n_576), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_547), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g785 ( .A(n_547), .B(n_625), .Y(n_785) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_548), .A2(n_616), .B(n_620), .Y(n_615) );
AND2x2_ASAP7_75t_L g696 ( .A(n_548), .B(n_579), .Y(n_696) );
OR2x2_ASAP7_75t_L g721 ( .A(n_548), .B(n_580), .Y(n_721) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx5_ASAP7_75t_L g575 ( .A(n_549), .Y(n_575) );
AND2x2_ASAP7_75t_L g662 ( .A(n_549), .B(n_644), .Y(n_662) );
AND2x2_ASAP7_75t_L g688 ( .A(n_549), .B(n_564), .Y(n_688) );
OR2x2_ASAP7_75t_L g691 ( .A(n_549), .B(n_578), .Y(n_691) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_549), .Y(n_709) );
AND2x4_ASAP7_75t_SL g766 ( .A(n_549), .B(n_643), .Y(n_766) );
OR2x2_ASAP7_75t_L g775 ( .A(n_549), .B(n_602), .Y(n_775) );
OR2x6_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g608 ( .A(n_557), .Y(n_608) );
AOI221xp5_ASAP7_75t_SL g726 ( .A1(n_557), .A2(n_610), .B1(n_727), .B2(n_729), .C(n_730), .Y(n_726) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_564), .Y(n_557) );
OR2x2_ASAP7_75t_L g665 ( .A(n_558), .B(n_635), .Y(n_665) );
OR2x2_ASAP7_75t_L g675 ( .A(n_558), .B(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g701 ( .A(n_558), .B(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g707 ( .A(n_558), .B(n_626), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_558), .B(n_690), .Y(n_719) );
INVx2_ASAP7_75t_L g732 ( .A(n_558), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g753 ( .A(n_558), .B(n_610), .Y(n_753) );
AND2x2_ASAP7_75t_L g757 ( .A(n_558), .B(n_579), .Y(n_757) );
AND2x2_ASAP7_75t_L g765 ( .A(n_558), .B(n_766), .Y(n_765) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g578 ( .A(n_559), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_564), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g609 ( .A(n_564), .B(n_578), .Y(n_609) );
INVx2_ASAP7_75t_L g626 ( .A(n_564), .Y(n_626) );
AND2x4_ASAP7_75t_L g643 ( .A(n_564), .B(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_564), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g755 ( .A(n_574), .B(n_577), .Y(n_755) );
AND2x4_ASAP7_75t_L g601 ( .A(n_575), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g642 ( .A(n_575), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g669 ( .A(n_575), .B(n_609), .Y(n_669) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
AND2x2_ASAP7_75t_L g773 ( .A(n_577), .B(n_774), .Y(n_773) );
BUFx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g625 ( .A(n_578), .B(n_626), .Y(n_625) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_579), .A2(n_646), .B(n_652), .Y(n_645) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_592), .Y(n_582) );
INVx1_ASAP7_75t_SL g699 ( .A(n_583), .Y(n_699) );
AND2x2_ASAP7_75t_L g729 ( .A(n_583), .B(n_639), .Y(n_729) );
AND2x4_ASAP7_75t_L g740 ( .A(n_583), .B(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g606 ( .A(n_584), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g613 ( .A(n_584), .Y(n_613) );
AND2x4_ASAP7_75t_L g619 ( .A(n_584), .B(n_605), .Y(n_619) );
INVx2_ASAP7_75t_L g630 ( .A(n_584), .Y(n_630) );
INVx1_ASAP7_75t_L g679 ( .A(n_584), .Y(n_679) );
OR2x2_ASAP7_75t_L g700 ( .A(n_584), .B(n_684), .Y(n_700) );
OR2x2_ASAP7_75t_L g714 ( .A(n_584), .B(n_594), .Y(n_714) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_584), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_584), .B(n_636), .Y(n_786) );
OR2x6_ASAP7_75t_L g584 ( .A(n_585), .B(n_591), .Y(n_584) );
INVx1_ASAP7_75t_L g631 ( .A(n_592), .Y(n_631) );
AND2x2_ASAP7_75t_L g764 ( .A(n_592), .B(n_630), .Y(n_764) );
AND2x2_ASAP7_75t_L g789 ( .A(n_592), .B(n_619), .Y(n_789) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g607 ( .A(n_594), .Y(n_607) );
BUFx3_ASAP7_75t_L g649 ( .A(n_594), .Y(n_649) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_594), .Y(n_676) );
INVx1_ASAP7_75t_L g685 ( .A(n_594), .Y(n_685) );
AOI33xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_603), .A3(n_608), .B1(n_609), .B2(n_610), .B3(n_611), .Y(n_600) );
AOI21x1_ASAP7_75t_SL g703 ( .A1(n_601), .A2(n_625), .B(n_687), .Y(n_703) );
INVx2_ASAP7_75t_L g733 ( .A(n_601), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_601), .B(n_732), .Y(n_739) );
AND2x2_ASAP7_75t_L g687 ( .A(n_602), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AND2x2_ASAP7_75t_L g650 ( .A(n_605), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g751 ( .A(n_606), .Y(n_751) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_607), .Y(n_741) );
OAI32xp33_ASAP7_75t_L g790 ( .A1(n_608), .A2(n_610), .A3(n_786), .B1(n_791), .B2(n_793), .Y(n_790) );
AND2x2_ASAP7_75t_L g708 ( .A(n_609), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_SL g698 ( .A(n_610), .Y(n_698) );
AND2x2_ASAP7_75t_L g763 ( .A(n_610), .B(n_707), .Y(n_763) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_624), .B1(n_627), .B2(n_641), .C(n_645), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_618), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_619), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_619), .B(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_619), .B(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g668 ( .A(n_623), .Y(n_668) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_632), .C(n_637), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_629), .A2(n_691), .B1(n_731), .B2(n_734), .Y(n_730) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g634 ( .A(n_630), .Y(n_634) );
NOR2x1p5_ASAP7_75t_L g648 ( .A(n_630), .B(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_630), .Y(n_670) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI322xp33_ASAP7_75t_L g697 ( .A1(n_633), .A2(n_675), .A3(n_698), .B1(n_699), .B2(n_700), .C1(n_701), .C2(n_703), .Y(n_697) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g653 ( .A1(n_635), .A2(n_654), .B(n_655), .C(n_657), .Y(n_653) );
OR2x2_ASAP7_75t_L g745 ( .A(n_635), .B(n_699), .Y(n_745) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g652 ( .A(n_636), .B(n_640), .Y(n_652) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g658 ( .A(n_642), .B(n_659), .Y(n_658) );
INVx3_ASAP7_75t_SL g690 ( .A(n_643), .Y(n_690) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_647), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_SL g694 ( .A(n_650), .Y(n_694) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_651), .Y(n_736) );
OR2x6_ASAP7_75t_SL g791 ( .A(n_654), .B(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g781 ( .A1(n_659), .A2(n_782), .B(n_783), .C(n_790), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_663), .B(n_666), .C(n_670), .Y(n_660) );
OAI211xp5_ASAP7_75t_SL g672 ( .A1(n_661), .A2(n_673), .B(n_680), .C(n_704), .Y(n_672) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_717), .C(n_761), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_676), .Y(n_768) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g723 ( .A(n_679), .Y(n_723) );
NOR3xp33_ASAP7_75t_SL g680 ( .A(n_681), .B(n_693), .C(n_697), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_686), .B1(n_689), .B2(n_692), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g725 ( .A(n_685), .Y(n_725) );
INVxp67_ASAP7_75t_SL g792 ( .A(n_685), .Y(n_792) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_SL g778 ( .A(n_691), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
OR2x2_ASAP7_75t_L g728 ( .A(n_694), .B(n_714), .Y(n_728) );
OR2x2_ASAP7_75t_L g779 ( .A(n_694), .B(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g777 ( .A(n_702), .Y(n_777) );
OR2x2_ASAP7_75t_L g793 ( .A(n_702), .B(n_732), .Y(n_793) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B(n_710), .Y(n_704) );
OAI31xp33_ASAP7_75t_L g718 ( .A1(n_705), .A2(n_719), .A3(n_720), .B(n_722), .Y(n_718) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
AND2x4_ASAP7_75t_L g750 ( .A(n_715), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND4xp25_ASAP7_75t_SL g717 ( .A(n_718), .B(n_726), .C(n_737), .D(n_742), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_725), .Y(n_760) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_746), .B1(n_750), .B2(n_752), .C(n_754), .Y(n_742) );
NAND2xp33_ASAP7_75t_SL g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g787 ( .A(n_746), .Y(n_787) );
AND2x2_ASAP7_75t_SL g746 ( .A(n_747), .B(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g782 ( .A(n_756), .Y(n_782) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_762), .B(n_781), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B1(n_765), .B2(n_767), .C(n_771), .Y(n_762) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
AOI21xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_776), .B(n_779), .Y(n_771) );
INVxp33_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_786), .B1(n_787), .B2(n_788), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_795), .Y(n_799) );
CKINVDCx11_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_803), .B(n_824), .Y(n_800) );
INVx2_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B(n_819), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_804), .A2(n_820), .B(n_821), .Y(n_819) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g820 ( .A(n_808), .Y(n_820) );
XNOR2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_813), .Y(n_808) );
NAND3x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .C(n_812), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g818 ( .A(n_816), .Y(n_818) );
CKINVDCx11_ASAP7_75t_R g826 ( .A(n_821), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
BUFx3_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_SL g827 ( .A(n_828), .Y(n_827) );
endmodule