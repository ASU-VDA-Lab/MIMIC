module fake_netlist_5_726_n_1380 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1380);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1380;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_370;
wire n_976;
wire n_343;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1377;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_1332;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_132),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_216),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_3),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_332),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_98),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_42),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_213),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_184),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_290),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_62),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_259),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_65),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_75),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_272),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_53),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_90),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_93),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_77),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_193),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_115),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_138),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_145),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_335),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_162),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_313),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_30),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_331),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_30),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_28),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_17),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_186),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_276),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_51),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_245),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_163),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_43),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_142),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_87),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_268),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_223),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_278),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_69),
.Y(n_381)
);

BUFx10_ASAP7_75t_L g382 ( 
.A(n_18),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_126),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_74),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_28),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_229),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_92),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_249),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_173),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_89),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_182),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_224),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_205),
.Y(n_393)
);

BUFx10_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_73),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_219),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_82),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_305),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_106),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_295),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_102),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_104),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_252),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_256),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_66),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_155),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_273),
.Y(n_408)
);

BUFx10_ASAP7_75t_L g409 ( 
.A(n_50),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_156),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_140),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_26),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_19),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_169),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_279),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_127),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_210),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_22),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_171),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_53),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_207),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_120),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_303),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_329),
.Y(n_424)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_188),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_137),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_3),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_315),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_21),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_55),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_262),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_58),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_266),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_24),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_14),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_64),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_22),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_267),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_228),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_217),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_280),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_203),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_327),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_101),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_284),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_122),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_144),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_76),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_158),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_55),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_79),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_176),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_13),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_47),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_7),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_97),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_67),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_239),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_238),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_174),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_32),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_129),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_153),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_78),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_200),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_227),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_326),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_215),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_71),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_11),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_299),
.Y(n_471)
);

BUFx2_ASAP7_75t_SL g472 ( 
.A(n_248),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_237),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_51),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_25),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_37),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_177),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_59),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_110),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_152),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_328),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_119),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_160),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_17),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_139),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_149),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_24),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_288),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_34),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_226),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_121),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_95),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_125),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_165),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_312),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_35),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_170),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_88),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_19),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_180),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_192),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_307),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_94),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_281),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_232),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_33),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_118),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_181),
.Y(n_508)
);

BUFx5_ASAP7_75t_L g509 ( 
.A(n_146),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_179),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_52),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_195),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_128),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_214),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_21),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_117),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_135),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_269),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_330),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_401),
.B(n_0),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_386),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_365),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_366),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_382),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_391),
.B(n_0),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_386),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_401),
.B(n_1),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_342),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_365),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_487),
.Y(n_530)
);

CKINVDCx11_ASAP7_75t_R g531 ( 
.A(n_382),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_487),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_486),
.B(n_1),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_386),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_386),
.Y(n_535)
);

BUFx8_ASAP7_75t_SL g536 ( 
.A(n_364),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_406),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_487),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_406),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_406),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_487),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_486),
.B(n_2),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_418),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_2),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_501),
.B(n_4),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_406),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_454),
.B(n_4),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_407),
.B(n_448),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_444),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_336),
.Y(n_550)
);

BUFx8_ASAP7_75t_SL g551 ( 
.A(n_430),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_418),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_418),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_515),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_515),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_393),
.B(n_5),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_444),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_431),
.B(n_5),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_355),
.B(n_6),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_384),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_503),
.B(n_6),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_355),
.B(n_7),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_444),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_346),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_515),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_369),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_346),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_447),
.B(n_8),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_350),
.B(n_8),
.Y(n_570)
);

BUFx12f_ASAP7_75t_L g571 ( 
.A(n_409),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_509),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_372),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_414),
.B(n_9),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_414),
.B(n_9),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_368),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_412),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_366),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_358),
.B(n_10),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_377),
.B(n_383),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_392),
.B(n_10),
.Y(n_581)
);

BUFx8_ASAP7_75t_SL g582 ( 
.A(n_437),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_346),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_425),
.B(n_11),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_380),
.B(n_12),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_507),
.B(n_12),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_420),
.B(n_13),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_387),
.B(n_400),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_470),
.B(n_14),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_475),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_357),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_476),
.B(n_15),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_499),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_341),
.B(n_15),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_349),
.B(n_16),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_511),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_384),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_409),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_351),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_357),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_337),
.Y(n_604)
);

CKINVDCx6p67_ASAP7_75t_R g605 ( 
.A(n_434),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_353),
.B(n_354),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_356),
.B(n_16),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_360),
.B(n_18),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_394),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_357),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_367),
.B(n_20),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_370),
.B(n_63),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_376),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_340),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_394),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_509),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_509),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_379),
.B(n_20),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_388),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_530),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_543),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_520),
.A2(n_427),
.B1(n_352),
.B2(n_375),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_520),
.A2(n_496),
.B1(n_385),
.B2(n_413),
.Y(n_623)
);

OA22x2_ASAP7_75t_L g624 ( 
.A1(n_523),
.A2(n_429),
.B1(n_432),
.B2(n_338),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_576),
.Y(n_625)
);

OAI22xp33_ASAP7_75t_L g626 ( 
.A1(n_527),
.A2(n_453),
.B1(n_474),
.B2(n_450),
.Y(n_626)
);

AO22x2_ASAP7_75t_L g627 ( 
.A1(n_542),
.A2(n_472),
.B1(n_390),
.B2(n_402),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_588),
.B(n_528),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_604),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_SL g630 ( 
.A1(n_527),
.A2(n_544),
.B1(n_548),
.B2(n_575),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_579),
.A2(n_362),
.B1(n_458),
.B2(n_363),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_584),
.A2(n_374),
.B1(n_404),
.B2(n_339),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_532),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_533),
.A2(n_545),
.B1(n_585),
.B2(n_544),
.Y(n_634)
);

OR2x6_ASAP7_75t_L g635 ( 
.A(n_524),
.B(n_399),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_560),
.A2(n_446),
.B1(n_469),
.B2(n_411),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_614),
.B(n_421),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_L g638 ( 
.A1(n_599),
.A2(n_484),
.B1(n_489),
.B2(n_478),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_563),
.A2(n_504),
.B1(n_483),
.B2(n_506),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_550),
.A2(n_419),
.B1(n_433),
.B2(n_405),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_614),
.B(n_421),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_522),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_L g643 ( 
.A1(n_599),
.A2(n_438),
.B1(n_439),
.B2(n_436),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g644 ( 
.A1(n_575),
.A2(n_449),
.B1(n_456),
.B2(n_440),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_538),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_529),
.B(n_435),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_568),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_536),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_568),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_541),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_523),
.B(n_23),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_574),
.A2(n_605),
.B1(n_571),
.B2(n_607),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_561),
.B(n_435),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_562),
.A2(n_578),
.B1(n_548),
.B2(n_581),
.Y(n_654)
);

AO22x2_ASAP7_75t_L g655 ( 
.A1(n_525),
.A2(n_457),
.B1(n_471),
.B2(n_463),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_553),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_555),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_618),
.A2(n_556),
.B1(n_559),
.B2(n_525),
.Y(n_658)
);

NAND3x1_ASAP7_75t_L g659 ( 
.A(n_562),
.B(n_481),
.C(n_477),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_556),
.A2(n_344),
.B1(n_345),
.B2(n_343),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_568),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_R g662 ( 
.A(n_531),
.B(n_347),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_578),
.A2(n_490),
.B1(n_500),
.B2(n_488),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_552),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_559),
.A2(n_359),
.B1(n_361),
.B2(n_348),
.Y(n_665)
);

OAI22xp5_ASAP7_75t_L g666 ( 
.A1(n_581),
.A2(n_373),
.B1(n_378),
.B2(n_371),
.Y(n_666)
);

AND2x2_ASAP7_75t_SL g667 ( 
.A(n_569),
.B(n_570),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_583),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_L g669 ( 
.A1(n_587),
.A2(n_510),
.B1(n_512),
.B2(n_502),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_598),
.B(n_23),
.Y(n_670)
);

AO22x2_ASAP7_75t_L g671 ( 
.A1(n_569),
.A2(n_516),
.B1(n_519),
.B2(n_514),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_L g672 ( 
.A1(n_587),
.A2(n_389),
.B1(n_395),
.B2(n_381),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_594),
.A2(n_397),
.B1(n_398),
.B2(n_396),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_609),
.B(n_455),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_615),
.B(n_455),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_L g676 ( 
.A1(n_589),
.A2(n_408),
.B1(n_410),
.B2(n_403),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_547),
.B(n_415),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_583),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_583),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_606),
.B(n_461),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_606),
.B(n_461),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_589),
.A2(n_417),
.B1(n_422),
.B2(n_416),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_591),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_594),
.A2(n_424),
.B1(n_426),
.B2(n_423),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_592),
.A2(n_441),
.B1(n_442),
.B2(n_428),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_570),
.B(n_68),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_592),
.A2(n_445),
.B1(n_451),
.B2(n_443),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_590),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_591),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_591),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_595),
.A2(n_608),
.B1(n_611),
.B2(n_586),
.Y(n_691)
);

AO22x2_ASAP7_75t_L g692 ( 
.A1(n_586),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_554),
.B(n_452),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_554),
.B(n_459),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_590),
.B(n_27),
.Y(n_695)
);

BUFx10_ASAP7_75t_L g696 ( 
.A(n_595),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_597),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_608),
.A2(n_485),
.B1(n_517),
.B2(n_513),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_566),
.B(n_460),
.Y(n_699)
);

AO22x2_ASAP7_75t_L g700 ( 
.A1(n_611),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_700)
);

OAI22xp33_ASAP7_75t_L g701 ( 
.A1(n_597),
.A2(n_518),
.B1(n_508),
.B2(n_505),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_521),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_580),
.B(n_462),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_702),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_683),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_661),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_683),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_678),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_628),
.B(n_566),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_648),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_647),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_679),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_690),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_668),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_689),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_633),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_645),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_630),
.A2(n_612),
.B(n_580),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_SL g719 ( 
.A(n_623),
.B(n_464),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_650),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_662),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_620),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_629),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_664),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_642),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_621),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_657),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_680),
.B(n_567),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_647),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_647),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_649),
.Y(n_731)
);

BUFx5_ASAP7_75t_L g732 ( 
.A(n_686),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_649),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_649),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_656),
.Y(n_735)
);

XOR2xp5_ASAP7_75t_L g736 ( 
.A(n_632),
.B(n_465),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_636),
.B(n_565),
.Y(n_737)
);

XOR2xp5_ASAP7_75t_L g738 ( 
.A(n_639),
.B(n_466),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_688),
.B(n_600),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_703),
.B(n_613),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_697),
.B(n_577),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_693),
.Y(n_742)
);

INVxp33_ASAP7_75t_L g743 ( 
.A(n_625),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_652),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_694),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_699),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_681),
.B(n_577),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_635),
.Y(n_748)
);

XNOR2xp5_ASAP7_75t_L g749 ( 
.A(n_640),
.B(n_551),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_634),
.B(n_619),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_696),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_696),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_654),
.B(n_619),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_646),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_667),
.Y(n_755)
);

XOR2x2_ASAP7_75t_L g756 ( 
.A(n_624),
.B(n_582),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_691),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_658),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_670),
.B(n_565),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_655),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_655),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_671),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_635),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_686),
.B(n_572),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_686),
.B(n_596),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_686),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_660),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_701),
.B(n_619),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_671),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_R g770 ( 
.A(n_653),
.B(n_467),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_677),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_677),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_674),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_R g774 ( 
.A(n_675),
.B(n_468),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_651),
.B(n_573),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_644),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_627),
.Y(n_777)
);

XNOR2x2_ASAP7_75t_L g778 ( 
.A(n_692),
.B(n_700),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_627),
.B(n_601),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_695),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_695),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_665),
.B(n_565),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_637),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_641),
.B(n_593),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_692),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_659),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_673),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_684),
.B(n_535),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_631),
.B(n_535),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_698),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_672),
.B(n_565),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_700),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_666),
.B(n_603),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_643),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_741),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_716),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_709),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_740),
.B(n_750),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_718),
.A2(n_682),
.B(n_676),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_740),
.B(n_750),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_771),
.B(n_612),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_718),
.A2(n_685),
.B(n_626),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_717),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_R g804 ( 
.A(n_710),
.B(n_473),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_742),
.B(n_612),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_755),
.B(n_687),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_721),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_758),
.B(n_638),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_766),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_747),
.B(n_745),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_786),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_722),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_746),
.B(n_612),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_739),
.B(n_753),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_783),
.B(n_622),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_705),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_753),
.B(n_602),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_766),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_728),
.B(n_616),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_728),
.B(n_617),
.Y(n_820)
);

BUFx12f_ASAP7_75t_SL g821 ( 
.A(n_789),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_707),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_720),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_743),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_724),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_757),
.B(n_521),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_784),
.B(n_521),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_766),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_732),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_726),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_764),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_788),
.B(n_669),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_727),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_711),
.Y(n_834)
);

HB1xp67_ASAP7_75t_L g835 ( 
.A(n_779),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_764),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_732),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_768),
.B(n_479),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_784),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_768),
.B(n_480),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_765),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_754),
.B(n_663),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_775),
.B(n_534),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_765),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_706),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_779),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_735),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_787),
.B(n_738),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_704),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_708),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_770),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_712),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_737),
.B(n_482),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_777),
.B(n_534),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_760),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_761),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_791),
.B(n_491),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_773),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_713),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_791),
.B(n_492),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_772),
.B(n_534),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_729),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_714),
.Y(n_863)
);

AND2x2_ASAP7_75t_SL g864 ( 
.A(n_785),
.B(n_537),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_730),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_794),
.B(n_537),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_715),
.Y(n_867)
);

AND2x2_ASAP7_75t_SL g868 ( 
.A(n_792),
.B(n_762),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_769),
.B(n_537),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_793),
.B(n_776),
.Y(n_870)
);

INVx3_ASAP7_75t_SL g871 ( 
.A(n_725),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_711),
.B(n_493),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_759),
.B(n_539),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_734),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_759),
.B(n_539),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_732),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_732),
.B(n_494),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_780),
.Y(n_878)
);

BUFx4f_ASAP7_75t_L g879 ( 
.A(n_782),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_732),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_782),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_751),
.B(n_539),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_731),
.B(n_733),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_752),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_781),
.B(n_540),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_778),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_723),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_814),
.B(n_736),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_867),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_816),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_807),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_814),
.B(n_767),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_818),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_839),
.B(n_790),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_887),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_839),
.B(n_744),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_818),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_816),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_855),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_798),
.B(n_495),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_867),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_822),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_822),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_887),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_800),
.B(n_497),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_797),
.B(n_748),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_818),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_824),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_824),
.B(n_719),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_817),
.B(n_498),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_797),
.B(n_763),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_828),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_887),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_795),
.B(n_749),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_795),
.B(n_29),
.Y(n_915)
);

OR2x6_ASAP7_75t_L g916 ( 
.A(n_881),
.B(n_756),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_796),
.Y(n_917)
);

CKINVDCx14_ASAP7_75t_R g918 ( 
.A(n_804),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_817),
.B(n_540),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_821),
.Y(n_920)
);

NOR2x1_ASAP7_75t_SL g921 ( 
.A(n_829),
.B(n_526),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_810),
.B(n_774),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_812),
.Y(n_923)
);

AND2x6_ASAP7_75t_L g924 ( 
.A(n_829),
.B(n_540),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_809),
.B(n_546),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_858),
.B(n_70),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_810),
.B(n_31),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_870),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_835),
.B(n_33),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_846),
.B(n_34),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_851),
.B(n_35),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_808),
.B(n_36),
.Y(n_932)
);

AND2x2_ASAP7_75t_SL g933 ( 
.A(n_879),
.B(n_546),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_812),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_828),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_809),
.B(n_828),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_881),
.B(n_546),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_871),
.Y(n_938)
);

BUFx4f_ASAP7_75t_L g939 ( 
.A(n_871),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_807),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_881),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_809),
.Y(n_942)
);

BUFx12f_ASAP7_75t_L g943 ( 
.A(n_858),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_796),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_871),
.B(n_36),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_830),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_832),
.B(n_37),
.Y(n_947)
);

AND2x6_ASAP7_75t_L g948 ( 
.A(n_829),
.B(n_549),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_884),
.B(n_72),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_809),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_803),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_830),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_803),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_836),
.B(n_549),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_843),
.B(n_870),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_884),
.B(n_80),
.Y(n_956)
);

BUFx12f_ASAP7_75t_L g957 ( 
.A(n_908),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_942),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_890),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_889),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_943),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_941),
.B(n_837),
.Y(n_962)
);

CKINVDCx8_ASAP7_75t_R g963 ( 
.A(n_891),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_954),
.A2(n_799),
.B(n_802),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_940),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_932),
.B(n_886),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_955),
.B(n_847),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_938),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_900),
.B(n_866),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_918),
.Y(n_970)
);

INVxp67_ASAP7_75t_SL g971 ( 
.A(n_942),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_895),
.Y(n_972)
);

INVxp67_ASAP7_75t_SL g973 ( 
.A(n_942),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_950),
.Y(n_974)
);

CKINVDCx8_ASAP7_75t_R g975 ( 
.A(n_920),
.Y(n_975)
);

NAND2x1p5_ASAP7_75t_L g976 ( 
.A(n_941),
.B(n_837),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_932),
.B(n_886),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_904),
.Y(n_978)
);

OR2x6_ASAP7_75t_L g979 ( 
.A(n_913),
.B(n_881),
.Y(n_979)
);

NAND2x1p5_ASAP7_75t_L g980 ( 
.A(n_941),
.B(n_950),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_950),
.Y(n_981)
);

BUFx2_ASAP7_75t_R g982 ( 
.A(n_909),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_897),
.Y(n_983)
);

INVx3_ASAP7_75t_SL g984 ( 
.A(n_896),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_897),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_901),
.B(n_847),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_893),
.B(n_837),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_917),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_939),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_899),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_898),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_903),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_897),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_900),
.B(n_866),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_899),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_907),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_922),
.B(n_831),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_928),
.Y(n_998)
);

INVx3_ASAP7_75t_SL g999 ( 
.A(n_896),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_907),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_939),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_907),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_936),
.Y(n_1003)
);

CKINVDCx11_ASAP7_75t_R g1004 ( 
.A(n_916),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_928),
.Y(n_1005)
);

BUFx4f_ASAP7_75t_SL g1006 ( 
.A(n_894),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_906),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_893),
.Y(n_1008)
);

BUFx2_ASAP7_75t_SL g1009 ( 
.A(n_906),
.Y(n_1009)
);

INVxp67_ASAP7_75t_SL g1010 ( 
.A(n_936),
.Y(n_1010)
);

CKINVDCx6p67_ASAP7_75t_R g1011 ( 
.A(n_916),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_894),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_915),
.A2(n_848),
.B(n_815),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_892),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_945),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_912),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_944),
.Y(n_1017)
);

INVx6_ASAP7_75t_L g1018 ( 
.A(n_957),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_957),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_966),
.A2(n_879),
.B1(n_840),
.B2(n_838),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_974),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_970),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_960),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_988),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_985),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_968),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_974),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1017),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_1013),
.A2(n_888),
.B1(n_802),
.B2(n_806),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_968),
.Y(n_1030)
);

BUFx8_ASAP7_75t_SL g1031 ( 
.A(n_970),
.Y(n_1031)
);

BUFx2_ASAP7_75t_SL g1032 ( 
.A(n_963),
.Y(n_1032)
);

OAI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_966),
.A2(n_947),
.B1(n_916),
.B2(n_930),
.Y(n_1033)
);

CKINVDCx8_ASAP7_75t_R g1034 ( 
.A(n_965),
.Y(n_1034)
);

OAI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_977),
.A2(n_929),
.B1(n_953),
.B2(n_951),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_977),
.A2(n_821),
.B1(n_931),
.B2(n_860),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_1012),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_965),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_959),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_1014),
.B(n_914),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_967),
.A2(n_931),
.B1(n_857),
.B2(n_811),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_969),
.B(n_905),
.Y(n_1042)
);

CKINVDCx11_ASAP7_75t_R g1043 ( 
.A(n_975),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_959),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_991),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_991),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_SL g1047 ( 
.A1(n_1006),
.A2(n_915),
.B1(n_914),
.B2(n_927),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_SL g1048 ( 
.A1(n_1015),
.A2(n_918),
.B(n_911),
.Y(n_1048)
);

BUFx4f_ASAP7_75t_L g1049 ( 
.A(n_984),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_974),
.Y(n_1050)
);

OAI21xp33_ASAP7_75t_L g1051 ( 
.A1(n_994),
.A2(n_905),
.B(n_910),
.Y(n_1051)
);

CKINVDCx16_ASAP7_75t_R g1052 ( 
.A(n_1005),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_967),
.A2(n_926),
.B1(n_842),
.B2(n_911),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_967),
.A2(n_926),
.B1(n_879),
.B2(n_949),
.Y(n_1054)
);

AOI22xp33_ASAP7_75t_L g1055 ( 
.A1(n_1007),
.A2(n_949),
.B1(n_956),
.B2(n_878),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_998),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_972),
.Y(n_1057)
);

OAI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1006),
.A2(n_910),
.B1(n_884),
.B2(n_902),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_1007),
.A2(n_956),
.B1(n_819),
.B2(n_820),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_986),
.B(n_843),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_986),
.A2(n_819),
.B1(n_820),
.B2(n_823),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_986),
.A2(n_823),
.B1(n_825),
.B2(n_827),
.Y(n_1062)
);

CKINVDCx14_ASAP7_75t_R g1063 ( 
.A(n_1005),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_974),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_964),
.A2(n_826),
.B1(n_825),
.B2(n_923),
.Y(n_1065)
);

CKINVDCx6p67_ASAP7_75t_R g1066 ( 
.A(n_989),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_990),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_SL g1068 ( 
.A1(n_1009),
.A2(n_933),
.B1(n_864),
.B2(n_868),
.Y(n_1068)
);

BUFx4f_ASAP7_75t_SL g1069 ( 
.A(n_989),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_992),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_1047),
.A2(n_984),
.B1(n_999),
.B2(n_964),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1023),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1029),
.A2(n_1004),
.B1(n_1011),
.B2(n_997),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1047),
.A2(n_1004),
.B1(n_1011),
.B2(n_997),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1024),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1028),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1033),
.A2(n_826),
.B1(n_999),
.B2(n_946),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1042),
.B(n_995),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_1064),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_1067),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1046),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_1026),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1039),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1030),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_1069),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1033),
.A2(n_882),
.B1(n_853),
.B2(n_861),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1040),
.A2(n_882),
.B1(n_861),
.B2(n_863),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1036),
.B(n_978),
.Y(n_1088)
);

OAI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_1035),
.A2(n_979),
.B1(n_934),
.B2(n_952),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1044),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1020),
.A2(n_863),
.B1(n_833),
.B2(n_827),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_SL g1092 ( 
.A1(n_1032),
.A2(n_933),
.B1(n_1018),
.B2(n_1049),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1051),
.A2(n_833),
.B1(n_852),
.B2(n_850),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1035),
.A2(n_992),
.B1(n_859),
.B2(n_849),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_SL g1095 ( 
.A1(n_1048),
.A2(n_1068),
.B(n_1041),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1068),
.A2(n_850),
.B1(n_852),
.B2(n_849),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1037),
.A2(n_859),
.B1(n_885),
.B2(n_805),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1045),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1070),
.Y(n_1099)
);

BUFx4f_ASAP7_75t_SL g1100 ( 
.A(n_1056),
.Y(n_1100)
);

OAI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1053),
.A2(n_982),
.B(n_885),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_SL g1102 ( 
.A1(n_1018),
.A2(n_1001),
.B1(n_961),
.B2(n_972),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_SL g1103 ( 
.A1(n_1018),
.A2(n_1001),
.B1(n_961),
.B2(n_1010),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1059),
.A2(n_813),
.B1(n_831),
.B2(n_979),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1043),
.Y(n_1105)
);

INVx5_ASAP7_75t_SL g1106 ( 
.A(n_1066),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1055),
.A2(n_831),
.B1(n_979),
.B2(n_845),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1060),
.A2(n_831),
.B1(n_845),
.B2(n_872),
.Y(n_1108)
);

OAI222xp33_ASAP7_75t_L g1109 ( 
.A1(n_1062),
.A2(n_841),
.B1(n_844),
.B2(n_836),
.C1(n_919),
.C2(n_937),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1054),
.A2(n_937),
.B1(n_973),
.B2(n_971),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1061),
.A2(n_831),
.B1(n_844),
.B2(n_841),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_1049),
.A2(n_1003),
.B1(n_864),
.B2(n_1016),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1058),
.A2(n_854),
.B1(n_801),
.B2(n_874),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1058),
.A2(n_854),
.B1(n_801),
.B2(n_874),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_1034),
.B(n_1008),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1065),
.A2(n_919),
.B1(n_864),
.B2(n_868),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_SL g1117 ( 
.A1(n_1069),
.A2(n_1003),
.B1(n_1016),
.B2(n_1008),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1065),
.A2(n_937),
.B1(n_1008),
.B2(n_987),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1038),
.B(n_868),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_SL g1120 ( 
.A1(n_1052),
.A2(n_1003),
.B1(n_980),
.B2(n_962),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_SL g1121 ( 
.A(n_1064),
.B(n_1025),
.Y(n_1121)
);

INVx6_ASAP7_75t_L g1122 ( 
.A(n_1064),
.Y(n_1122)
);

CKINVDCx14_ASAP7_75t_R g1123 ( 
.A(n_1063),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1021),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1021),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1019),
.A2(n_801),
.B1(n_873),
.B2(n_875),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1050),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1022),
.A2(n_801),
.B1(n_873),
.B2(n_875),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1050),
.A2(n_877),
.B(n_954),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1057),
.A2(n_987),
.B1(n_834),
.B2(n_980),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1027),
.A2(n_869),
.B1(n_996),
.B2(n_983),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1064),
.B(n_856),
.Y(n_1132)
);

OAI222xp33_ASAP7_75t_L g1133 ( 
.A1(n_1074),
.A2(n_883),
.B1(n_1002),
.B2(n_1027),
.C1(n_996),
.C2(n_983),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1072),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1092),
.A2(n_1002),
.B1(n_962),
.B2(n_976),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1074),
.A2(n_1031),
.B1(n_869),
.B2(n_1002),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1101),
.A2(n_1000),
.B1(n_993),
.B2(n_985),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_1079),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1073),
.A2(n_862),
.B1(n_1000),
.B2(n_993),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_SL g1140 ( 
.A1(n_1115),
.A2(n_976),
.B1(n_981),
.B2(n_958),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1075),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1073),
.A2(n_862),
.B1(n_1000),
.B2(n_993),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1071),
.A2(n_1077),
.B1(n_1088),
.B2(n_1086),
.Y(n_1143)
);

AND2x2_ASAP7_75t_SL g1144 ( 
.A(n_1077),
.B(n_985),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_SL g1145 ( 
.A1(n_1119),
.A2(n_958),
.B1(n_981),
.B2(n_993),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1128),
.A2(n_862),
.B1(n_1000),
.B2(n_985),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1118),
.A2(n_981),
.B1(n_958),
.B2(n_1025),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1078),
.B(n_1025),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1112),
.A2(n_862),
.B1(n_865),
.B2(n_935),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1095),
.A2(n_865),
.B1(n_862),
.B2(n_948),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_L g1151 ( 
.A(n_1087),
.B(n_865),
.C(n_935),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1076),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1107),
.A2(n_935),
.B1(n_948),
.B2(n_924),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1129),
.A2(n_1098),
.B(n_1090),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1126),
.A2(n_948),
.B1(n_924),
.B2(n_912),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1102),
.A2(n_880),
.B1(n_876),
.B2(n_925),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1103),
.A2(n_948),
.B1(n_924),
.B2(n_876),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_1080),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1097),
.A2(n_924),
.B1(n_880),
.B2(n_925),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1081),
.B(n_81),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1104),
.A2(n_880),
.B1(n_549),
.B2(n_557),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1083),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1116),
.A2(n_557),
.B1(n_558),
.B2(n_564),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1105),
.A2(n_564),
.B1(n_558),
.B2(n_557),
.Y(n_1164)
);

AOI222xp33_ASAP7_75t_L g1165 ( 
.A1(n_1116),
.A2(n_1089),
.B1(n_1094),
.B2(n_1100),
.C1(n_1096),
.C2(n_1109),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1089),
.A2(n_558),
.B1(n_564),
.B2(n_603),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1091),
.A2(n_603),
.B1(n_610),
.B2(n_526),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1099),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1100),
.A2(n_1094),
.B1(n_1111),
.B2(n_1084),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1082),
.A2(n_603),
.B1(n_610),
.B2(n_526),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1108),
.A2(n_921),
.B(n_610),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1120),
.A2(n_610),
.B1(n_526),
.B2(n_40),
.Y(n_1172)
);

INVx4_ASAP7_75t_R g1173 ( 
.A(n_1085),
.Y(n_1173)
);

OAI222xp33_ASAP7_75t_L g1174 ( 
.A1(n_1131),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.C1(n_41),
.C2(n_42),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_1113),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.C(n_43),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1117),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1132),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1110),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1114),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1106),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1123),
.A2(n_1106),
.B1(n_1130),
.B2(n_1093),
.Y(n_1181)
);

CKINVDCx6p67_ASAP7_75t_R g1182 ( 
.A(n_1079),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1124),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1106),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1127),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1125),
.B(n_83),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1122),
.A2(n_60),
.B1(n_61),
.B2(n_334),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1122),
.A2(n_60),
.B1(n_61),
.B2(n_84),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1122),
.A2(n_85),
.B1(n_86),
.B2(n_91),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1079),
.B(n_1121),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1079),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1101),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_1192)
);

OA21x2_ASAP7_75t_L g1193 ( 
.A1(n_1154),
.A2(n_1171),
.B(n_1150),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1133),
.B(n_108),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1134),
.B(n_109),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_L g1196 ( 
.A(n_1187),
.B(n_111),
.C(n_112),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1141),
.B(n_113),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1163),
.A2(n_114),
.B(n_116),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1165),
.B(n_123),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1148),
.B(n_124),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1152),
.B(n_1162),
.Y(n_1201)
);

NAND4xp25_ASAP7_75t_L g1202 ( 
.A(n_1184),
.B(n_130),
.C(n_131),
.D(n_133),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1136),
.A2(n_134),
.B1(n_136),
.B2(n_141),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1168),
.B(n_143),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1158),
.B(n_147),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1144),
.B(n_333),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1183),
.B(n_148),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1144),
.B(n_1181),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1187),
.B(n_150),
.C(n_151),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1143),
.B(n_154),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1147),
.B(n_157),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1145),
.B(n_159),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1140),
.B(n_161),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1188),
.B(n_164),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1175),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1174),
.A2(n_172),
.B(n_175),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1169),
.B(n_178),
.Y(n_1217)
);

AOI221xp5_ASAP7_75t_L g1218 ( 
.A1(n_1177),
.A2(n_1180),
.B1(n_1178),
.B2(n_1179),
.C(n_1176),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1137),
.B(n_1160),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1136),
.B(n_183),
.Y(n_1220)
);

NAND3xp33_ASAP7_75t_L g1221 ( 
.A(n_1188),
.B(n_185),
.C(n_187),
.Y(n_1221)
);

AOI221xp5_ASAP7_75t_L g1222 ( 
.A1(n_1185),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.C(n_194),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1186),
.B(n_196),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1137),
.B(n_197),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1139),
.B(n_198),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1142),
.B(n_1190),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1163),
.B(n_199),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1146),
.B(n_201),
.Y(n_1228)
);

NAND4xp25_ASAP7_75t_L g1229 ( 
.A(n_1164),
.B(n_202),
.C(n_204),
.D(n_206),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1138),
.B(n_208),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1151),
.B(n_209),
.Y(n_1231)
);

OAI221xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1192),
.A2(n_211),
.B1(n_212),
.B2(n_218),
.C(n_220),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1138),
.B(n_221),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1191),
.B(n_222),
.C(n_225),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1172),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1191),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1166),
.B(n_1149),
.Y(n_1237)
);

OA211x2_ASAP7_75t_L g1238 ( 
.A1(n_1153),
.A2(n_240),
.B(n_241),
.C(n_242),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1189),
.B(n_243),
.C(n_244),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1157),
.A2(n_246),
.B(n_247),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1208),
.B(n_1182),
.Y(n_1241)
);

OA211x2_ASAP7_75t_L g1242 ( 
.A1(n_1194),
.A2(n_1159),
.B(n_1161),
.C(n_1155),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1201),
.B(n_1135),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_1205),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1195),
.B(n_1173),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1199),
.A2(n_1156),
.B1(n_1170),
.B2(n_1167),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1226),
.B(n_250),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1195),
.B(n_251),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1199),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_1249)
);

NAND3xp33_ASAP7_75t_L g1250 ( 
.A(n_1216),
.B(n_257),
.C(n_258),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1219),
.B(n_260),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1193),
.B(n_261),
.Y(n_1252)
);

INVx5_ASAP7_75t_L g1253 ( 
.A(n_1230),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1197),
.B(n_263),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1206),
.B(n_264),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1193),
.B(n_265),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1193),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1197),
.B(n_270),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1194),
.B(n_271),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1204),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1196),
.B(n_274),
.C(n_275),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1218),
.A2(n_282),
.B1(n_283),
.B2(n_285),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1200),
.B(n_286),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1230),
.Y(n_1264)
);

NAND4xp75_ASAP7_75t_L g1265 ( 
.A(n_1238),
.B(n_287),
.C(n_289),
.D(n_291),
.Y(n_1265)
);

NOR3xp33_ASAP7_75t_L g1266 ( 
.A(n_1209),
.B(n_292),
.C(n_293),
.Y(n_1266)
);

NAND3xp33_ASAP7_75t_L g1267 ( 
.A(n_1221),
.B(n_296),
.C(n_297),
.Y(n_1267)
);

NAND4xp75_ASAP7_75t_L g1268 ( 
.A(n_1242),
.B(n_1213),
.C(n_1214),
.D(n_1231),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1260),
.B(n_1207),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1243),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1257),
.Y(n_1271)
);

NAND4xp75_ASAP7_75t_SL g1272 ( 
.A(n_1255),
.B(n_1212),
.C(n_1214),
.D(n_1211),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1260),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1264),
.B(n_1212),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1244),
.B(n_1237),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1253),
.B(n_1233),
.Y(n_1276)
);

XOR2x2_ASAP7_75t_L g1277 ( 
.A(n_1250),
.B(n_1234),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1253),
.B(n_1237),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1252),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1241),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1253),
.Y(n_1281)
);

XNOR2xp5_ASAP7_75t_L g1282 ( 
.A(n_1245),
.B(n_1202),
.Y(n_1282)
);

AND4x1_ASAP7_75t_L g1283 ( 
.A(n_1249),
.B(n_1239),
.C(n_1236),
.D(n_1222),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1256),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1245),
.B(n_1233),
.Y(n_1285)
);

XOR2x2_ASAP7_75t_L g1286 ( 
.A(n_1259),
.B(n_1232),
.Y(n_1286)
);

INVx4_ASAP7_75t_L g1287 ( 
.A(n_1248),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1273),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1270),
.B(n_1279),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1284),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1273),
.Y(n_1291)
);

XOR2x2_ASAP7_75t_L g1292 ( 
.A(n_1286),
.B(n_1265),
.Y(n_1292)
);

XOR2x2_ASAP7_75t_L g1293 ( 
.A(n_1286),
.B(n_1267),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1271),
.Y(n_1294)
);

XNOR2x2_ASAP7_75t_L g1295 ( 
.A(n_1268),
.B(n_1213),
.Y(n_1295)
);

XNOR2xp5_ASAP7_75t_L g1296 ( 
.A(n_1282),
.B(n_1248),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1276),
.B(n_1251),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1271),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1269),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1278),
.Y(n_1300)
);

XNOR2xp5_ASAP7_75t_L g1301 ( 
.A(n_1282),
.B(n_1247),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1294),
.Y(n_1302)
);

OA22x2_ASAP7_75t_L g1303 ( 
.A1(n_1301),
.A2(n_1287),
.B1(n_1280),
.B2(n_1274),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1292),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1297),
.B(n_1276),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1290),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1290),
.Y(n_1307)
);

OA22x2_ASAP7_75t_L g1308 ( 
.A1(n_1296),
.A2(n_1287),
.B1(n_1274),
.B2(n_1285),
.Y(n_1308)
);

XOR2x2_ASAP7_75t_L g1309 ( 
.A(n_1293),
.B(n_1272),
.Y(n_1309)
);

OA22x2_ASAP7_75t_L g1310 ( 
.A1(n_1295),
.A2(n_1287),
.B1(n_1285),
.B2(n_1275),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1292),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1294),
.Y(n_1312)
);

XNOR2xp5_ASAP7_75t_L g1313 ( 
.A(n_1293),
.B(n_1268),
.Y(n_1313)
);

AOI22x1_ASAP7_75t_L g1314 ( 
.A1(n_1300),
.A2(n_1277),
.B1(n_1227),
.B2(n_1198),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1289),
.A2(n_1281),
.B1(n_1277),
.B2(n_1220),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1298),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1302),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1308),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1302),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1306),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1307),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1312),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1303),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1312),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1316),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1311),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1317),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1317),
.Y(n_1328)
);

NAND4xp75_ASAP7_75t_L g1329 ( 
.A(n_1320),
.B(n_1313),
.C(n_1311),
.D(n_1304),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1323),
.A2(n_1304),
.B1(n_1310),
.B2(n_1309),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1321),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1318),
.A2(n_1314),
.B1(n_1310),
.B2(n_1315),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1326),
.A2(n_1308),
.B1(n_1303),
.B2(n_1266),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1327),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1330),
.A2(n_1281),
.B1(n_1305),
.B2(n_1325),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1328),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1332),
.A2(n_1319),
.B(n_1322),
.C(n_1324),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1331),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1333),
.A2(n_1329),
.B1(n_1331),
.B2(n_1319),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1327),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1339),
.A2(n_1324),
.B1(n_1299),
.B2(n_1298),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1334),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1335),
.A2(n_1240),
.B1(n_1261),
.B2(n_1262),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1338),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1336),
.B(n_1291),
.Y(n_1345)
);

NOR2x1_ASAP7_75t_L g1346 ( 
.A(n_1337),
.B(n_1229),
.Y(n_1346)
);

NOR2x1_ASAP7_75t_L g1347 ( 
.A(n_1340),
.B(n_1288),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1346),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1341),
.B(n_1283),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1347),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1344),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1342),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1345),
.Y(n_1353)
);

AND4x1_ASAP7_75t_L g1354 ( 
.A(n_1352),
.B(n_1343),
.C(n_1235),
.D(n_1217),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1350),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1351),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1348),
.A2(n_1258),
.B1(n_1254),
.B2(n_1210),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1349),
.A2(n_1246),
.B1(n_1215),
.B2(n_1263),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1355),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1356),
.A2(n_1353),
.B1(n_1223),
.B2(n_1203),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1354),
.Y(n_1361)
);

OA22x2_ASAP7_75t_L g1362 ( 
.A1(n_1357),
.A2(n_1231),
.B1(n_1223),
.B2(n_1224),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1358),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1359),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1361),
.A2(n_1227),
.B1(n_1225),
.B2(n_1228),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1363),
.Y(n_1366)
);

AO22x1_ASAP7_75t_L g1367 ( 
.A1(n_1362),
.A2(n_298),
.B1(n_300),
.B2(n_301),
.Y(n_1367)
);

OAI22x1_ASAP7_75t_L g1368 ( 
.A1(n_1360),
.A2(n_302),
.B1(n_304),
.B2(n_306),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1366),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1364),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1368),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1367),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1369),
.A2(n_1370),
.B1(n_1371),
.B2(n_1372),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1369),
.A2(n_1365),
.B1(n_310),
.B2(n_311),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1373),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1374),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1375),
.A2(n_308),
.B1(n_314),
.B2(n_316),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1377),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1378),
.A2(n_1376),
.B1(n_318),
.B2(n_320),
.C(n_321),
.Y(n_1379)
);

AOI211xp5_ASAP7_75t_L g1380 ( 
.A1(n_1379),
.A2(n_317),
.B(n_323),
.C(n_325),
.Y(n_1380)
);


endmodule