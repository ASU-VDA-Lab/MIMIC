module fake_jpeg_5737_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_4),
.B(n_6),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_26),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_27),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_28),
.B1(n_14),
.B2(n_9),
.Y(n_37)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_25),
.Y(n_31)
);

NOR3xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_16),
.C(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_5),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_11),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_32),
.C(n_20),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_38),
.B1(n_30),
.B2(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_30),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_40),
.C(n_42),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_48),
.C(n_43),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_44),
.B(n_46),
.C(n_41),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_61),
.B1(n_55),
.B2(n_52),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_53),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_54),
.B(n_44),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_60),
.C(n_62),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_46),
.B1(n_13),
.B2(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_13),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_51),
.C(n_15),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_65),
.Y(n_69)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.C(n_8),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_8),
.Y(n_72)
);


endmodule