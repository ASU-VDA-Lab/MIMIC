module fake_ibex_1974_n_14 (n_3, n_1, n_4, n_2, n_0, n_14);

input n_3;
input n_1;
input n_4;
input n_2;
input n_0;

output n_14;



endmodule