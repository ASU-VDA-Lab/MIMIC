module fake_jpeg_2978_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_54),
.Y(n_62)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_42),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_67),
.Y(n_73)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_39),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_55),
.Y(n_76)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_48),
.C(n_39),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_44),
.B1(n_48),
.B2(n_53),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_52),
.B1(n_55),
.B2(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_52),
.B1(n_57),
.B2(n_43),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_41),
.B(n_37),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_65),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_73),
.B(n_72),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_87),
.B(n_47),
.Y(n_99)
);

OA21x2_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_60),
.B(n_47),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_53),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_15),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_49),
.C(n_40),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_1),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_93),
.B(n_95),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_0),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_47),
.B1(n_45),
.B2(n_3),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_97),
.A2(n_103),
.B1(n_8),
.B2(n_11),
.Y(n_123)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_1),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_107),
.C(n_108),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_2),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_110),
.B(n_112),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_5),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_21),
.B1(n_33),
.B2(n_30),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_87),
.B(n_88),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_122),
.B(n_124),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_83),
.B(n_90),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_109),
.B(n_97),
.Y(n_126)
);

AOI221xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_103),
.B1(n_111),
.B2(n_26),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_13),
.B(n_16),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_111),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_120),
.B(n_125),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.C(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_131),
.B1(n_114),
.B2(n_117),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_130),
.B(n_121),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_129),
.B(n_122),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_113),
.C(n_24),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_22),
.Y(n_141)
);


endmodule