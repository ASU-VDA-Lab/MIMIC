module fake_ariane_2271_n_1668 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1668);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1668;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_85),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_139),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_0),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_46),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_55),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_127),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_29),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_48),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_9),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_121),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_34),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_93),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_103),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_69),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_61),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_25),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_77),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_60),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_19),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_29),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_2),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_136),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_14),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_35),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_34),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_40),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_90),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_72),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_17),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_49),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_4),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_107),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_1),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_14),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_37),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_73),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_71),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_33),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_131),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_57),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_62),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_94),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_13),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_81),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_70),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_25),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_109),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_116),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_78),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_27),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_100),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_28),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_132),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_75),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_2),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_147),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_63),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_0),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_112),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_130),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_87),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_122),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_1),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_115),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_42),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_110),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_52),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_11),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_54),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_145),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_58),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_68),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_44),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_74),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_91),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_19),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_11),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_114),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_18),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_146),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_64),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_10),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_26),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_89),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_96),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_124),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_129),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_15),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_6),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_118),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_21),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_88),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_111),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_123),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_92),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_59),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_39),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_128),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_137),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_48),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_53),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_120),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_99),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_28),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_41),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_105),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_12),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_7),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_41),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_22),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_20),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_22),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_143),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_43),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_36),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_15),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_20),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_32),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_138),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_43),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_23),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_24),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_18),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_3),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_47),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_83),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_7),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_133),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_67),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_104),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_51),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_84),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_213),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_198),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_161),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_177),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_192),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_153),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_168),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_226),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_271),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_271),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_152),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_174),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_152),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_246),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_198),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_232),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_176),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_180),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_154),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_181),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_274),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_182),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_179),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g332 ( 
.A(n_195),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_196),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_185),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_169),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_204),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_188),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_190),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_210),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_268),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_221),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_235),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_237),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_250),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_258),
.Y(n_347)
);

INVxp33_ASAP7_75t_SL g348 ( 
.A(n_159),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_279),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_232),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_157),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_178),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_160),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_186),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_156),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_187),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_189),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_209),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_191),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_214),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_215),
.Y(n_363)
);

BUFx6f_ASAP7_75t_SL g364 ( 
.A(n_156),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_220),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_208),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_295),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_305),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_295),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_313),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_296),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_315),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_303),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_296),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_298),
.B(n_276),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_309),
.B(n_175),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_299),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_298),
.B(n_276),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_307),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_311),
.B(n_225),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_316),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_316),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_354),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_317),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_318),
.Y(n_388)
);

BUFx8_ASAP7_75t_L g389 ( 
.A(n_364),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_299),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_304),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_300),
.A2(n_185),
.B1(n_201),
.B2(n_240),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_304),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_360),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_294),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_326),
.B(n_227),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_334),
.A2(n_201),
.B1(n_170),
.B2(n_160),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_326),
.B(n_238),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_356),
.B(n_294),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_302),
.A2(n_163),
.B1(n_170),
.B2(n_173),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_329),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_358),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_320),
.Y(n_413)
);

OA21x2_ASAP7_75t_L g414 ( 
.A1(n_358),
.A2(n_293),
.B(n_244),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_359),
.B(n_280),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_308),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_332),
.B(n_156),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_359),
.B(n_184),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_337),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_320),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_326),
.B(n_242),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_326),
.B(n_254),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_350),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_297),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_350),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_335),
.B(n_260),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_357),
.A2(n_163),
.B1(n_173),
.B2(n_275),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_362),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_363),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_363),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_308),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g434 ( 
.A(n_361),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_310),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_367),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_301),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_367),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_416),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_375),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_385),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_306),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_368),
.B(n_327),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_416),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_385),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_370),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_434),
.B(n_348),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_385),
.B(n_365),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_385),
.B(n_314),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_419),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_400),
.B(n_324),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_364),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_412),
.B(n_340),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_372),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_429),
.Y(n_468)
);

INVx8_ASAP7_75t_L g469 ( 
.A(n_400),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_400),
.A2(n_364),
.B1(n_355),
.B2(n_339),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_416),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_430),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_376),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_430),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_400),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_416),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_431),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_395),
.B(n_150),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_408),
.B(n_349),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_432),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_408),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_408),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_390),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_406),
.B(n_151),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_411),
.B(n_150),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

AOI21x1_ASAP7_75t_L g492 ( 
.A1(n_414),
.A2(n_267),
.B(n_263),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_432),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_409),
.B(n_325),
.C(n_322),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_394),
.B(n_341),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_SL g496 ( 
.A(n_411),
.B(n_275),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_381),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_392),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_408),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_409),
.A2(n_277),
.B1(n_278),
.B2(n_269),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_436),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_436),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_369),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_421),
.B(n_344),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_392),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_422),
.B(n_323),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_397),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_423),
.B(n_323),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_369),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_415),
.B(n_328),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_423),
.B(n_277),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_390),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_371),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_415),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_390),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_415),
.B(n_328),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_371),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_378),
.B(n_330),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_413),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_390),
.Y(n_522)
);

AND3x2_ASAP7_75t_L g523 ( 
.A(n_415),
.B(n_333),
.C(n_330),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_373),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_414),
.A2(n_233),
.B1(n_255),
.B2(n_257),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g527 ( 
.A(n_394),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_433),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_414),
.A2(n_233),
.B1(n_255),
.B2(n_257),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_389),
.B(n_155),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_418),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_413),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_373),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_435),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_382),
.B(n_333),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_374),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_418),
.B(n_336),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_418),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_424),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_403),
.B(n_336),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_374),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_389),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_383),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_410),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_426),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_425),
.Y(n_549)
);

BUFx6f_ASAP7_75t_SL g550 ( 
.A(n_377),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_389),
.B(n_377),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_403),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_403),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_377),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_407),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_428),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_383),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_407),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_407),
.Y(n_559)
);

INVxp33_ASAP7_75t_SL g560 ( 
.A(n_428),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_414),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_407),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_380),
.B(n_278),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_L g564 ( 
.A(n_384),
.B(n_151),
.Y(n_564)
);

INVx8_ASAP7_75t_L g565 ( 
.A(n_380),
.Y(n_565)
);

OAI21xp33_ASAP7_75t_SL g566 ( 
.A1(n_384),
.A2(n_352),
.B(n_343),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_420),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_420),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_380),
.A2(n_257),
.B1(n_255),
.B2(n_288),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_380),
.B(n_342),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_386),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_402),
.B(n_398),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_386),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_387),
.B(n_155),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_420),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_420),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_387),
.Y(n_577)
);

BUFx4f_ASAP7_75t_L g578 ( 
.A(n_398),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_388),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_388),
.Y(n_580)
);

INVx8_ASAP7_75t_L g581 ( 
.A(n_399),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_449),
.B(n_458),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_443),
.A2(n_391),
.B1(n_396),
.B2(n_393),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_581),
.Y(n_584)
);

INVx8_ASAP7_75t_L g585 ( 
.A(n_469),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_520),
.B(n_399),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_507),
.B(n_391),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_537),
.B(n_393),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_477),
.A2(n_396),
.B1(n_158),
.B2(n_172),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_575),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_575),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_477),
.B(n_158),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_528),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_485),
.B(n_162),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_458),
.B(n_162),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_556),
.A2(n_560),
.B1(n_527),
.B2(n_495),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_471),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_485),
.B(n_164),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_486),
.B(n_164),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_458),
.B(n_540),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_486),
.A2(n_172),
.B1(n_171),
.B2(n_217),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_442),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_540),
.B(n_165),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_499),
.B(n_516),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_463),
.B(n_343),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_540),
.B(n_165),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_439),
.B(n_216),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_444),
.B(n_509),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_581),
.B(n_166),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_528),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_509),
.B(n_166),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_554),
.B(n_532),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_505),
.B(n_457),
.C(n_501),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_554),
.B(n_171),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_463),
.B(n_345),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_489),
.A2(n_290),
.B(n_291),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_528),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_516),
.B(n_461),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_457),
.B(n_233),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_554),
.B(n_217),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_532),
.B(n_518),
.Y(n_622)
);

AND2x2_ASAP7_75t_SL g623 ( 
.A(n_556),
.B(n_184),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_469),
.B(n_231),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_570),
.B(n_346),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_560),
.A2(n_495),
.B1(n_447),
.B2(n_462),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_581),
.B(n_234),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_455),
.B(n_247),
.Y(n_628)
);

BUFx5_ASAP7_75t_L g629 ( 
.A(n_454),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_469),
.B(n_248),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_469),
.B(n_261),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_452),
.A2(n_273),
.B1(n_287),
.B2(n_286),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_581),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_528),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_550),
.A2(n_183),
.B1(n_292),
.B2(n_149),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_497),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_529),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_565),
.B(n_265),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_565),
.B(n_266),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_482),
.B(n_270),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_539),
.B(n_347),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_490),
.B(n_565),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_500),
.B(n_347),
.Y(n_643)
);

BUFx8_ASAP7_75t_L g644 ( 
.A(n_549),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_500),
.B(n_351),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_539),
.B(n_351),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_438),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_565),
.B(n_272),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_459),
.B(n_281),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_563),
.A2(n_229),
.B1(n_194),
.B2(n_197),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_454),
.B(n_352),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_529),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_529),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_483),
.B(n_284),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_470),
.B(n_288),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_551),
.B(n_288),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_444),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_574),
.B(n_3),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_464),
.B(n_199),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_464),
.B(n_200),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_549),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_523),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_468),
.B(n_184),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_468),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_473),
.B(n_202),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_473),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_446),
.B(n_5),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_547),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_529),
.Y(n_669)
);

INVxp33_ASAP7_75t_L g670 ( 
.A(n_445),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_474),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_529),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_511),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_476),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_476),
.B(n_203),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_494),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_479),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_572),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_578),
.A2(n_228),
.B1(n_264),
.B2(n_262),
.Y(n_679)
);

OAI21xp33_ASAP7_75t_L g680 ( 
.A1(n_479),
.A2(n_312),
.B(n_224),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_481),
.B(n_205),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_451),
.B(n_312),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_559),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_559),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_493),
.B(n_5),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_481),
.B(n_222),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_533),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_484),
.B(n_502),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_578),
.B(n_230),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_578),
.B(n_219),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_533),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_484),
.B(n_151),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_545),
.B(n_206),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_533),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_572),
.B(n_6),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_502),
.A2(n_259),
.B1(n_167),
.B2(n_193),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_496),
.B(n_236),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_545),
.B(n_8),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_541),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_SL g700 ( 
.A(n_572),
.B(n_561),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_503),
.B(n_239),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_503),
.B(n_8),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_571),
.B(n_573),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_580),
.B(n_218),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_504),
.B(n_243),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_438),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_513),
.B(n_253),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_504),
.B(n_252),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_542),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_541),
.Y(n_710)
);

NAND2x1_ASAP7_75t_L g711 ( 
.A(n_517),
.B(n_259),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_510),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_541),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_510),
.B(n_211),
.Y(n_714)
);

BUFx6f_ASAP7_75t_SL g715 ( 
.A(n_572),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_515),
.B(n_251),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_566),
.A2(n_249),
.B(n_245),
.C(n_259),
.Y(n_717)
);

NAND3xp33_ASAP7_75t_L g718 ( 
.A(n_569),
.B(n_259),
.C(n_212),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_515),
.B(n_151),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_519),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_519),
.B(n_151),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_531),
.B(n_10),
.C(n_12),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_525),
.B(n_151),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_555),
.B(n_13),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_536),
.Y(n_725)
);

OAI221xp5_ASAP7_75t_L g726 ( 
.A1(n_526),
.A2(n_212),
.B1(n_207),
.B2(n_193),
.C(n_167),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_525),
.A2(n_151),
.B1(n_212),
.B2(n_193),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_534),
.B(n_212),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_536),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_438),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_555),
.B(n_16),
.Y(n_731)
);

NAND2x1p5_ASAP7_75t_L g732 ( 
.A(n_555),
.B(n_207),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_538),
.B(n_207),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_538),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_544),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_544),
.B(n_193),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_623),
.B(n_558),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_734),
.A2(n_577),
.B1(n_546),
.B2(n_557),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_608),
.B(n_530),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_623),
.B(n_676),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_608),
.B(n_546),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_657),
.B(n_557),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_598),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_629),
.B(n_438),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_725),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_729),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_668),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_603),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_628),
.B(n_577),
.Y(n_749)
);

AND2x6_ASAP7_75t_SL g750 ( 
.A(n_695),
.B(n_521),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_628),
.B(n_579),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_629),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_629),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_585),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_585),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_700),
.A2(n_564),
.B1(n_562),
.B2(n_558),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_588),
.B(n_586),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_629),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_661),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_644),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_629),
.Y(n_761)
);

AND2x4_ASAP7_75t_SL g762 ( 
.A(n_643),
.B(n_558),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_657),
.B(n_579),
.Y(n_763)
);

AO22x1_ASAP7_75t_L g764 ( 
.A1(n_695),
.A2(n_562),
.B1(n_561),
.B2(n_524),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_664),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_629),
.Y(n_766)
);

BUFx8_ASAP7_75t_L g767 ( 
.A(n_715),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_585),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_606),
.B(n_562),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_584),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_687),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_620),
.A2(n_561),
.B1(n_568),
.B2(n_567),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_633),
.B(n_438),
.Y(n_773)
);

AND2x6_ASAP7_75t_SL g774 ( 
.A(n_640),
.B(n_16),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_R g775 ( 
.A(n_644),
.B(n_489),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_597),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_676),
.B(n_614),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_709),
.B(n_441),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_666),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_616),
.B(n_734),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_633),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_587),
.B(n_524),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_688),
.A2(n_564),
.B(n_568),
.C(n_567),
.Y(n_784)
);

BUFx10_ASAP7_75t_L g785 ( 
.A(n_648),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_584),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_678),
.B(n_441),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_671),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_SL g789 ( 
.A(n_612),
.B(n_17),
.C(n_21),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_649),
.B(n_535),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_709),
.B(n_441),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_584),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_609),
.B(n_535),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_649),
.B(n_576),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_691),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_626),
.A2(n_543),
.B1(n_548),
.B2(n_453),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_654),
.B(n_576),
.Y(n_797)
);

AND3x2_ASAP7_75t_SL g798 ( 
.A(n_715),
.B(n_553),
.C(n_552),
.Y(n_798)
);

AND2x6_ASAP7_75t_SL g799 ( 
.A(n_640),
.B(n_23),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_654),
.B(n_553),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_584),
.B(n_480),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_694),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_706),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_699),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_674),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_596),
.A2(n_543),
.B1(n_548),
.B2(n_466),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_625),
.B(n_552),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_656),
.A2(n_478),
.B1(n_437),
.B2(n_440),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_647),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_SL g810 ( 
.A(n_632),
.B(n_24),
.C(n_26),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_619),
.B(n_480),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_710),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_706),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_656),
.A2(n_475),
.B1(n_465),
.B2(n_466),
.Y(n_814)
);

AO22x1_ASAP7_75t_L g815 ( 
.A1(n_670),
.A2(n_448),
.B1(n_460),
.B2(n_472),
.Y(n_815)
);

BUFx12f_ASAP7_75t_L g816 ( 
.A(n_643),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_677),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_590),
.B(n_448),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_673),
.B(n_437),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_712),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_688),
.B(n_480),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_642),
.A2(n_460),
.B1(n_472),
.B2(n_517),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_720),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_645),
.B(n_517),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_735),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_726),
.A2(n_450),
.B1(n_475),
.B2(n_512),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_662),
.B(n_480),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_703),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_641),
.B(n_488),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_646),
.A2(n_453),
.B(n_465),
.C(n_467),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_658),
.A2(n_467),
.B1(n_478),
.B2(n_512),
.Y(n_831)
);

AND2x4_ASAP7_75t_SL g832 ( 
.A(n_698),
.B(n_480),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_713),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_658),
.A2(n_498),
.B1(n_508),
.B2(n_506),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_706),
.B(n_730),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_622),
.B(n_498),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_713),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_591),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_635),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_682),
.Y(n_840)
);

AO21x1_ASAP7_75t_L g841 ( 
.A1(n_702),
.A2(n_492),
.B(n_506),
.Y(n_841)
);

INVx5_ASAP7_75t_L g842 ( 
.A(n_706),
.Y(n_842)
);

AND2x2_ASAP7_75t_SL g843 ( 
.A(n_722),
.B(n_167),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_593),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_730),
.B(n_605),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_648),
.B(n_514),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_730),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_651),
.B(n_514),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_702),
.B(n_522),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_SL g850 ( 
.A(n_722),
.B(n_27),
.C(n_30),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_642),
.B(n_522),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_647),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_583),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_582),
.A2(n_522),
.B(n_491),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_611),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_667),
.B(n_522),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_730),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_618),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_667),
.B(n_522),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_724),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_634),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_663),
.Y(n_862)
);

OAI22xp33_ASAP7_75t_L g863 ( 
.A1(n_602),
.A2(n_491),
.B1(n_487),
.B2(n_456),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_637),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_683),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_R g866 ( 
.A(n_610),
.B(n_492),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_601),
.B(n_456),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_663),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_685),
.B(n_491),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_685),
.B(n_491),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_592),
.B(n_491),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_704),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_594),
.B(n_487),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_652),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_653),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_684),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_669),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_653),
.B(n_487),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_599),
.B(n_487),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_627),
.A2(n_487),
.B1(n_456),
.B2(n_167),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_672),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_689),
.A2(n_456),
.B(n_66),
.Y(n_882)
);

NOR2x2_ASAP7_75t_L g883 ( 
.A(n_624),
.B(n_30),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_719),
.Y(n_884)
);

AND2x6_ASAP7_75t_SL g885 ( 
.A(n_731),
.B(n_600),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_647),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_589),
.B(n_659),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_660),
.B(n_456),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_665),
.B(n_31),
.Y(n_889)
);

AOI211xp5_ASAP7_75t_L g890 ( 
.A1(n_655),
.A2(n_31),
.B(n_32),
.C(n_35),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_647),
.B(n_36),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_721),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_675),
.B(n_37),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_723),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_731),
.B(n_38),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_711),
.Y(n_896)
);

O2A1O1Ixp5_ASAP7_75t_L g897 ( 
.A1(n_690),
.A2(n_38),
.B(n_39),
.C(n_42),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_693),
.B(n_44),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_733),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_736),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_L g901 ( 
.A(n_630),
.B(n_45),
.C(n_46),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_681),
.Y(n_902)
);

BUFx12f_ASAP7_75t_L g903 ( 
.A(n_663),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_686),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_732),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_613),
.A2(n_98),
.B(n_141),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_732),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_663),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_697),
.Y(n_909)
);

NAND2x1p5_ASAP7_75t_L g910 ( 
.A(n_638),
.B(n_97),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_663),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_741),
.B(n_650),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_778),
.A2(n_617),
.B(n_714),
.C(n_708),
.Y(n_913)
);

AND2x2_ASAP7_75t_SL g914 ( 
.A(n_843),
.B(n_740),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_757),
.A2(n_692),
.B(n_615),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_747),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_828),
.B(n_716),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_747),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_748),
.B(n_718),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_743),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_749),
.A2(n_621),
.B(n_705),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_740),
.B(n_701),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_817),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_849),
.A2(n_639),
.B(n_631),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_751),
.A2(n_595),
.B(n_604),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_838),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_754),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_744),
.A2(n_607),
.B(n_707),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_777),
.B(n_679),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_778),
.B(n_680),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_742),
.B(n_717),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_840),
.B(n_727),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_784),
.A2(n_728),
.B(n_696),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_754),
.B(n_696),
.Y(n_934)
);

OA21x2_ASAP7_75t_L g935 ( 
.A1(n_841),
.A2(n_101),
.B(n_140),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_744),
.A2(n_80),
.B(n_117),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_817),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_784),
.A2(n_45),
.B(n_47),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_820),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_793),
.B(n_56),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_776),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_853),
.A2(n_65),
.B1(n_76),
.B2(n_79),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_739),
.A2(n_102),
.B(n_108),
.C(n_113),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_895),
.A2(n_142),
.B(n_887),
.C(n_902),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_R g945 ( 
.A(n_760),
.B(n_759),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_820),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_872),
.B(n_839),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_823),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_737),
.A2(n_843),
.B(n_904),
.C(n_895),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_763),
.B(n_737),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_754),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_856),
.A2(n_869),
.B(n_859),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_738),
.A2(n_823),
.B1(n_825),
.B2(n_780),
.Y(n_953)
);

AOI21x1_ASAP7_75t_L g954 ( 
.A1(n_811),
.A2(n_821),
.B(n_845),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_765),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_825),
.B(n_788),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_754),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_785),
.B(n_816),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_SL g959 ( 
.A(n_890),
.B(n_901),
.C(n_810),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_865),
.A2(n_876),
.B1(n_806),
.B2(n_824),
.Y(n_960)
);

BUFx8_ASAP7_75t_L g961 ( 
.A(n_776),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_805),
.B(n_762),
.Y(n_962)
);

OR2x6_ASAP7_75t_SL g963 ( 
.A(n_760),
.B(n_889),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_SL g964 ( 
.A(n_903),
.B(n_782),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_785),
.B(n_755),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_755),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_750),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_785),
.A2(n_824),
.B1(n_762),
.B2(n_827),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_860),
.A2(n_769),
.B1(n_783),
.B2(n_893),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_807),
.A2(n_829),
.B1(n_870),
.B2(n_791),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_767),
.Y(n_971)
);

BUFx10_ASAP7_75t_L g972 ( 
.A(n_885),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_768),
.B(n_827),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_779),
.A2(n_791),
.B(n_790),
.C(n_794),
.Y(n_974)
);

AND2x4_ASAP7_75t_SL g975 ( 
.A(n_827),
.B(n_782),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_821),
.A2(n_800),
.B(n_797),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_745),
.Y(n_977)
);

NAND2x1p5_ASAP7_75t_L g978 ( 
.A(n_768),
.B(n_813),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_779),
.A2(n_846),
.B(n_756),
.C(n_884),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_787),
.B(n_819),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_767),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_894),
.A2(n_818),
.B(n_911),
.C(n_908),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_782),
.Y(n_983)
);

INVx1_ASAP7_75t_SL g984 ( 
.A(n_832),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_832),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_888),
.A2(n_879),
.B(n_873),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_787),
.B(n_909),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_789),
.B(n_787),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_775),
.Y(n_989)
);

INVx3_ASAP7_75t_SL g990 ( 
.A(n_883),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_770),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_818),
.A2(n_911),
.B(n_908),
.C(n_830),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_772),
.B(n_813),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_764),
.B(n_796),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_774),
.Y(n_995)
);

AO21x1_ASAP7_75t_L g996 ( 
.A1(n_845),
.A2(n_851),
.B(n_891),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_833),
.B(n_837),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_871),
.A2(n_766),
.B(n_752),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_833),
.B(n_837),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_813),
.B(n_842),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_771),
.B(n_795),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_836),
.B(n_771),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_746),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_908),
.A2(n_911),
.B(n_850),
.C(n_897),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_848),
.A2(n_892),
.B(n_854),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_892),
.B(n_812),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_891),
.A2(n_898),
.B(n_822),
.Y(n_1007)
);

BUFx2_ASAP7_75t_SL g1008 ( 
.A(n_813),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_752),
.A2(n_753),
.B(n_758),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_770),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_795),
.B(n_804),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_753),
.A2(n_758),
.B1(n_761),
.B2(n_766),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_799),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_802),
.B(n_812),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_802),
.B(n_804),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_761),
.A2(n_878),
.B(n_835),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_878),
.A2(n_910),
.B(n_863),
.C(n_835),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_906),
.A2(n_868),
.B(n_862),
.C(n_880),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_775),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_903),
.A2(n_875),
.B1(n_815),
.B2(n_867),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_844),
.B(n_855),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_746),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_842),
.B(n_770),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_910),
.A2(n_834),
.B1(n_831),
.B2(n_814),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_801),
.A2(n_773),
.B(n_900),
.Y(n_1026)
);

NAND3xp33_ASAP7_75t_L g1027 ( 
.A(n_808),
.B(n_882),
.C(n_801),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_773),
.A2(n_900),
.B(n_899),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_867),
.A2(n_852),
.B1(n_847),
.B2(n_857),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_899),
.A2(n_847),
.B(n_842),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_844),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_847),
.A2(n_867),
.B(n_858),
.C(n_881),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_886),
.B(n_842),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_861),
.B(n_877),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_864),
.B(n_874),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_905),
.Y(n_1036)
);

INVx3_ASAP7_75t_SL g1037 ( 
.A(n_883),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_803),
.B(n_857),
.Y(n_1038)
);

OAI22x1_ASAP7_75t_L g1039 ( 
.A1(n_798),
.A2(n_907),
.B1(n_905),
.B2(n_852),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_803),
.B(n_770),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_786),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_786),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_786),
.B(n_792),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_907),
.A2(n_792),
.B1(n_809),
.B2(n_896),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_826),
.A2(n_798),
.B(n_866),
.C(n_809),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_792),
.B(n_896),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_792),
.A2(n_896),
.B(n_866),
.C(n_809),
.Y(n_1047)
);

OR2x6_ASAP7_75t_SL g1048 ( 
.A(n_896),
.B(n_457),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_817),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_926),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_950),
.B(n_922),
.Y(n_1051)
);

INVx6_ASAP7_75t_L g1052 ( 
.A(n_961),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_949),
.B(n_917),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_974),
.A2(n_970),
.B(n_952),
.Y(n_1054)
);

AOI31xp67_ASAP7_75t_L g1055 ( 
.A1(n_993),
.A2(n_912),
.A3(n_1029),
.B(n_1043),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_1033),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_955),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_1033),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_970),
.A2(n_979),
.B(n_915),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_SL g1061 ( 
.A1(n_969),
.A2(n_938),
.B(n_942),
.C(n_953),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_978),
.Y(n_1062)
);

OA22x2_ASAP7_75t_L g1063 ( 
.A1(n_990),
.A2(n_1037),
.B1(n_968),
.B2(n_929),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_920),
.B(n_918),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_956),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_938),
.A2(n_953),
.B1(n_931),
.B2(n_969),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_913),
.A2(n_921),
.B(n_976),
.Y(n_1067)
);

AO21x2_ASAP7_75t_L g1068 ( 
.A1(n_1005),
.A2(n_976),
.B(n_996),
.Y(n_1068)
);

AO21x2_ASAP7_75t_L g1069 ( 
.A1(n_1028),
.A2(n_954),
.B(n_1025),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1002),
.B(n_937),
.Y(n_1070)
);

AO31x2_ASAP7_75t_L g1071 ( 
.A1(n_1012),
.A2(n_1025),
.A3(n_1039),
.B(n_982),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_939),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1002),
.B(n_946),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_944),
.A2(n_1007),
.B(n_925),
.C(n_924),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_SL g1075 ( 
.A(n_964),
.B(n_1045),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1026),
.A2(n_1017),
.B(n_1009),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1004),
.A2(n_992),
.B(n_1027),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_948),
.B(n_1049),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_916),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_SL g1080 ( 
.A1(n_988),
.A2(n_942),
.B(n_943),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_928),
.A2(n_1018),
.B(n_933),
.Y(n_1081)
);

AO32x2_ASAP7_75t_L g1082 ( 
.A1(n_1012),
.A2(n_1041),
.A3(n_966),
.B1(n_935),
.B2(n_963),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_964),
.B(n_1021),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_980),
.B(n_1006),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1019),
.A2(n_1047),
.B(n_1030),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_973),
.B(n_975),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_951),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_951),
.B(n_973),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_SL g1089 ( 
.A1(n_958),
.A2(n_932),
.B(n_967),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_977),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_933),
.A2(n_983),
.B(n_936),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1032),
.A2(n_987),
.B(n_994),
.C(n_940),
.Y(n_1092)
);

NAND2x1_ASAP7_75t_L g1093 ( 
.A(n_983),
.B(n_1041),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1003),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_SL g1095 ( 
.A1(n_965),
.A2(n_1000),
.B(n_1024),
.C(n_962),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_941),
.Y(n_1096)
);

NOR2xp67_ASAP7_75t_L g1097 ( 
.A(n_1020),
.B(n_966),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_935),
.A2(n_999),
.B(n_997),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1014),
.A2(n_1016),
.B(n_1035),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_960),
.A2(n_1023),
.B1(n_1031),
.B2(n_1036),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1001),
.B(n_1011),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1022),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1044),
.A2(n_1038),
.B(n_1046),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1034),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_919),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_934),
.A2(n_1040),
.B(n_978),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_972),
.B(n_1015),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1008),
.A2(n_1042),
.B(n_1010),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_984),
.A2(n_985),
.B(n_1042),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_984),
.A2(n_985),
.B1(n_951),
.B2(n_927),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1013),
.B(n_995),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_991),
.A2(n_1042),
.B(n_1010),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_991),
.A2(n_1010),
.B(n_951),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_991),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_927),
.B(n_957),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_971),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_927),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_957),
.B(n_961),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_SL g1119 ( 
.A1(n_957),
.A2(n_945),
.B(n_981),
.Y(n_1119)
);

AO21x1_ASAP7_75t_L g1120 ( 
.A1(n_930),
.A2(n_739),
.B(n_895),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_986),
.A2(n_952),
.B(n_970),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_912),
.A2(n_608),
.B(n_959),
.C(n_949),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_914),
.B(n_785),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_979),
.A2(n_974),
.B(n_913),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_973),
.B(n_755),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_979),
.A2(n_974),
.B(n_913),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_974),
.A2(n_741),
.B(n_757),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_986),
.A2(n_952),
.B(n_976),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_914),
.B(n_785),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_974),
.A2(n_741),
.B(n_757),
.Y(n_1131)
);

BUFx8_ASAP7_75t_SL g1132 ( 
.A(n_989),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_951),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_947),
.B(n_560),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_996),
.A2(n_841),
.A3(n_986),
.B(n_1012),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_SL g1138 ( 
.A1(n_949),
.A2(n_734),
.B(n_781),
.Y(n_1138)
);

AO22x2_ASAP7_75t_L g1139 ( 
.A1(n_1025),
.A2(n_739),
.B1(n_969),
.B2(n_938),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_916),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_961),
.Y(n_1141)
);

BUFx4_ASAP7_75t_SL g1142 ( 
.A(n_989),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_979),
.A2(n_974),
.B(n_913),
.Y(n_1143)
);

AO21x1_ASAP7_75t_L g1144 ( 
.A1(n_930),
.A2(n_739),
.B(n_895),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_914),
.B(n_785),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_950),
.B(n_757),
.Y(n_1146)
);

CKINVDCx11_ASAP7_75t_R g1147 ( 
.A(n_1048),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_914),
.A2(n_781),
.B1(n_757),
.B2(n_741),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_947),
.B(n_626),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_974),
.A2(n_741),
.B(n_749),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_SL g1151 ( 
.A1(n_949),
.A2(n_734),
.B(n_781),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_923),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_974),
.A2(n_741),
.B(n_757),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_914),
.A2(n_781),
.B1(n_757),
.B2(n_741),
.Y(n_1159)
);

INVx3_ASAP7_75t_SL g1160 ( 
.A(n_971),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_SL g1161 ( 
.A1(n_912),
.A2(n_741),
.B(n_749),
.C(n_913),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_947),
.B(n_560),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_974),
.A2(n_741),
.B(n_757),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_950),
.B(n_757),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_914),
.B(n_785),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_R g1168 ( 
.A(n_945),
.B(n_457),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_926),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_912),
.A2(n_608),
.B(n_959),
.C(n_949),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_996),
.A2(n_841),
.A3(n_986),
.B(n_1012),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_947),
.B(n_560),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_996),
.A2(n_841),
.A3(n_986),
.B(n_1012),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1005),
.A2(n_998),
.B(n_986),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_912),
.A2(n_608),
.B(n_959),
.C(n_949),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_973),
.B(n_755),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_950),
.B(n_757),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_930),
.B(n_608),
.C(n_614),
.Y(n_1179)
);

OAI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_990),
.A2(n_620),
.B1(n_556),
.B2(n_560),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_923),
.Y(n_1181)
);

NAND2x1_ASAP7_75t_L g1182 ( 
.A(n_983),
.B(n_809),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_961),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1064),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1135),
.A2(n_1153),
.B(n_1152),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1136),
.B(n_1162),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1057),
.B(n_1059),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1154),
.A2(n_1156),
.B(n_1155),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1087),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1050),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1094),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1171),
.A2(n_1176),
.B(n_1150),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1066),
.A2(n_1120),
.A3(n_1144),
.B(n_1074),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1161),
.A2(n_1066),
.B(n_1173),
.C(n_1080),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1086),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1163),
.A2(n_1175),
.B(n_1170),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_1132),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1089),
.B(n_1058),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1086),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1139),
.A2(n_1159),
.B1(n_1148),
.B2(n_1063),
.Y(n_1201)
);

BUFx4f_ASAP7_75t_L g1202 ( 
.A(n_1052),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1166),
.A2(n_1067),
.B(n_1121),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1079),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1099),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1057),
.B(n_1059),
.Y(n_1206)
);

CKINVDCx11_ASAP7_75t_R g1207 ( 
.A(n_1160),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1087),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1140),
.B(n_1096),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1072),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1119),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1076),
.A2(n_1060),
.B(n_1091),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1054),
.A2(n_1085),
.B(n_1081),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1133),
.Y(n_1214)
);

CKINVDCx16_ASAP7_75t_R g1215 ( 
.A(n_1168),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1077),
.A2(n_1143),
.B(n_1127),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1150),
.A2(n_1164),
.B(n_1158),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1169),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1128),
.A2(n_1131),
.B(n_1053),
.C(n_1125),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1068),
.Y(n_1220)
);

AND2x2_ASAP7_75t_SL g1221 ( 
.A(n_1075),
.B(n_1139),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_1133),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_SL g1223 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1143),
.Y(n_1223)
);

AO21x2_ASAP7_75t_L g1224 ( 
.A1(n_1077),
.A2(n_1069),
.B(n_1092),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1061),
.A2(n_1129),
.B(n_1106),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1157),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1181),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1139),
.A2(n_1063),
.B1(n_1180),
.B2(n_1146),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1051),
.B(n_1178),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1107),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1069),
.Y(n_1231)
);

AO21x2_ASAP7_75t_L g1232 ( 
.A1(n_1106),
.A2(n_1083),
.B(n_1073),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1146),
.A2(n_1178),
.B(n_1165),
.C(n_1105),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1129),
.A2(n_1103),
.B(n_1108),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1147),
.Y(n_1235)
);

INVxp67_ASAP7_75t_SL g1236 ( 
.A(n_1101),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1078),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1126),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1138),
.A2(n_1151),
.B(n_1165),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1104),
.A2(n_1101),
.B(n_1065),
.C(n_1102),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1078),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1142),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1070),
.A2(n_1073),
.B(n_1084),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_SL g1244 ( 
.A1(n_1182),
.A2(n_1093),
.B(n_1130),
.C(n_1167),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1124),
.A2(n_1145),
.B1(n_1084),
.B2(n_1100),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1062),
.B(n_1177),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1052),
.A2(n_1068),
.B1(n_1183),
.B2(n_1141),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1137),
.Y(n_1248)
);

AOI22x1_ASAP7_75t_L g1249 ( 
.A1(n_1116),
.A2(n_1113),
.B1(n_1112),
.B2(n_1109),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1114),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1118),
.A2(n_1095),
.B(n_1110),
.C(n_1088),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1113),
.A2(n_1110),
.B(n_1115),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1062),
.A2(n_1115),
.B(n_1117),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1111),
.A2(n_1116),
.B1(n_1097),
.B2(n_1082),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1082),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1137),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1082),
.B(n_1071),
.Y(n_1257)
);

INVx4_ASAP7_75t_L g1258 ( 
.A(n_1055),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1137),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1174),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1071),
.Y(n_1261)
);

INVx5_ASAP7_75t_L g1262 ( 
.A(n_1071),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1172),
.B(n_1174),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1172),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1174),
.A2(n_1179),
.B(n_608),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1168),
.Y(n_1266)
);

NAND2xp33_ASAP7_75t_SL g1267 ( 
.A(n_1066),
.B(n_781),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1179),
.A2(n_608),
.B(n_1122),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1087),
.Y(n_1271)
);

OA21x2_ASAP7_75t_L g1272 ( 
.A1(n_1067),
.A2(n_1054),
.B(n_1081),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1050),
.Y(n_1273)
);

BUFx2_ASAP7_75t_R g1274 ( 
.A(n_1132),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1148),
.B(n_1159),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1149),
.A2(n_623),
.B1(n_914),
.B2(n_626),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_1101),
.Y(n_1278)
);

BUFx2_ASAP7_75t_R g1279 ( 
.A(n_1132),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1050),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1090),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1090),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_1079),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1057),
.B(n_1059),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_SL g1286 ( 
.A(n_1052),
.B(n_457),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1168),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1168),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_1116),
.B(n_958),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1111),
.Y(n_1292)
);

AND2x6_ASAP7_75t_L g1293 ( 
.A(n_1053),
.B(n_1021),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1294)
);

AOI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1150),
.A2(n_1098),
.B(n_1121),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1068),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1056),
.A2(n_1134),
.B(n_1123),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1136),
.A2(n_1162),
.B1(n_1173),
.B2(n_560),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1087),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1067),
.A2(n_1054),
.B(n_1081),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1218),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1236),
.B(n_1278),
.Y(n_1303)
);

BUFx4f_ASAP7_75t_SL g1304 ( 
.A(n_1198),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1207),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1220),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_SL g1307 ( 
.A1(n_1209),
.A2(n_1263),
.B(n_1185),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1239),
.B(n_1275),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1192),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1220),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1233),
.A2(n_1195),
.B(n_1269),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1187),
.A2(n_1299),
.B1(n_1201),
.B2(n_1275),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1212),
.A2(n_1203),
.B(n_1217),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1220),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_SL g1315 ( 
.A1(n_1265),
.A2(n_1193),
.B(n_1286),
.C(n_1271),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1229),
.B(n_1240),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1240),
.B(n_1216),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1199),
.B(n_1191),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1184),
.A2(n_1290),
.B(n_1186),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1202),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1216),
.B(n_1284),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1267),
.A2(n_1219),
.B(n_1223),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1251),
.A2(n_1216),
.B(n_1219),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1204),
.B(n_1238),
.Y(n_1324)
);

OA22x2_ASAP7_75t_L g1325 ( 
.A1(n_1255),
.A2(n_1266),
.B1(n_1287),
.B2(n_1288),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1238),
.B(n_1188),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1198),
.Y(n_1327)
);

AOI31xp33_ASAP7_75t_L g1328 ( 
.A1(n_1201),
.A2(n_1228),
.A3(n_1254),
.B(n_1288),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1189),
.A2(n_1291),
.B(n_1281),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1273),
.B(n_1280),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1277),
.A2(n_1221),
.B1(n_1245),
.B2(n_1254),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1202),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1247),
.B(n_1206),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1243),
.B(n_1250),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1293),
.B(n_1245),
.Y(n_1335)
);

BUFx12f_ASAP7_75t_L g1336 ( 
.A(n_1207),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_SL g1337 ( 
.A1(n_1211),
.A2(n_1266),
.B(n_1287),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1230),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1244),
.A2(n_1224),
.B(n_1301),
.C(n_1272),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1243),
.A2(n_1232),
.B(n_1224),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1296),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1221),
.A2(n_1215),
.B1(n_1247),
.B2(n_1289),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_R g1343 ( 
.A(n_1235),
.B(n_1200),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1243),
.A2(n_1232),
.B(n_1196),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1213),
.A2(n_1257),
.B(n_1261),
.C(n_1262),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1197),
.A2(n_1270),
.B(n_1268),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1262),
.A2(n_1264),
.B(n_1225),
.C(n_1252),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1196),
.A2(n_1200),
.B(n_1301),
.Y(n_1349)
);

OA22x2_ASAP7_75t_L g1350 ( 
.A1(n_1246),
.A2(n_1253),
.B1(n_1237),
.B2(n_1242),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1241),
.B(n_1194),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1241),
.B(n_1194),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1293),
.B(n_1227),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1235),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1285),
.A2(n_1190),
.B1(n_1222),
.B2(n_1262),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1274),
.Y(n_1356)
);

OA22x2_ASAP7_75t_L g1357 ( 
.A1(n_1258),
.A2(n_1259),
.B1(n_1260),
.B2(n_1256),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1222),
.A2(n_1262),
.B1(n_1271),
.B2(n_1208),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1214),
.B(n_1194),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1279),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1214),
.B(n_1222),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1296),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1300),
.B(n_1226),
.Y(n_1363)
);

OA22x2_ASAP7_75t_L g1364 ( 
.A1(n_1258),
.A2(n_1260),
.B1(n_1259),
.B2(n_1256),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1249),
.A2(n_1276),
.B(n_1298),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1210),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1268),
.A2(n_1291),
.B(n_1297),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1234),
.B(n_1248),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1295),
.A2(n_1205),
.B1(n_1231),
.B2(n_1292),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1294),
.B(n_1297),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1292),
.B(n_1294),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1292),
.A2(n_1212),
.B(n_1203),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_SL g1373 ( 
.A1(n_1233),
.A2(n_1066),
.B(n_1122),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1212),
.A2(n_1203),
.B(n_1217),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1216),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1334),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1309),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1340),
.A2(n_1348),
.B(n_1317),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1344),
.B(n_1350),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1371),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1373),
.A2(n_1311),
.B(n_1322),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1372),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1348),
.A2(n_1375),
.B(n_1345),
.Y(n_1383)
);

AO21x1_ASAP7_75t_SL g1384 ( 
.A1(n_1335),
.A2(n_1321),
.B(n_1310),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1303),
.B(n_1375),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1350),
.B(n_1349),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1359),
.B(n_1368),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1345),
.A2(n_1339),
.B(n_1331),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1372),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1369),
.A2(n_1328),
.B(n_1353),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1308),
.B(n_1370),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1351),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1302),
.B(n_1352),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1330),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1372),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1308),
.B(n_1313),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1346),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1338),
.Y(n_1398)
);

AO21x1_ASAP7_75t_SL g1399 ( 
.A1(n_1306),
.A2(n_1341),
.B(n_1314),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1316),
.B(n_1308),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1357),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1312),
.A2(n_1342),
.B1(n_1325),
.B2(n_1333),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1323),
.B(n_1325),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1310),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1313),
.B(n_1374),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_1314),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1355),
.A2(n_1358),
.B(n_1320),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1318),
.B(n_1362),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1313),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1324),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1357),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1374),
.B(n_1319),
.Y(n_1412)
);

NOR2x1_ASAP7_75t_R g1413 ( 
.A(n_1327),
.B(n_1336),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1315),
.A2(n_1363),
.B(n_1366),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1364),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1361),
.B(n_1363),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1364),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1381),
.A2(n_1356),
.B1(n_1343),
.B2(n_1320),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1385),
.B(n_1329),
.Y(n_1419)
);

OR2x2_ASAP7_75t_SL g1420 ( 
.A(n_1383),
.B(n_1307),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1404),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1387),
.B(n_1396),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1376),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1381),
.B(n_1326),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1377),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1377),
.Y(n_1426)
);

AO21x2_ASAP7_75t_L g1427 ( 
.A1(n_1388),
.A2(n_1367),
.B(n_1365),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1384),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1396),
.B(n_1347),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1384),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1414),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1404),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1412),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1412),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1406),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1405),
.B(n_1391),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1389),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1405),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1406),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1398),
.B(n_1337),
.Y(n_1440)
);

AOI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1419),
.A2(n_1402),
.B1(n_1403),
.B2(n_1389),
.C(n_1388),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1435),
.B(n_1398),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1421),
.B(n_1408),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1428),
.B(n_1430),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1428),
.B(n_1391),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1424),
.A2(n_1402),
.B1(n_1388),
.B2(n_1403),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1422),
.B(n_1391),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1427),
.A2(n_1378),
.B(n_1388),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1430),
.B(n_1386),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1425),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1431),
.B(n_1400),
.C(n_1393),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1431),
.A2(n_1390),
.B1(n_1417),
.B2(n_1415),
.Y(n_1452)
);

OAI321xp33_ASAP7_75t_L g1453 ( 
.A1(n_1418),
.A2(n_1379),
.A3(n_1386),
.B1(n_1411),
.B2(n_1415),
.C(n_1417),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1422),
.B(n_1399),
.Y(n_1454)
);

CKINVDCx16_ASAP7_75t_R g1455 ( 
.A(n_1440),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1425),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1425),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1422),
.B(n_1399),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1424),
.A2(n_1386),
.B1(n_1379),
.B2(n_1383),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1420),
.A2(n_1407),
.B1(n_1380),
.B2(n_1386),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1426),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1431),
.A2(n_1390),
.B1(n_1411),
.B2(n_1401),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1427),
.A2(n_1378),
.B(n_1409),
.Y(n_1463)
);

AOI222xp33_ASAP7_75t_L g1464 ( 
.A1(n_1429),
.A2(n_1401),
.B1(n_1395),
.B2(n_1382),
.C1(n_1397),
.C2(n_1392),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1418),
.A2(n_1390),
.B1(n_1378),
.B2(n_1383),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1408),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1436),
.B(n_1380),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1436),
.B(n_1410),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1420),
.A2(n_1379),
.B1(n_1394),
.B2(n_1416),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1432),
.B(n_1393),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1437),
.A2(n_1383),
.B1(n_1382),
.B2(n_1395),
.Y(n_1471)
);

INVx4_ASAP7_75t_SL g1472 ( 
.A(n_1449),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1442),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1446),
.A2(n_1439),
.B(n_1435),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1448),
.B(n_1437),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1450),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1450),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1456),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1471),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1456),
.B(n_1423),
.Y(n_1480)
);

INVxp67_ASAP7_75t_SL g1481 ( 
.A(n_1446),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1465),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1457),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1457),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1448),
.B(n_1433),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1463),
.Y(n_1486)
);

OA21x2_ASAP7_75t_L g1487 ( 
.A1(n_1441),
.A2(n_1419),
.B(n_1434),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1463),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1461),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1444),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1454),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1455),
.B(n_1413),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_SL g1493 ( 
.A1(n_1460),
.A2(n_1439),
.B(n_1433),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1454),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1470),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1474),
.B(n_1491),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1486),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1476),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1474),
.B(n_1458),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1476),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1479),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1491),
.B(n_1458),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1495),
.B(n_1479),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1472),
.B(n_1449),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1491),
.B(n_1494),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_SL g1506 ( 
.A(n_1493),
.B(n_1354),
.C(n_1464),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1481),
.B(n_1451),
.C(n_1452),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1477),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1490),
.B(n_1447),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1473),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1473),
.B(n_1443),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1490),
.B(n_1447),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1477),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1478),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1492),
.B(n_1444),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1481),
.B(n_1438),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1486),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1493),
.B(n_1433),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1487),
.B(n_1433),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1487),
.B(n_1467),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1487),
.B(n_1467),
.Y(n_1521)
);

OAI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1482),
.A2(n_1453),
.B1(n_1459),
.B2(n_1379),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1486),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1480),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1472),
.B(n_1445),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1488),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1480),
.B(n_1443),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1483),
.B(n_1470),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1515),
.B(n_1445),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1482),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1501),
.B(n_1503),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1514),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1514),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1519),
.Y(n_1534)
);

AOI211xp5_ASAP7_75t_L g1535 ( 
.A1(n_1506),
.A2(n_1475),
.B(n_1485),
.C(n_1469),
.Y(n_1535)
);

OAI21xp33_ASAP7_75t_L g1536 ( 
.A1(n_1503),
.A2(n_1485),
.B(n_1475),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1515),
.B(n_1445),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1511),
.B(n_1466),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1510),
.B(n_1487),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1525),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1498),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1511),
.B(n_1483),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1525),
.B(n_1475),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1525),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1498),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1500),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1527),
.B(n_1484),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1527),
.B(n_1484),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1509),
.B(n_1468),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1525),
.B(n_1472),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1509),
.B(n_1468),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1528),
.B(n_1524),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1519),
.Y(n_1553)
);

NAND2x1_ASAP7_75t_L g1554 ( 
.A(n_1525),
.B(n_1485),
.Y(n_1554)
);

NAND2x2_ASAP7_75t_L g1555 ( 
.A(n_1506),
.B(n_1332),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1520),
.B(n_1487),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1528),
.B(n_1489),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1500),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1508),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1509),
.B(n_1489),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1519),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1508),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1505),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1512),
.B(n_1502),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1564),
.B(n_1520),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1564),
.B(n_1520),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1556),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1529),
.B(n_1521),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1541),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1531),
.Y(n_1570)
);

NOR2xp67_ASAP7_75t_L g1571 ( 
.A(n_1563),
.B(n_1496),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1531),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1550),
.B(n_1505),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1530),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1534),
.Y(n_1575)
);

NAND2xp33_ASAP7_75t_L g1576 ( 
.A(n_1529),
.B(n_1360),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1544),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1545),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1546),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1540),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1537),
.B(n_1521),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1540),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1558),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1560),
.B(n_1513),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1534),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1532),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1563),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1537),
.B(n_1496),
.Y(n_1588)
);

AOI222xp33_ASAP7_75t_L g1589 ( 
.A1(n_1539),
.A2(n_1507),
.B1(n_1516),
.B2(n_1522),
.C1(n_1496),
.C2(n_1462),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1555),
.A2(n_1507),
.B1(n_1499),
.B2(n_1504),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1586),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1586),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1571),
.A2(n_1535),
.B(n_1536),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1572),
.B(n_1533),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_L g1595 ( 
.A1(n_1590),
.A2(n_1552),
.B(n_1505),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1572),
.B(n_1560),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1587),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1569),
.Y(n_1598)
);

OAI31xp33_ASAP7_75t_L g1599 ( 
.A1(n_1574),
.A2(n_1516),
.A3(n_1543),
.B(n_1553),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_L g1600 ( 
.A(n_1589),
.B(n_1552),
.C(n_1559),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1588),
.B(n_1573),
.Y(n_1601)
);

AOI21xp33_ASAP7_75t_L g1602 ( 
.A1(n_1589),
.A2(n_1542),
.B(n_1562),
.Y(n_1602)
);

OAI211xp5_ASAP7_75t_L g1603 ( 
.A1(n_1574),
.A2(n_1543),
.B(n_1554),
.C(n_1561),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1588),
.B(n_1549),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1549),
.Y(n_1605)
);

OAI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1567),
.A2(n_1555),
.B1(n_1561),
.B2(n_1553),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1570),
.A2(n_1499),
.B(n_1550),
.Y(n_1607)
);

AOI32xp33_ASAP7_75t_L g1608 ( 
.A1(n_1565),
.A2(n_1499),
.A3(n_1475),
.B1(n_1518),
.B2(n_1485),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1570),
.B(n_1551),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1569),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1602),
.B(n_1577),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1604),
.B(n_1588),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1601),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1605),
.B(n_1573),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1609),
.B(n_1580),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1591),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1607),
.B(n_1573),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1592),
.B(n_1304),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1596),
.B(n_1580),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1597),
.B(n_1582),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_R g1621 ( 
.A(n_1594),
.B(n_1573),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1611),
.A2(n_1600),
.B1(n_1593),
.B2(n_1567),
.C(n_1599),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1611),
.A2(n_1571),
.B1(n_1603),
.B2(n_1607),
.Y(n_1623)
);

OAI21xp33_ASAP7_75t_L g1624 ( 
.A1(n_1618),
.A2(n_1595),
.B(n_1608),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1617),
.A2(n_1603),
.B(n_1567),
.Y(n_1625)
);

AND2x2_ASAP7_75t_SL g1626 ( 
.A(n_1619),
.B(n_1576),
.Y(n_1626)
);

AOI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1615),
.A2(n_1610),
.B1(n_1598),
.B2(n_1606),
.C(n_1565),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_L g1628 ( 
.A(n_1620),
.B(n_1582),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1612),
.A2(n_1577),
.B(n_1566),
.Y(n_1629)
);

OAI211xp5_ASAP7_75t_L g1630 ( 
.A1(n_1613),
.A2(n_1578),
.B(n_1583),
.C(n_1579),
.Y(n_1630)
);

AOI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1616),
.A2(n_1566),
.B1(n_1565),
.B2(n_1578),
.C(n_1579),
.Y(n_1631)
);

OAI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1622),
.A2(n_1618),
.B1(n_1585),
.B2(n_1575),
.C(n_1566),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1629),
.Y(n_1633)
);

NAND4xp25_ASAP7_75t_L g1634 ( 
.A(n_1625),
.B(n_1614),
.C(n_1573),
.D(n_1621),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1623),
.A2(n_1585),
.B(n_1575),
.C(n_1583),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1626),
.B(n_1568),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1627),
.A2(n_1585),
.B1(n_1575),
.B2(n_1581),
.C(n_1568),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1624),
.A2(n_1581),
.B1(n_1568),
.B2(n_1550),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1634),
.B(n_1628),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1636),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1633),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1638),
.B(n_1631),
.Y(n_1642)
);

NOR2xp67_ASAP7_75t_SL g1643 ( 
.A(n_1632),
.B(n_1305),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1635),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1637),
.B(n_1630),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1640),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1641),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_R g1648 ( 
.A(n_1639),
.B(n_1327),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1644),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1639),
.B(n_1584),
.Y(n_1650)
);

NOR2x1_ASAP7_75t_L g1651 ( 
.A(n_1646),
.B(n_1645),
.Y(n_1651)
);

NOR3xp33_ASAP7_75t_SL g1652 ( 
.A(n_1648),
.B(n_1642),
.C(n_1643),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1650),
.A2(n_1647),
.B(n_1649),
.Y(n_1653)
);

AOI31xp33_ASAP7_75t_L g1654 ( 
.A1(n_1653),
.A2(n_1581),
.A3(n_1584),
.B(n_1304),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1654),
.B(n_1651),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1655),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1655),
.Y(n_1657)
);

AOI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1652),
.B(n_1542),
.Y(n_1658)
);

OAI31xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1656),
.A2(n_1499),
.A3(n_1518),
.B(n_1551),
.Y(n_1659)
);

AO22x2_ASAP7_75t_L g1660 ( 
.A1(n_1658),
.A2(n_1548),
.B1(n_1547),
.B2(n_1557),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1659),
.B(n_1512),
.Y(n_1661)
);

OAI22x1_ASAP7_75t_L g1662 ( 
.A1(n_1661),
.A2(n_1499),
.B1(n_1548),
.B2(n_1547),
.Y(n_1662)
);

OAI22xp33_ASAP7_75t_SL g1663 ( 
.A1(n_1660),
.A2(n_1526),
.B1(n_1523),
.B2(n_1497),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1663),
.A2(n_1557),
.B(n_1538),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1664),
.B(n_1662),
.C(n_1517),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1517),
.B(n_1497),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1666),
.A2(n_1526),
.B1(n_1523),
.B2(n_1517),
.Y(n_1667)
);

AOI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1526),
.B(n_1523),
.C(n_1497),
.Y(n_1668)
);


endmodule