module real_jpeg_2469_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_23),
.B1(n_37),
.B2(n_45),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_28),
.B1(n_37),
.B2(n_49),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_37),
.B1(n_60),
.B2(n_61),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_27),
.C(n_28),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_23),
.B1(n_39),
.B2(n_45),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_3),
.A2(n_28),
.B1(n_39),
.B2(n_49),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_3),
.A2(n_39),
.B1(n_60),
.B2(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_3),
.B(n_48),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_3),
.B(n_57),
.C(n_61),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_3),
.B(n_35),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_75),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_34),
.C(n_76),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_3),
.B(n_63),
.Y(n_170)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_84),
.Y(n_203)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_10),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_127),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_209),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_188),
.B(n_208),
.Y(n_14)
);

OAI211xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_107),
.B(n_130),
.C(n_187),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_17),
.B(n_96),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_67),
.B2(n_68),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_18),
.B(n_70),
.C(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_40),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_20),
.B(n_42),
.C(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_21),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_45),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_28),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_28),
.B(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_30),
.A2(n_31),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_31),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_31),
.B(n_158),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_31),
.B(n_129),
.C(n_170),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_32),
.B(n_38),
.Y(n_86)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_33),
.A2(n_34),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_34),
.B(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_38),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_52),
.B2(n_66),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_41),
.A2(n_42),
.B1(n_89),
.B2(n_100),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_41),
.B(n_89),
.C(n_194),
.Y(n_231)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_44),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_46),
.B(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_46),
.Y(n_223)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_51),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_104),
.C(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_52),
.A2(n_66),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_52),
.A2(n_227),
.B(n_230),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_52),
.B(n_227),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_52)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_63),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_65),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_55),
.A2(n_59),
.B(n_65),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

AOI22x1_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_61),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_61),
.B(n_163),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_87),
.B2(n_88),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_81),
.B2(n_82),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_82),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_71),
.A2(n_72),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_71),
.B(n_164),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_71),
.A2(n_72),
.B1(n_89),
.B2(n_100),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_71),
.B(n_89),
.C(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_74),
.B(n_79),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_73),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_74),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_75),
.A2(n_206),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_79),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_85),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_86),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_85),
.B(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.C(n_92),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_91),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_93),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_93),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_92),
.B(n_115),
.C(n_120),
.Y(n_191)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_94),
.B(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.C(n_103),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_103),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_105),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_131),
.C(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_109),
.B(n_110),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_111),
.B(n_113),
.C(n_122),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_121),
.B2(n_122),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_124),
.B(n_128),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_126),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_129),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_128),
.A2(n_129),
.B1(n_142),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_137),
.C(n_142),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_149),
.B(n_186),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_136),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_161),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_180),
.B(n_185),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_174),
.B(n_179),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_166),
.B(n_173),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_160),
.B(n_165),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_157),
.B(n_159),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_162),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_172),
.Y(n_173)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_176),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_184),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_190),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_193),
.C(n_198),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_207),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_202),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_207),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_232),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_213),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_231),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_225),
.B2(n_226),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);


endmodule