module fake_jpeg_1712_n_213 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_213);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_4),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_23),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_82),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_51),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_51),
.B1(n_60),
.B2(n_53),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_80),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_94),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_66),
.B1(n_65),
.B2(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_74),
.B1(n_62),
.B2(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_63),
.B1(n_52),
.B2(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_68),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_104),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_57),
.B1(n_76),
.B2(n_50),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_77),
.B(n_72),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_105),
.Y(n_120)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_61),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_65),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_110),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_0),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_31),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_115),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_2),
.C(n_3),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_5),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_2),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_7),
.Y(n_145)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_135),
.B1(n_113),
.B2(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_70),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_58),
.C(n_55),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_101),
.A2(n_70),
.B1(n_71),
.B2(n_58),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_3),
.CI(n_4),
.CON(n_136),
.SN(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_5),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_150),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_142),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_154),
.B1(n_155),
.B2(n_158),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_6),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_34),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_7),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_145),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_8),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_9),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_55),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_33),
.C(n_41),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_32),
.B1(n_47),
.B2(n_45),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_29),
.B1(n_44),
.B2(n_43),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_137),
.B(n_10),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_124),
.B(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_13),
.B(n_14),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_157),
.B(n_155),
.Y(n_166)
);

XOR2x1_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_136),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_169),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_133),
.B(n_15),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_13),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_15),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_151),
.Y(n_179)
);

AO221x1_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_181),
.B1(n_154),
.B2(n_17),
.C(n_16),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_182),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_143),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_188),
.Y(n_203)
);

AO221x1_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_174),
.B1(n_171),
.B2(n_175),
.C(n_164),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_198),
.B1(n_186),
.B2(n_183),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_166),
.B(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_197),
.C(n_180),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_178),
.C(n_165),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_172),
.B(n_146),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_188),
.C(n_190),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_203),
.B1(n_192),
.B2(n_170),
.Y(n_206)
);

OAI31xp33_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_163),
.A3(n_177),
.B(n_194),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_16),
.C(n_19),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_199),
.Y(n_207)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_208),
.B(n_206),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_204),
.C(n_24),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_210),
.Y(n_211)
);

OAI221xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_20),
.B1(n_30),
.B2(n_35),
.C(n_36),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_212),
.B(n_39),
.Y(n_213)
);


endmodule