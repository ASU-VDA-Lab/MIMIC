module fake_jpeg_4062_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_17),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_16),
.B1(n_26),
.B2(n_28),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx9p33_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_2),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_32),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_16),
.B1(n_25),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_50),
.B1(n_57),
.B2(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_18),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_33),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_33),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_16),
.B1(n_21),
.B2(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_63),
.Y(n_95)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_64),
.B(n_67),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_41),
.B1(n_25),
.B2(n_29),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_69),
.A2(n_35),
.B1(n_34),
.B2(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_73),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_19),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_79),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_41),
.B1(n_31),
.B2(n_22),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_18),
.B1(n_22),
.B2(n_34),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_51),
.A2(n_30),
.B1(n_17),
.B2(n_27),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_82),
.A2(n_92),
.B1(n_15),
.B2(n_6),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_24),
.B1(n_35),
.B2(n_4),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_84),
.B(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_90),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_23),
.B1(n_20),
.B2(n_24),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_2),
.B(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_5),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_53),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_97),
.B1(n_110),
.B2(n_81),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_35),
.B1(n_34),
.B2(n_38),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_20),
.B(n_24),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_102),
.B(n_106),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_35),
.B(n_34),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_109),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_63),
.B1(n_68),
.B2(n_90),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_24),
.B(n_3),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_106),
.B1(n_102),
.B2(n_120),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_64),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_119),
.B1(n_75),
.B2(n_73),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_5),
.B(n_7),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_67),
.B(n_62),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_67),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_124),
.B1(n_129),
.B2(n_110),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_127),
.B1(n_111),
.B2(n_115),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_86),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_130),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_86),
.B1(n_84),
.B2(n_59),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_125),
.A2(n_98),
.B1(n_99),
.B2(n_114),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_59),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_113),
.B1(n_118),
.B2(n_109),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_59),
.Y(n_133)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_62),
.C(n_64),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_99),
.C(n_117),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_142),
.B(n_149),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_97),
.B(n_62),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_139),
.B(n_141),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_96),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_95),
.Y(n_144)
);

CKINVDCx11_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_108),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_105),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_94),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_78),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_162),
.B1(n_169),
.B2(n_149),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_170),
.C(n_136),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_161),
.Y(n_182)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

OR2x6_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_117),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_138),
.B(n_137),
.Y(n_190)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_167),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_106),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_125),
.Y(n_191)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_116),
.B1(n_105),
.B2(n_119),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_173),
.Y(n_198)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_175),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_178),
.B(n_110),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_181),
.A2(n_187),
.B1(n_197),
.B2(n_200),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_128),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_193),
.Y(n_217)
);

XOR2x2_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_166),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_191),
.Y(n_207)
);

AO22x2_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_135),
.B1(n_127),
.B2(n_129),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_189),
.B(n_190),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_135),
.B(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_194),
.B(n_196),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_201),
.C(n_158),
.Y(n_218)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_121),
.B1(n_142),
.B2(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_199),
.B(n_175),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_140),
.B(n_145),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_136),
.C(n_126),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_221),
.Y(n_231)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_178),
.B1(n_162),
.B2(n_152),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_189),
.B1(n_197),
.B2(n_179),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_174),
.B1(n_151),
.B2(n_163),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_164),
.B1(n_171),
.B2(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_167),
.B1(n_152),
.B2(n_159),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_153),
.B1(n_150),
.B2(n_134),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_195),
.C(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_194),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_153),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_220),
.A2(n_200),
.B(n_187),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_182),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_208),
.C(n_132),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_225),
.C(n_205),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_183),
.C(n_190),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_228),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_234),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_210),
.A2(n_193),
.B1(n_184),
.B2(n_202),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_232),
.A2(n_235),
.B1(n_203),
.B2(n_220),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_176),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_134),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_216),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_202),
.B1(n_180),
.B2(n_141),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_208),
.B1(n_211),
.B2(n_209),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_240),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_244),
.C(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_225),
.C(n_224),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_100),
.B(n_10),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_204),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_100),
.C(n_10),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_205),
.C(n_207),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_233),
.C(n_222),
.Y(n_253)
);

OAI321xp33_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_227),
.A3(n_233),
.B1(n_237),
.B2(n_226),
.C(n_220),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_253),
.B(n_255),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_156),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_SL g255 ( 
.A1(n_249),
.A2(n_231),
.B(n_176),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_156),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_242),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_9),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_9),
.Y(n_261)
);

AOI221xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_263),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_248),
.B1(n_241),
.B2(n_78),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_266),
.B(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_270),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_260),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_250),
.B(n_241),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_250),
.C(n_14),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_272),
.A2(n_273),
.B(n_101),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_269),
.C(n_101),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_277),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_276),
.B(n_72),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_66),
.Y(n_280)
);


endmodule