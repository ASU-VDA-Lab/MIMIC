module fake_jpeg_282_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_0),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_38),
.B1(n_37),
.B2(n_45),
.Y(n_56)
);

AO21x2_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_4),
.B(n_6),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_47),
.B1(n_45),
.B2(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_46),
.B1(n_2),
.B2(n_3),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_43),
.B1(n_40),
.B2(n_35),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_47),
.B1(n_40),
.B2(n_35),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_50),
.Y(n_59)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_67),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_48),
.B(n_36),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_14),
.Y(n_68)
);

AOI32xp33_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_73),
.A3(n_61),
.B1(n_59),
.B2(n_27),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_71),
.B(n_76),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_6),
.Y(n_89)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_16),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_62),
.B(n_8),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_55),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_88),
.C(n_62),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_60),
.C(n_62),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_7),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_100),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_18),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_97),
.C(n_102),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_20),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_103),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_15),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_7),
.B(n_9),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_9),
.B(n_10),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_30),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_21),
.C(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_78),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_11),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_11),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_12),
.Y(n_111)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_13),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_112),
.C(n_114),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_22),
.B(n_24),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_29),
.B1(n_94),
.B2(n_112),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_95),
.C(n_97),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_109),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_109),
.C(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_125),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_108),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_126),
.B(n_123),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_117),
.C(n_116),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_104),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_116),
.Y(n_132)
);


endmodule