module fake_jpeg_20409_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_SL g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_17),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_17),
.B1(n_15),
.B2(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_10),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_23),
.B(n_13),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_19),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_14),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_29),
.B1(n_21),
.B2(n_22),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_50),
.B1(n_35),
.B2(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_51),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_12),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_57),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_42),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_55),
.B(n_44),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_38),
.B(n_42),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_36),
.B1(n_27),
.B2(n_40),
.Y(n_56)
);

INVxp67_ASAP7_75t_SL g60 ( 
.A(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_9),
.Y(n_57)
);

AOI221xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_51),
.B1(n_49),
.B2(n_46),
.C(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_62),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_53),
.C(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_60),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_55),
.C(n_54),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_67),
.C(n_20),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_20),
.C(n_11),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_70),
.C(n_20),
.Y(n_71)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_12),
.B(n_11),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B1(n_3),
.B2(n_4),
.Y(n_73)
);

AOI332xp33_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_1),
.A3(n_3),
.B1(n_6),
.B2(n_8),
.B3(n_11),
.C1(n_72),
.C2(n_40),
.Y(n_74)
);


endmodule