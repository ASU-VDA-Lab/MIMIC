module real_jpeg_31503_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_0),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_0),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_0),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_533),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_1),
.B(n_534),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_4),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_4),
.Y(n_225)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_4),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_5),
.A2(n_205),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g268 ( 
.A1(n_5),
.A2(n_209),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g414 ( 
.A1(n_5),
.A2(n_209),
.B1(n_415),
.B2(n_418),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_5),
.A2(n_209),
.B1(n_458),
.B2(n_461),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_6),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_6),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

AO22x2_ASAP7_75t_L g153 ( 
.A1(n_8),
.A2(n_57),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_8),
.A2(n_57),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_8),
.A2(n_57),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_9),
.Y(n_124)
);

AOI22x1_ASAP7_75t_SL g95 ( 
.A1(n_10),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_10),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_10),
.A2(n_99),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g259 ( 
.A1(n_10),
.A2(n_99),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g435 ( 
.A(n_10),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_10),
.B(n_65),
.Y(n_453)
);

OAI32xp33_ASAP7_75t_L g472 ( 
.A1(n_10),
.A2(n_226),
.A3(n_473),
.B1(n_477),
.B2(n_484),
.Y(n_472)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_11),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_12),
.A2(n_27),
.B1(n_181),
.B2(n_185),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_12),
.A2(n_27),
.B1(n_222),
.B2(n_226),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_12),
.A2(n_27),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_13),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_193),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_191),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_160),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_19),
.B(n_161),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_62),
.B1(n_103),
.B2(n_104),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_21),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_30),
.B(n_52),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_23),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_31),
.B(n_53),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_31),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_31),
.B(n_204),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_SL g342 ( 
.A1(n_31),
.A2(n_107),
.B(n_171),
.Y(n_342)
);

NOR2x1p5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_44),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_34),
.Y(n_278)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_38),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_44),
.B(n_204),
.Y(n_203)
);

AO22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_45),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_46),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_48),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_49),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_49),
.Y(n_431)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_52),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_52),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_60),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_55),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_56),
.Y(n_174)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_56),
.Y(n_208)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_59),
.B(n_99),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_60),
.B(n_171),
.Y(n_318)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_61),
.B(n_99),
.Y(n_400)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_62),
.B(n_298),
.C(n_300),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_63),
.B(n_202),
.Y(n_201)
);

AOI21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_80),
.B(n_95),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_65),
.B(n_151),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g190 ( 
.A(n_65),
.B(n_153),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_65),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_SL g387 ( 
.A(n_65),
.B(n_268),
.Y(n_387)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AO21x2_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_81),
.B(n_88),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_74),
.B2(n_78),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_69),
.Y(n_420)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_79),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_79),
.Y(n_252)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g316 ( 
.A(n_80),
.B(n_95),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_88),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_98),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_98),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_99),
.A2(n_172),
.B(n_175),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g427 ( 
.A1(n_99),
.A2(n_428),
.A3(n_432),
.B1(n_434),
.B2(n_435),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_99),
.B(n_485),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_R g496 ( 
.A(n_99),
.B(n_115),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_99),
.B(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.C(n_148),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_106),
.B(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_111),
.B(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_168),
.C(n_177),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_113),
.A2(n_149),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_113),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g385 ( 
.A(n_113),
.B(n_386),
.C(n_388),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_113),
.A2(n_167),
.B1(n_386),
.B2(n_395),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_127),
.B(n_141),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_114),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_114),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_114),
.B(n_141),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_114),
.B(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_128),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B1(n_122),
.B2(n_125),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_117),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_120),
.Y(n_501)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_121),
.Y(n_261)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_126),
.Y(n_239)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_126),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_127),
.B(n_141),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_127),
.B(n_215),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_127),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_127),
.B(n_414),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_131),
.B1(n_134),
.B2(n_139),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_138),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_143),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_150),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_152),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_152),
.B(n_387),
.Y(n_386)
);

NAND2x1_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_159),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.C(n_176),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_369)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_167),
.B(n_178),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_168),
.A2(n_169),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_170),
.B(n_203),
.Y(n_388)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_175),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_176),
.B(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B(n_189),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_180),
.Y(n_335)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_189),
.B(n_267),
.Y(n_401)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NOR2x1_ASAP7_75t_L g315 ( 
.A(n_190),
.B(n_316),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21x1_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_376),
.B(n_528),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_352),
.B(n_355),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_321),
.B(n_323),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_296),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_198),
.B(n_296),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_242),
.C(n_264),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_200),
.B(n_242),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_211),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_202),
.Y(n_300)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_211),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_212),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_213),
.B(n_413),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_214),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_214),
.B(n_441),
.Y(n_451)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_217),
.Y(n_417)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_218),
.Y(n_433)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_L g389 ( 
.A(n_220),
.B(n_390),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_228),
.B(n_232),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_221),
.A2(n_255),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_227),
.Y(n_460)
);

AO21x2_ASAP7_75t_L g308 ( 
.A1(n_228),
.A2(n_230),
.B(n_309),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g506 ( 
.A1(n_228),
.A2(n_309),
.B(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_229),
.B(n_237),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_229),
.A2(n_259),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_229),
.B(n_457),
.Y(n_456)
);

INVx4_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_232),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_232),
.B(n_456),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_236),
.Y(n_295)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_SL g462 ( 
.A(n_239),
.Y(n_462)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2x2_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_254),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_244),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_313)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_252),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_253),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_253),
.B(n_413),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_255),
.B(n_507),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_256),
.B(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_264),
.B(n_380),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_272),
.C(n_274),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_265),
.A2(n_266),
.B1(n_272),
.B2(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_272),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_318),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_273),
.B(n_318),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_274),
.B(n_383),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_285),
.B(n_293),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_276),
.B(n_286),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.C(n_281),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_290),
.B(n_292),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_293),
.B(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_301),
.Y(n_296)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_311),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_307),
.B1(n_308),
.B2(n_310),
.Y(n_302)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_307),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_307),
.A2(n_308),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_342),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_308),
.A2(n_366),
.B(n_367),
.Y(n_365)
);

NOR2x1_ASAP7_75t_SL g442 ( 
.A(n_308),
.B(n_427),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_311),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

AOI22x1_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_314)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_319),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_320),
.Y(n_350)
);

NOR4xp25_ASAP7_75t_L g522 ( 
.A(n_321),
.B(n_353),
.C(n_523),
.D(n_526),
.Y(n_522)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_329),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_347),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_339),
.B1(n_345),
.B2(n_346),
.Y(n_330)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_331),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_348),
.C(n_372),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_334),
.B(n_338),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_334),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_333),
.B(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B(n_337),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_343),
.B2(n_344),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_346),
.Y(n_372)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.C(n_351),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_370),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_368),
.Y(n_357)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_358),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_363),
.C(n_365),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_359),
.A2(n_360),
.B1(n_363),
.B2(n_364),
.Y(n_375)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_365),
.Y(n_374)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_368),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_371),
.B(n_373),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_406),
.B(n_522),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_391),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_378),
.B(n_525),
.Y(n_524)
);

NAND2x1_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_379),
.B(n_381),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.C(n_389),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_405),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_389),
.Y(n_405)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_386),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_423),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_394),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_404),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_392),
.B(n_404),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.C(n_402),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_393),
.B(n_520),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_396),
.B(n_402),
.Y(n_520)
);

MAJx2_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_399),
.C(n_401),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_397),
.A2(n_399),
.B1(n_400),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_397),
.Y(n_445)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_401),
.Y(n_446)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

AO21x1_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_517),
.B(n_521),
.Y(n_407)
);

OAI21x1_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_447),
.B(n_516),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_438),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_410),
.B(n_438),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_421),
.C(n_424),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_422),
.Y(n_464)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_425),
.B(n_464),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_443),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_442),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_440),
.B(n_442),
.C(n_443),
.Y(n_518)
);

XOR2x2_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

AOI21x1_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_465),
.B(n_515),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_463),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_SL g515 ( 
.A(n_449),
.B(n_463),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.C(n_454),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_451),
.A2(n_452),
.B1(n_453),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_451),
.Y(n_469)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_504),
.Y(n_507)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_492),
.B(n_514),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_467),
.B(n_470),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_490),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_SL g511 ( 
.A(n_471),
.B(n_491),
.Y(n_511)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_472),
.B(n_490),
.Y(n_512)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

AOI21x1_ASAP7_75t_SL g492 ( 
.A1(n_493),
.A2(n_509),
.B(n_513),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_497),
.B(n_508),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_496),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_506),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

BUFx4f_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_511),
.C(n_512),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_510),
.A2(n_511),
.B(n_512),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_519),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_518),
.B(n_519),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

BUFx2_ASAP7_75t_SL g528 ( 
.A(n_529),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_531),
.C(n_532),
.Y(n_529)
);


endmodule