module fake_jpeg_22292_n_48 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_48);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_48;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_40;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_13),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_0),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_3),
.C(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_1),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_7),
.B(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_25),
.A3(n_27),
.B1(n_5),
.B2(n_6),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_36),
.B(n_37),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI22x1_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_33),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_16),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_17),
.C(n_18),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_19),
.C(n_20),
.Y(n_48)
);


endmodule