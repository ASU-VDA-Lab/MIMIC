module fake_jpeg_26482_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_66),
.Y(n_73)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_53),
.B1(n_55),
.B2(n_47),
.Y(n_79)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_57),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_60),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_0),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_48),
.B1(n_43),
.B2(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_52),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_58),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_63),
.B1(n_56),
.B2(n_46),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_92),
.B1(n_97),
.B2(n_81),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_61),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_51),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_56),
.B1(n_54),
.B2(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_96),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_4),
.B(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_45),
.B(n_5),
.C(n_7),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_107),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_90),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_111),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_113),
.B(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_86),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_22),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_24),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_21),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_26),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_120),
.B(n_121),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_70),
.C(n_106),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_119),
.B1(n_106),
.B2(n_118),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_107),
.B1(n_83),
.B2(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_4),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_8),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_29),
.C(n_37),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_117),
.B1(n_28),
.B2(n_15),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_125),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_25),
.B(n_35),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_20),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_17),
.B(n_19),
.C(n_31),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_34),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_39),
.Y(n_135)
);


endmodule