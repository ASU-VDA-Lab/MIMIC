module fake_netlist_1_6266_n_21 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_21;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
INVxp33_ASAP7_75t_SL g11 ( .A(n_3), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_1), .B(n_0), .Y(n_12) );
INVx3_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
AO21x1_ASAP7_75t_L g14 ( .A1(n_5), .A2(n_7), .B(n_8), .Y(n_14) );
INVx5_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
OR2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_0), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_16), .B(n_15), .Y(n_17) );
AOI211xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_14), .B(n_12), .C(n_11), .Y(n_18) );
NOR2x1_ASAP7_75t_L g19 ( .A(n_18), .B(n_4), .Y(n_19) );
XOR2x1_ASAP7_75t_L g20 ( .A(n_19), .B(n_6), .Y(n_20) );
OAI21xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_9), .B(n_10), .Y(n_21) );
endmodule