module fake_jpeg_4857_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_16),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_22),
.B1(n_32),
.B2(n_21),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_54),
.B(n_55),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_21),
.B1(n_32),
.B2(n_24),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_20),
.Y(n_87)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_22),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_82),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_43),
.B1(n_38),
.B2(n_39),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_85),
.B1(n_91),
.B2(n_92),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_78),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_43),
.B1(n_42),
.B2(n_45),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_60),
.B1(n_56),
.B2(n_47),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_21),
.B(n_16),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_94),
.B(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_25),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_93),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_44),
.B1(n_43),
.B2(n_35),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_42),
.B1(n_25),
.B2(n_18),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_42),
.B1(n_35),
.B2(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_18),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_33),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_99),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_51),
.A2(n_30),
.B(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_26),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_101),
.B(n_104),
.Y(n_147)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_103),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_110),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_70),
.B1(n_90),
.B2(n_73),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_86),
.C(n_74),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_111),
.C(n_113),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_41),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_41),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_115),
.B(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_124),
.Y(n_136)
);

NAND2x1_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_44),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_82),
.B(n_77),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_30),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_128),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_47),
.B1(n_66),
.B2(n_58),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_80),
.B1(n_89),
.B2(n_70),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_142),
.B1(n_151),
.B2(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_132),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_72),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_144),
.B(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_139),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_146),
.B1(n_152),
.B2(n_119),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_87),
.C(n_71),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_148),
.C(n_41),
.Y(n_181)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_106),
.B1(n_118),
.B2(n_114),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_121),
.A2(n_95),
.B1(n_98),
.B2(n_83),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_90),
.B(n_88),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_92),
.B1(n_76),
.B2(n_89),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_109),
.C(n_116),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_73),
.B1(n_24),
.B2(n_20),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_73),
.B1(n_88),
.B2(n_76),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_124),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_105),
.B(n_101),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_105),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_160),
.B(n_167),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_177),
.B1(n_159),
.B2(n_138),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_127),
.B(n_112),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_171),
.B(n_191),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_154),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_181),
.C(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_173),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_125),
.B(n_104),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_151),
.B1(n_134),
.B2(n_157),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_179),
.B1(n_184),
.B2(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_135),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_123),
.A3(n_103),
.B1(n_115),
.B2(n_120),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_178),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_137),
.B1(n_152),
.B2(n_150),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_35),
.B1(n_32),
.B2(n_20),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_35),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_103),
.B1(n_24),
.B2(n_36),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_44),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_186),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_133),
.A2(n_36),
.B1(n_58),
.B2(n_44),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_44),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_41),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_41),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_150),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_36),
.B1(n_31),
.B2(n_27),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_17),
.B(n_27),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_27),
.B(n_17),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_149),
.B(n_27),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_193),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_194),
.B(n_196),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_211),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_213),
.C(n_214),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_154),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_209),
.B(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_212),
.B1(n_218),
.B2(n_170),
.Y(n_235)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_31),
.B1(n_27),
.B2(n_17),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_27),
.C(n_17),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_17),
.C(n_31),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_217),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_186),
.B(n_31),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_SL g218 ( 
.A1(n_169),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_219),
.A2(n_179),
.B1(n_170),
.B2(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_161),
.A2(n_2),
.B(n_3),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_194),
.B(n_165),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_225),
.B(n_236),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_161),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_167),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_240),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_197),
.B(n_219),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_196),
.B(n_160),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_169),
.B(n_192),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_248),
.B(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_239),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_174),
.B1(n_171),
.B2(n_163),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_247),
.B1(n_218),
.B2(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_243),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_202),
.B(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_188),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_244),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_195),
.A2(n_164),
.B1(n_189),
.B2(n_5),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_245),
.A2(n_235),
.B1(n_240),
.B2(n_232),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_206),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_200),
.A2(n_3),
.B(n_4),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_205),
.C(n_214),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_259),
.C(n_264),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_255),
.B(n_248),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

AO221x1_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_269),
.B1(n_233),
.B2(n_223),
.C(n_198),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_215),
.C(n_216),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_211),
.C(n_220),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_270),
.B1(n_4),
.B2(n_5),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_207),
.B(n_195),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_262),
.A2(n_223),
.B(n_234),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_207),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_218),
.C(n_217),
.Y(n_267)
);

OAI322xp33_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_229),
.A3(n_224),
.B1(n_239),
.B2(n_12),
.C1(n_9),
.C2(n_10),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_198),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_238),
.Y(n_271)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_276),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_266),
.A2(n_245),
.B1(n_242),
.B2(n_233),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_277),
.B1(n_282),
.B2(n_284),
.Y(n_302)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_285),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_281),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_255),
.A2(n_244),
.B1(n_231),
.B2(n_247),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_280),
.C(n_261),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_9),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_4),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_287),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_286),
.B1(n_253),
.B2(n_262),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_5),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_254),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_264),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_298),
.B1(n_290),
.B2(n_299),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_290),
.A2(n_10),
.B(n_12),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_292),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_259),
.C(n_250),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_296),
.C(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_302),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_251),
.C(n_252),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_277),
.A2(n_258),
.B1(n_265),
.B2(n_257),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_301),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_276),
.B(n_252),
.C(n_263),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_278),
.B1(n_287),
.B2(n_279),
.Y(n_301)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_286),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_309),
.B(n_311),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_294),
.A2(n_272),
.B(n_274),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_312),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_285),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_272),
.C(n_281),
.Y(n_312)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_13),
.B(n_14),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_6),
.C(n_7),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_7),
.Y(n_322)
);

AOI21x1_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_291),
.B(n_293),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_317),
.A2(n_318),
.B(n_322),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_300),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_14),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_328),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_312),
.Y(n_327)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_303),
.C(n_306),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_314),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_329),
.B(n_330),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_316),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_315),
.B(n_316),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_303),
.C(n_331),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_330),
.C(n_326),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_324),
.Y(n_338)
);


endmodule