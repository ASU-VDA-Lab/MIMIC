module fake_jpeg_30719_n_93 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx4f_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_1),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_52),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_8),
.B(n_10),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_59),
.B(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_4),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_56),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_53),
.Y(n_71)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_27),
.B(n_5),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_58),
.Y(n_72)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_6),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_33),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_28),
.B(n_21),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_26),
.Y(n_64)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_77),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_52),
.B1(n_48),
.B2(n_54),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_75),
.A2(n_76),
.B(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_46),
.B1(n_45),
.B2(n_55),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_76),
.Y(n_81)
);

XOR2x1_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_75),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_70),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_83),
.C(n_68),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_70),
.C(n_72),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_67),
.Y(n_86)
);

AOI221xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_49),
.B1(n_34),
.B2(n_79),
.C(n_42),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_87),
.C(n_32),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_89),
.C(n_34),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_40),
.C(n_39),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_51),
.B1(n_34),
.B2(n_42),
.Y(n_93)
);


endmodule