module fake_jpeg_29993_n_195 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_195);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_12),
.B(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_6),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_13),
.B(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_23),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_28),
.B1(n_17),
.B2(n_26),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_47),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_23),
.B1(n_22),
.B2(n_25),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_50),
.A2(n_61),
.B1(n_51),
.B2(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_15),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_32),
.A2(n_28),
.B1(n_18),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_16),
.B1(n_27),
.B2(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_31),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_49),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_23),
.B1(n_22),
.B2(n_27),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_67),
.B1(n_44),
.B2(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_89),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_92),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_73),
.B1(n_79),
.B2(n_84),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_30),
.B1(n_35),
.B2(n_27),
.Y(n_73)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_24),
.B(n_21),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_78),
.B(n_86),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_19),
.B1(n_24),
.B2(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_16),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_87),
.C(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_35),
.B1(n_19),
.B2(n_2),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_8),
.B1(n_11),
.B2(n_2),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_35),
.C(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_3),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_46),
.C(n_63),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_3),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_87),
.B1(n_73),
.B2(n_76),
.Y(n_122)
);

NOR2x1_ASAP7_75t_R g98 ( 
.A(n_61),
.B(n_0),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_1),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_49),
.B1(n_54),
.B2(n_4),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_120),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_98),
.B1(n_74),
.B2(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_113),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_9),
.B1(n_11),
.B2(n_0),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_78),
.B(n_83),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_102),
.B(n_117),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_1),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_86),
.A2(n_82),
.B1(n_93),
.B2(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_84),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_68),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_76),
.B1(n_90),
.B2(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_103),
.Y(n_138)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_75),
.C(n_68),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_132),
.C(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_134),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_133),
.A2(n_102),
.B(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_109),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_105),
.B1(n_123),
.B2(n_110),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_145),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_105),
.B(n_115),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_112),
.Y(n_161)
);

OAI221xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_101),
.B1(n_100),
.B2(n_108),
.C(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_134),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_106),
.B1(n_114),
.B2(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_112),
.B1(n_126),
.B2(n_130),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_124),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_112),
.C(n_127),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_131),
.C(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_152),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_155),
.B(n_154),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_164),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_130),
.C(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_160),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_161),
.A2(n_150),
.B1(n_146),
.B2(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_144),
.B(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_163),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_153),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_154),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_172),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_159),
.A2(n_149),
.B1(n_143),
.B2(n_141),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_142),
.B(n_143),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_156),
.C(n_166),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_167),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_175),
.B1(n_168),
.B2(n_173),
.Y(n_184)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_164),
.C(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_181),
.B(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_173),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_183),
.A2(n_186),
.B(n_177),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_184),
.A2(n_185),
.B1(n_180),
.B2(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_187),
.A2(n_186),
.B(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_189),
.B(n_180),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_188),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_192),
.Y(n_195)
);


endmodule