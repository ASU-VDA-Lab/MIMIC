module fake_netlist_6_4344_n_763 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_763);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_763;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_544;
wire n_468;
wire n_372;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_550;
wire n_487;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx2_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_86),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_50),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_21),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_11),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_65),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_87),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_5),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_25),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_69),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_89),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_56),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_116),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_28),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_97),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_73),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_67),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_90),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_24),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_55),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_115),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_15),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_77),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_111),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_70),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_99),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_68),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_47),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_80),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_118),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_0),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_34),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_81),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_51),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_71),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_15),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_22),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_91),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_126),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_121),
.Y(n_192)
);

BUFx4f_ASAP7_75t_SL g193 ( 
.A(n_38),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_24),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_22),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_62),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_0),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_146),
.B(n_144),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_1),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_173),
.B(n_2),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_2),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_26),
.Y(n_207)
);

BUFx8_ASAP7_75t_SL g208 ( 
.A(n_165),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_156),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_148),
.B(n_3),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_3),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_4),
.Y(n_212)
);

BUFx8_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_27),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_161),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_4),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_5),
.Y(n_219)
);

BUFx8_ASAP7_75t_SL g220 ( 
.A(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_171),
.B(n_6),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

BUFx8_ASAP7_75t_SL g225 ( 
.A(n_188),
.Y(n_225)
);

BUFx8_ASAP7_75t_SL g226 ( 
.A(n_189),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_6),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_7),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_183),
.B(n_7),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_159),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_196),
.B1(n_172),
.B2(n_145),
.Y(n_237)
);

AO22x2_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_8),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_145),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_201),
.A2(n_196),
.B1(n_172),
.B2(n_192),
.Y(n_244)
);

AO22x2_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_201),
.A2(n_174),
.B1(n_191),
.B2(n_186),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_160),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_235),
.A2(n_185),
.B1(n_180),
.B2(n_179),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_209),
.B1(n_217),
.B2(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_204),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_211),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_166),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_170),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_177),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_193),
.B1(n_13),
.B2(n_14),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_12),
.B1(n_16),
.B2(n_17),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_219),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_L g264 ( 
.A1(n_198),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_202),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_198),
.A2(n_23),
.B1(n_29),
.B2(n_30),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_219),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_33),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_200),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_39),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_40),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_200),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_202),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_212),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_224),
.B(n_48),
.Y(n_275)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_199),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_212),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_223),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_223),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_281)
);

AO22x2_ASAP7_75t_L g282 ( 
.A1(n_203),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_229),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_250),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_247),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_236),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_256),
.A2(n_207),
.B(n_214),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_228),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_254),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_240),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_239),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_280),
.B(n_207),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_255),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_243),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_222),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_246),
.B(n_228),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_249),
.A2(n_207),
.B(n_214),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_244),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_281),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_R g314 ( 
.A(n_282),
.B(n_207),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_236),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_260),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_276),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_260),
.B(n_214),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_269),
.A2(n_214),
.B(n_233),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_238),
.Y(n_327)
);

OR2x2_ASAP7_75t_SL g328 ( 
.A(n_245),
.B(n_218),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_272),
.B(n_203),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_264),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_261),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_279),
.A2(n_227),
.B(n_222),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_274),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_253),
.A2(n_210),
.B(n_229),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_242),
.B(n_236),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_275),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_257),
.B(n_233),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_251),
.Y(n_342)
);

OR2x6_ASAP7_75t_L g343 ( 
.A(n_238),
.B(n_197),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_251),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

BUFx4f_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_292),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_289),
.B(n_286),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_290),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_285),
.B(n_210),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_321),
.B(n_233),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_342),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_286),
.B(n_226),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_321),
.B(n_233),
.Y(n_364)
);

NAND2x1p5_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_215),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_340),
.B(n_233),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_304),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_306),
.B(n_233),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_310),
.B(n_225),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_284),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_313),
.B(n_227),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_227),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_308),
.B(n_227),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_284),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_287),
.B(n_227),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_309),
.B(n_227),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_315),
.B(n_222),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_222),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_305),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_299),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_222),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_301),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_334),
.B(n_222),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_213),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_337),
.B(n_215),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_326),
.B(n_215),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_296),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_297),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_298),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_323),
.A2(n_206),
.B(n_213),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_215),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_331),
.B(n_215),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

AND2x4_ASAP7_75t_L g403 ( 
.A(n_329),
.B(n_88),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_330),
.B(n_213),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

AND2x4_ASAP7_75t_SL g406 ( 
.A(n_322),
.B(n_215),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_325),
.B(n_213),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_316),
.B(n_319),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_311),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_336),
.B(n_230),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_317),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_387),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_374),
.B(n_324),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

BUFx4f_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_324),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_343),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_312),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_291),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

BUFx4f_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_353),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_354),
.B(n_208),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_291),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_349),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_349),
.B(n_343),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_386),
.B(n_327),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_358),
.B(n_327),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_358),
.B(n_332),
.Y(n_439)
);

NAND2x1p5_ASAP7_75t_L g440 ( 
.A(n_348),
.B(n_206),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

HB1xp67_ASAP7_75t_SL g442 ( 
.A(n_410),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_387),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_352),
.Y(n_444)
);

BUFx5_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_L g446 ( 
.A(n_369),
.B(n_230),
.Y(n_446)
);

AND2x2_ASAP7_75t_SL g447 ( 
.A(n_348),
.B(n_220),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_343),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_387),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_392),
.B(n_314),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

OR2x6_ASAP7_75t_L g454 ( 
.A(n_347),
.B(n_230),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_347),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_357),
.B(n_92),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_357),
.B(n_93),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_355),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_405),
.B(n_314),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_355),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_405),
.B(n_206),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_359),
.B(n_362),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_375),
.B(n_197),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_393),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_348),
.B(n_197),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_363),
.B(n_94),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_443),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_415),
.B(n_375),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_360),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g475 ( 
.A(n_429),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_444),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_416),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_443),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_451),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_416),
.Y(n_480)
);

INVx5_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_451),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_462),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_448),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_453),
.Y(n_487)
);

CKINVDCx11_ASAP7_75t_R g488 ( 
.A(n_454),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_462),
.Y(n_491)
);

INVx3_ASAP7_75t_SL g492 ( 
.A(n_442),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_459),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_455),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_439),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_461),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_417),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_425),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_428),
.Y(n_503)
);

INVx8_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_415),
.B(n_381),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_437),
.Y(n_507)
);

BUFx12f_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

INVx3_ASAP7_75t_SL g509 ( 
.A(n_442),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_418),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_360),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_419),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

NAND2x1p5_ASAP7_75t_L g514 ( 
.A(n_428),
.B(n_387),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_425),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_494),
.Y(n_517)
);

BUFx12f_ASAP7_75t_L g518 ( 
.A(n_488),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_475),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_510),
.Y(n_520)
);

OAI22x1_ASAP7_75t_L g521 ( 
.A1(n_492),
.A2(n_431),
.B1(n_426),
.B2(n_423),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_506),
.A2(n_348),
.B1(n_423),
.B2(n_431),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_510),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_492),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_506),
.A2(n_426),
.B1(n_347),
.B2(n_382),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_490),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_492),
.Y(n_527)
);

INVx8_ASAP7_75t_L g528 ( 
.A(n_504),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_490),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_SL g530 ( 
.A1(n_495),
.A2(n_430),
.B1(n_447),
.B2(n_347),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_473),
.A2(n_347),
.B1(n_382),
.B2(n_381),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_476),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g533 ( 
.A1(n_504),
.A2(n_347),
.B1(n_468),
.B2(n_367),
.Y(n_533)
);

INVx6_ASAP7_75t_L g534 ( 
.A(n_475),
.Y(n_534)
);

CKINVDCx11_ASAP7_75t_R g535 ( 
.A(n_509),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_509),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_471),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_507),
.A2(n_403),
.B1(n_469),
.B2(n_452),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_485),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_504),
.A2(n_468),
.B1(n_465),
.B2(n_439),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_504),
.A2(n_452),
.B1(n_460),
.B2(n_435),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_478),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_485),
.Y(n_543)
);

BUFx4f_ASAP7_75t_SL g544 ( 
.A(n_509),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_507),
.B(n_435),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_511),
.A2(n_356),
.B(n_378),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_504),
.A2(n_460),
.B1(n_387),
.B2(n_414),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_511),
.A2(n_464),
.B1(n_467),
.B2(n_450),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_511),
.A2(n_414),
.B1(n_407),
.B2(n_450),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_476),
.Y(n_551)
);

CKINVDCx11_ASAP7_75t_R g552 ( 
.A(n_499),
.Y(n_552)
);

CKINVDCx11_ASAP7_75t_R g553 ( 
.A(n_499),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_511),
.A2(n_371),
.B1(n_446),
.B2(n_434),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_496),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_512),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_486),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_521),
.A2(n_408),
.B1(n_390),
.B2(n_456),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_522),
.A2(n_457),
.B1(n_449),
.B2(n_364),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_513),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_457),
.B1(n_364),
.B2(n_434),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_544),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_520),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_523),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_555),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_548),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_526),
.B(n_513),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_530),
.A2(n_454),
.B1(n_368),
.B2(n_411),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_535),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_540),
.A2(n_454),
.B1(n_368),
.B2(n_411),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_549),
.A2(n_391),
.B1(n_432),
.B2(n_496),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_549),
.A2(n_391),
.B1(n_373),
.B2(n_370),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_555),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_538),
.A2(n_380),
.B(n_389),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_524),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_533),
.A2(n_373),
.B1(n_362),
.B2(n_370),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_545),
.A2(n_359),
.B1(n_372),
.B2(n_436),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_538),
.A2(n_436),
.B1(n_421),
.B2(n_500),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_545),
.A2(n_372),
.B1(n_474),
.B2(n_498),
.Y(n_579)
);

INVx5_ASAP7_75t_SL g580 ( 
.A(n_537),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_529),
.B(n_525),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_554),
.A2(n_404),
.B1(n_498),
.B2(n_503),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_556),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_518),
.A2(n_398),
.B1(n_498),
.B2(n_501),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_525),
.A2(n_474),
.B1(n_498),
.B2(n_501),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_536),
.A2(n_508),
.B1(n_500),
.B2(n_516),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_546),
.A2(n_409),
.B(n_406),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_529),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_528),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_541),
.A2(n_531),
.B1(n_550),
.B2(n_527),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_531),
.A2(n_409),
.B(n_406),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_532),
.B(n_472),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_532),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_547),
.A2(n_474),
.B1(n_501),
.B2(n_498),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_539),
.A2(n_474),
.B1(n_501),
.B2(n_498),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_534),
.A2(n_433),
.B1(n_516),
.B2(n_400),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_543),
.A2(n_503),
.B1(n_501),
.B2(n_508),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_552),
.A2(n_501),
.B1(n_503),
.B2(n_366),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_537),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_551),
.Y(n_600)
);

BUFx12f_ASAP7_75t_L g601 ( 
.A(n_552),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_551),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_518),
.A2(n_503),
.B1(n_406),
.B2(n_494),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_557),
.B(n_472),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_568),
.A2(n_570),
.B1(n_559),
.B2(n_561),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_558),
.A2(n_503),
.B1(n_553),
.B2(n_388),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_578),
.A2(n_503),
.B1(n_388),
.B2(n_534),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_576),
.A2(n_534),
.B1(n_396),
.B2(n_515),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_579),
.A2(n_515),
.B1(n_519),
.B2(n_433),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_590),
.A2(n_515),
.B1(n_433),
.B2(n_400),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_577),
.A2(n_514),
.B1(n_402),
.B2(n_400),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_586),
.A2(n_528),
.B1(n_514),
.B2(n_517),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_571),
.A2(n_515),
.B1(n_402),
.B2(n_505),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_SL g614 ( 
.A1(n_601),
.A2(n_528),
.B1(n_514),
.B2(n_517),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_598),
.A2(n_587),
.B1(n_595),
.B2(n_597),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_572),
.A2(n_402),
.B1(n_494),
.B2(n_413),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_601),
.A2(n_515),
.B1(n_505),
.B2(n_383),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_591),
.A2(n_494),
.B1(n_502),
.B2(n_515),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_582),
.A2(n_584),
.B1(n_573),
.B2(n_585),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_594),
.A2(n_505),
.B1(n_383),
.B2(n_502),
.Y(n_620)
);

OAI222xp33_ASAP7_75t_L g621 ( 
.A1(n_603),
.A2(n_484),
.B1(n_493),
.B2(n_497),
.C1(n_365),
.C2(n_557),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_565),
.A2(n_413),
.B1(n_502),
.B2(n_497),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_574),
.A2(n_505),
.B1(n_502),
.B2(n_493),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_575),
.A2(n_379),
.B1(n_542),
.B2(n_484),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_575),
.A2(n_413),
.B1(n_377),
.B2(n_376),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_560),
.B(n_486),
.Y(n_626)
);

OAI211xp5_ASAP7_75t_SL g627 ( 
.A1(n_563),
.A2(n_413),
.B(n_384),
.C(n_385),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_569),
.A2(n_384),
.B1(n_365),
.B2(n_395),
.Y(n_628)
);

OAI221xp5_ASAP7_75t_SL g629 ( 
.A1(n_562),
.A2(n_487),
.B1(n_491),
.B2(n_470),
.C(n_463),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_564),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_SL g631 ( 
.A1(n_596),
.A2(n_542),
.B1(n_537),
.B2(n_365),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_SL g632 ( 
.A1(n_565),
.A2(n_487),
.B1(n_477),
.B2(n_480),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_581),
.A2(n_395),
.B1(n_445),
.B2(n_361),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_581),
.A2(n_395),
.B1(n_445),
.B2(n_361),
.Y(n_634)
);

OAI221xp5_ASAP7_75t_SL g635 ( 
.A1(n_562),
.A2(n_491),
.B1(n_470),
.B2(n_463),
.C(n_480),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_569),
.A2(n_478),
.B1(n_481),
.B2(n_470),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_566),
.A2(n_395),
.B1(n_445),
.B2(n_361),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_583),
.A2(n_567),
.B1(n_560),
.B2(n_589),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_567),
.A2(n_445),
.B1(n_361),
.B2(n_477),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_589),
.A2(n_445),
.B1(n_477),
.B2(n_480),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_630),
.B(n_602),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_624),
.B(n_606),
.C(n_625),
.Y(n_642)
);

OAI22xp33_ASAP7_75t_L g643 ( 
.A1(n_615),
.A2(n_589),
.B1(n_592),
.B2(n_604),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_630),
.B(n_588),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_638),
.B(n_593),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_626),
.B(n_600),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_619),
.B(n_604),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_607),
.B(n_592),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_625),
.B(n_599),
.Y(n_649)
);

OA211x2_ASAP7_75t_L g650 ( 
.A1(n_617),
.A2(n_580),
.B(n_599),
.C(n_537),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_605),
.A2(n_580),
.B1(n_599),
.B2(n_478),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_609),
.B(n_599),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_610),
.B(n_580),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_623),
.B(n_580),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_628),
.B(n_480),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_636),
.A2(n_479),
.B1(n_471),
.B2(n_483),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_631),
.B(n_477),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_628),
.B(n_618),
.Y(n_658)
);

NAND3xp33_ASAP7_75t_L g659 ( 
.A(n_629),
.B(n_483),
.C(n_482),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_613),
.B(n_491),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_612),
.B(n_95),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_608),
.A2(n_478),
.B1(n_481),
.B2(n_489),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_633),
.B(n_96),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_632),
.B(n_479),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_635),
.B(n_479),
.C(n_483),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_614),
.B(n_98),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_611),
.A2(n_479),
.B1(n_483),
.B2(n_482),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_616),
.A2(n_489),
.B1(n_478),
.B2(n_481),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_641),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_642),
.B(n_620),
.C(n_627),
.Y(n_670)
);

AO21x2_ASAP7_75t_L g671 ( 
.A1(n_664),
.A2(n_621),
.B(n_622),
.Y(n_671)
);

NAND4xp75_ASAP7_75t_L g672 ( 
.A(n_650),
.B(n_100),
.C(n_101),
.D(n_103),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_641),
.B(n_634),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_658),
.B(n_647),
.C(n_649),
.Y(n_674)
);

AOI221xp5_ASAP7_75t_L g675 ( 
.A1(n_643),
.A2(n_639),
.B1(n_637),
.B2(n_640),
.C(n_483),
.Y(n_675)
);

OAI211xp5_ASAP7_75t_SL g676 ( 
.A1(n_658),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_676)
);

NAND2x1_ASAP7_75t_L g677 ( 
.A(n_644),
.B(n_483),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_644),
.B(n_107),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_645),
.B(n_657),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_651),
.A2(n_489),
.B1(n_482),
.B2(n_479),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_661),
.B(n_109),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_645),
.B(n_110),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_659),
.B(n_482),
.C(n_479),
.Y(n_683)
);

NAND3xp33_ASAP7_75t_SL g684 ( 
.A(n_666),
.B(n_440),
.C(n_489),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_646),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_674),
.B(n_664),
.C(n_665),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_679),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_685),
.B(n_657),
.Y(n_688)
);

NAND4xp75_ASAP7_75t_L g689 ( 
.A(n_682),
.B(n_652),
.C(n_663),
.D(n_655),
.Y(n_689)
);

XNOR2x2_ASAP7_75t_L g690 ( 
.A(n_683),
.B(n_648),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_669),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_679),
.B(n_654),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_678),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_683),
.B(n_656),
.Y(n_694)
);

XNOR2xp5_ASAP7_75t_L g695 ( 
.A(n_670),
.B(n_663),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_692),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_688),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_R g698 ( 
.A(n_690),
.B(n_681),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_695),
.A2(n_670),
.B1(n_673),
.B2(n_672),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_687),
.B(n_677),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_698),
.A2(n_686),
.B1(n_689),
.B2(n_694),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_698),
.A2(n_694),
.B1(n_687),
.B2(n_684),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_700),
.Y(n_703)
);

OA22x2_ASAP7_75t_L g704 ( 
.A1(n_699),
.A2(n_693),
.B1(n_691),
.B2(n_653),
.Y(n_704)
);

OAI22x1_ASAP7_75t_L g705 ( 
.A1(n_696),
.A2(n_693),
.B1(n_671),
.B2(n_660),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_703),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_704),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_701),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_702),
.Y(n_709)
);

AOI221xp5_ASAP7_75t_L g710 ( 
.A1(n_708),
.A2(n_705),
.B1(n_697),
.B2(n_676),
.C(n_671),
.Y(n_710)
);

AOI32xp33_ASAP7_75t_L g711 ( 
.A1(n_709),
.A2(n_693),
.A3(n_680),
.B1(n_667),
.B2(n_675),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_706),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_712),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_711),
.Y(n_714)
);

OAI22x1_ASAP7_75t_L g715 ( 
.A1(n_710),
.A2(n_707),
.B1(n_706),
.B2(n_662),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_710),
.A2(n_668),
.B1(n_482),
.B2(n_471),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_714),
.B(n_482),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_713),
.B(n_113),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_715),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_716),
.Y(n_720)
);

AOI221xp5_ASAP7_75t_L g721 ( 
.A1(n_715),
.A2(n_471),
.B1(n_117),
.B2(n_120),
.C(n_122),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_714),
.B(n_471),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_713),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_722),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_723),
.Y(n_725)
);

NOR3xp33_ASAP7_75t_L g726 ( 
.A(n_718),
.B(n_114),
.C(n_123),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_720),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_719),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_717),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_721),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_728),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_724),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_725),
.Y(n_733)
);

NAND4xp25_ASAP7_75t_L g734 ( 
.A(n_730),
.B(n_124),
.C(n_127),
.D(n_128),
.Y(n_734)
);

INVxp67_ASAP7_75t_SL g735 ( 
.A(n_729),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_727),
.B(n_129),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_726),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_726),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_731),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_735),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_732),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_733),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_736),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_737),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_738),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_744),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_745),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_739),
.A2(n_734),
.B1(n_471),
.B2(n_478),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_741),
.A2(n_481),
.B1(n_440),
.B2(n_206),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_742),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_748),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_746),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_747),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_751),
.B(n_743),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_SL g756 ( 
.A1(n_753),
.A2(n_752),
.B1(n_754),
.B2(n_755),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_753),
.A2(n_749),
.B1(n_750),
.B2(n_481),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_756),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_757),
.Y(n_759)
);

AOI211xp5_ASAP7_75t_L g760 ( 
.A1(n_758),
.A2(n_133),
.B(n_135),
.C(n_136),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_760),
.Y(n_761)
);

AOI221xp5_ASAP7_75t_L g762 ( 
.A1(n_761),
.A2(n_759),
.B1(n_481),
.B2(n_139),
.C(n_140),
.Y(n_762)
);

AOI211xp5_ASAP7_75t_L g763 ( 
.A1(n_762),
.A2(n_137),
.B(n_138),
.C(n_142),
.Y(n_763)
);


endmodule