module fake_jpeg_28778_n_356 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_356);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_356;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_9),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_45),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_6),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_8),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx9p33_ASAP7_75t_R g101 ( 
.A(n_56),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_5),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_74),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_28),
.B(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_76),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_4),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_42),
.B1(n_43),
.B2(n_36),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_84),
.B1(n_127),
.B2(n_17),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_35),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_42),
.B1(n_78),
.B2(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_104),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_35),
.B1(n_34),
.B2(n_37),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_86),
.A2(n_31),
.B1(n_17),
.B2(n_19),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_44),
.B(n_27),
.C(n_16),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_93),
.B(n_11),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_37),
.B1(n_34),
.B2(n_39),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_99),
.B1(n_116),
.B2(n_29),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_37),
.B1(n_39),
.B2(n_29),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_44),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_61),
.B(n_16),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_46),
.B(n_27),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_119),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_58),
.A2(n_29),
.B1(n_23),
.B2(n_40),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_46),
.B(n_36),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_64),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_0),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_47),
.A2(n_19),
.B1(n_24),
.B2(n_20),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_120),
.B1(n_93),
.B2(n_95),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_143),
.B1(n_149),
.B2(n_154),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_136),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_23),
.C(n_31),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_92),
.Y(n_164)
);

BUFx2_ASAP7_75t_SL g132 ( 
.A(n_101),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_132),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_133),
.B(n_134),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_153),
.Y(n_170)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_89),
.Y(n_139)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_79),
.A2(n_23),
.B(n_20),
.C(n_30),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_88),
.CI(n_105),
.CON(n_174),
.SN(n_174)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_25),
.B1(n_23),
.B2(n_30),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_0),
.B(n_1),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_88),
.B(n_107),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_115),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_25),
.B1(n_11),
.B2(n_4),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_87),
.B(n_80),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_97),
.A2(n_12),
.B1(n_15),
.B2(n_2),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_99),
.A2(n_15),
.B1(n_12),
.B2(n_1),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_159),
.B1(n_162),
.B2(n_107),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_1),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_161),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_94),
.A2(n_12),
.B1(n_108),
.B2(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_108),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_94),
.A2(n_121),
.B1(n_98),
.B2(n_110),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_117),
.A2(n_122),
.B1(n_91),
.B2(n_90),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_163),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_141),
.C(n_155),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_132),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_169),
.B(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_102),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_174),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_178),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_105),
.B(n_122),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_189),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_154),
.B1(n_134),
.B2(n_135),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_115),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_182),
.B(n_174),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_184),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_91),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_133),
.A2(n_98),
.B1(n_110),
.B2(n_90),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_162),
.B1(n_151),
.B2(n_135),
.Y(n_198)
);

AO22x2_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_103),
.B1(n_117),
.B2(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_160),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_191),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_142),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_144),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_138),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_137),
.B(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_139),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_203),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_185),
.B1(n_183),
.B2(n_180),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_159),
.B1(n_152),
.B2(n_148),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_131),
.B1(n_155),
.B2(n_141),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_185),
.B1(n_197),
.B2(n_193),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_182),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_212),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_220),
.C(n_201),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_225),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_166),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_139),
.C(n_156),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_189),
.C(n_175),
.Y(n_249)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_223),
.Y(n_252)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_170),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_176),
.B(n_170),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_173),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_238),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_236),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_237),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_189),
.B1(n_168),
.B2(n_174),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_212),
.B(n_196),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_249),
.C(n_204),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_195),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_244),
.Y(n_264)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_202),
.B(n_189),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_205),
.A2(n_168),
.B(n_165),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_250),
.A2(n_233),
.B(n_243),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_189),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_181),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_231),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_258),
.C(n_265),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_205),
.B(n_199),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_257),
.A2(n_262),
.B(n_244),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_234),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_186),
.Y(n_280)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_223),
.B(n_210),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_268),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_226),
.C(n_211),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_198),
.B1(n_216),
.B2(n_203),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_266),
.A2(n_230),
.B1(n_240),
.B2(n_241),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_267),
.B(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_272),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_213),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_229),
.C(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_256),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_231),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_278),
.C(n_285),
.Y(n_300)
);

NOR4xp25_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_237),
.C(n_236),
.D(n_233),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_282),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_229),
.Y(n_278)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_274),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_216),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_293),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_257),
.B(n_260),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_246),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_292),
.C(n_272),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_271),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_253),
.B1(n_235),
.B2(n_264),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_267),
.B(n_252),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_252),
.B1(n_254),
.B2(n_256),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_289),
.Y(n_294)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_266),
.B1(n_273),
.B2(n_230),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_298),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_291),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_297),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_254),
.B1(n_264),
.B2(n_262),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_305),
.C(n_301),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_301),
.B(n_306),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_255),
.B(n_260),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_303),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_255),
.B1(n_269),
.B2(n_268),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_279),
.C(n_278),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_308),
.C(n_261),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_311),
.B(n_313),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_279),
.C(n_286),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_275),
.C(n_292),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_316),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_302),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_SL g319 ( 
.A1(n_303),
.A2(n_259),
.B(n_234),
.C(n_188),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_319),
.A2(n_294),
.B(n_297),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_304),
.B(n_213),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_320),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_307),
.B(n_227),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_309),
.Y(n_329)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_323),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_305),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_328),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_306),
.B1(n_295),
.B2(n_309),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_329),
.B(n_331),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_332),
.C(n_317),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_296),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_263),
.C(n_239),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_321),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_334),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_338),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g336 ( 
.A(n_326),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_336),
.B(n_319),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_317),
.Y(n_338)
);

AOI322xp5_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_325),
.A3(n_314),
.B1(n_327),
.B2(n_319),
.C1(n_324),
.C2(n_332),
.Y(n_342)
);

AOI21x1_ASAP7_75t_SL g347 ( 
.A1(n_342),
.A2(n_336),
.B(n_333),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_343),
.B(n_344),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_337),
.A2(n_247),
.B1(n_248),
.B2(n_245),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_340),
.A2(n_247),
.B(n_245),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_345),
.B(n_215),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_347),
.A2(n_349),
.B(n_350),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_219),
.C(n_206),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_348),
.A2(n_346),
.B(n_342),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_248),
.Y(n_353)
);

AOI322xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_351),
.A3(n_234),
.B1(n_206),
.B2(n_209),
.C1(n_222),
.C2(n_221),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_354),
.B(n_169),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g356 ( 
.A(n_355),
.B(n_218),
.CI(n_209),
.CON(n_356),
.SN(n_356)
);


endmodule