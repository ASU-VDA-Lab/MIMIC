module fake_jpeg_16584_n_353 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_50),
.Y(n_61)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_54),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_21),
.C(n_33),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_33),
.C(n_37),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_30),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_21),
.B1(n_23),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_21),
.B1(n_23),
.B2(n_32),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_27),
.B1(n_19),
.B2(n_25),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_32),
.B1(n_21),
.B2(n_23),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_21),
.B(n_39),
.C(n_29),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_71),
.Y(n_85)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_34),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_29),
.B1(n_24),
.B2(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_29),
.B1(n_30),
.B2(n_20),
.Y(n_109)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_81),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_83),
.Y(n_117)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_37),
.B1(n_35),
.B2(n_26),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_82),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_61),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_88),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

NAND2x1_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_38),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_59),
.B(n_69),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_100),
.Y(n_129)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_104),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_18),
.B1(n_19),
.B2(n_25),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_71),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_24),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_24),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_28),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_106),
.A2(n_109),
.B1(n_27),
.B2(n_20),
.Y(n_122)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_124),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_65),
.B(n_68),
.C(n_62),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_125),
.B(n_90),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_R g121 ( 
.A(n_93),
.B(n_55),
.C(n_28),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_133),
.Y(n_145)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_158)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

OAI22x1_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_59),
.C(n_75),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_59),
.C(n_92),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_77),
.B1(n_73),
.B2(n_64),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_108),
.B1(n_80),
.B2(n_77),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_85),
.B1(n_99),
.B2(n_94),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_167),
.B1(n_73),
.B2(n_64),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_79),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_148),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_83),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_153),
.B(n_161),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_85),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_104),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_166),
.C(n_31),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_154),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_151),
.A2(n_152),
.B1(n_162),
.B2(n_165),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_97),
.B1(n_87),
.B2(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_102),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_100),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_159),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_112),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_157),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_105),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_92),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_91),
.B1(n_70),
.B2(n_80),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_113),
.B1(n_111),
.B2(n_63),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_64),
.B1(n_66),
.B2(n_81),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_118),
.A2(n_125),
.B1(n_70),
.B2(n_127),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_118),
.B(n_109),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_185),
.Y(n_215)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_118),
.B(n_126),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_171),
.B(n_184),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_78),
.B(n_114),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_150),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_172),
.B(n_176),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_114),
.C(n_31),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_192),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_136),
.B1(n_124),
.B2(n_123),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_113),
.B1(n_111),
.B2(n_66),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_34),
.B(n_31),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_63),
.B1(n_37),
.B2(n_35),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_194),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_152),
.A2(n_35),
.B1(n_34),
.B2(n_31),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_0),
.C(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_161),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_141),
.A2(n_166),
.B1(n_140),
.B2(n_142),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_143),
.B1(n_14),
.B2(n_17),
.Y(n_201)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_151),
.B(n_156),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_0),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_200),
.B(n_206),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_192),
.B(n_199),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_143),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_207),
.C(n_219),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_180),
.B(n_147),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_178),
.B(n_171),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_198),
.A2(n_163),
.B1(n_146),
.B2(n_162),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_227),
.B1(n_228),
.B2(n_186),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_182),
.B(n_160),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_168),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_221),
.B(n_222),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_15),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_195),
.C(n_189),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_0),
.B(n_3),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_4),
.B(n_5),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_224),
.A2(n_181),
.B(n_5),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_181),
.B(n_9),
.Y(n_226)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_183),
.A2(n_169),
.B1(n_170),
.B2(n_175),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_193),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_230),
.A2(n_248),
.B1(n_211),
.B2(n_214),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_231),
.A2(n_237),
.B(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_175),
.B1(n_196),
.B2(n_177),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_233),
.A2(n_213),
.B1(n_228),
.B2(n_211),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_190),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_244),
.C(n_255),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_227),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_253),
.Y(n_257)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_243),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_187),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_245),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_196),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

XOR2x1_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_201),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_4),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_197),
.C(n_6),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_8),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_219),
.C(n_220),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_254),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_275),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_216),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_270),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_234),
.B(n_225),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_225),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_256),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_235),
.A2(n_221),
.B(n_224),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

XOR2x1_ASAP7_75t_SL g292 ( 
.A(n_274),
.B(n_223),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_217),
.C(n_204),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_223),
.C(n_6),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_251),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_246),
.B1(n_243),
.B2(n_245),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_285),
.B1(n_292),
.B2(n_253),
.Y(n_299)
);

AOI21x1_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_233),
.B(n_249),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_286),
.A2(n_271),
.B1(n_270),
.B2(n_242),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_262),
.B(n_249),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_295),
.B(n_236),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_241),
.Y(n_309)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_261),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_250),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_264),
.A2(n_247),
.B(n_238),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_275),
.C(n_258),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_300),
.Y(n_322)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_258),
.C(n_257),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_257),
.C(n_278),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_291),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_269),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_265),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_307),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_306),
.B(n_280),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_310),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_268),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_311),
.A2(n_288),
.B1(n_290),
.B2(n_281),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_255),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_314),
.B(n_300),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_283),
.Y(n_317)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_292),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_321),
.B(n_325),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_298),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_296),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_328),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_305),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_315),
.A2(n_311),
.B(n_302),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_334),
.C(n_324),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_297),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_320),
.B(n_313),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_335),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_307),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_8),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_11),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_322),
.C(n_321),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_341),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_325),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_327),
.A2(n_318),
.B(n_12),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_342),
.B(n_8),
.Y(n_344)
);

AND2x2_ASAP7_75t_SL g343 ( 
.A(n_337),
.B(n_327),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_343),
.B(n_344),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_346),
.B(n_338),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_345),
.C(n_336),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_347),
.B(n_11),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_4),
.C(n_6),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_351),
.A2(n_11),
.B(n_12),
.Y(n_352)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_352),
.Y(n_353)
);


endmodule