module real_jpeg_29044_n_13 (n_46, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_47, n_2, n_45, n_6, n_7, n_3, n_10, n_9, n_13);

input n_46;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_47;
input n_2;
input n_45;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_33;
wire n_29;
wire n_31;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_14;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;

NAND3xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_3),
.C(n_16),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_3),
.B(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_16),
.C(n_47),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_7),
.B(n_16),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_L g39 ( 
.A(n_5),
.B(n_7),
.C(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_12),
.B(n_16),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g33 ( 
.A(n_8),
.B(n_12),
.C(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_9),
.A2(n_28),
.B(n_29),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_35),
.B(n_36),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_35),
.C(n_36),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_9),
.A2(n_41),
.B(n_42),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_9),
.B(n_41),
.C(n_42),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_19),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_17),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_45),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_40),
.B(n_43),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_38),
.B(n_39),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_34),
.B(n_37),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_32),
.B(n_33),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B(n_30),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_46),
.Y(n_28)
);


endmodule