module fake_ariane_82_n_1009 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1009);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1009;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_821;
wire n_218;
wire n_770;
wire n_839;
wire n_928;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_939;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_976;
wire n_909;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_0),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_7),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_102),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_51),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_76),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_74),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_27),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_44),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_18),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_33),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_62),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_48),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_169),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_101),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_118),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_72),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_185),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_46),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_59),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_138),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_129),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_172),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_199),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_113),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_156),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_45),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_89),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_83),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_106),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_31),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_91),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_124),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_75),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_26),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_31),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_150),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_88),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_182),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_116),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_195),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_144),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_174),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_63),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_5),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_103),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_41),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_21),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_146),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_114),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_177),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_160),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_167),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_69),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_24),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_123),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_100),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_154),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_186),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_119),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_165),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_115),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_52),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_32),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_71),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_140),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_135),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_137),
.Y(n_281)
);

BUFx2_ASAP7_75t_SL g282 ( 
.A(n_159),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_6),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_134),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_60),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_20),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_90),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_9),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_58),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_197),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_25),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_180),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_0),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_194),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_201),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_14),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_259),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_206),
.B(n_1),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_220),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_227),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_207),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_253),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_273),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_274),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_216),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_245),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_R g319 ( 
.A(n_249),
.B(n_38),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_205),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_297),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_212),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_215),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_242),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_210),
.B(n_1),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_246),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_247),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_267),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_291),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_286),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_213),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_2),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_219),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_221),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_294),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_295),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_240),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_241),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_243),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_220),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_244),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_208),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_263),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_265),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_209),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_211),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_217),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_218),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_222),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_224),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_303),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_307),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_309),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_214),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_310),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_311),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_341),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_315),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_298),
.B(n_276),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_304),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_328),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_299),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_R g372 ( 
.A(n_348),
.B(n_296),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_332),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_343),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_334),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_343),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_299),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_349),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_305),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_287),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_320),
.B(n_282),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_321),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_335),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_290),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_337),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_347),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_301),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_345),
.B(n_223),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_322),
.B(n_223),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_347),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_350),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_330),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_350),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_317),
.B(n_225),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_351),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_324),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_356),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_358),
.B(n_326),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_318),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_397),
.B(n_226),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_356),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_369),
.B(n_331),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_394),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_363),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_364),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_364),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_363),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_354),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_371),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_351),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_354),
.Y(n_430)
);

OR2x6_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_226),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_327),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_386),
.Y(n_433)
);

AND2x2_ASAP7_75t_SL g434 ( 
.A(n_395),
.B(n_268),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_394),
.B(n_327),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_333),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

INVx4_ASAP7_75t_SL g438 ( 
.A(n_394),
.Y(n_438)
);

NOR2x1p5_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_336),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_359),
.Y(n_440)
);

OR2x6_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_268),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_394),
.B(n_398),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_394),
.B(n_336),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_375),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_373),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_404),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_373),
.B(n_278),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_398),
.B(n_228),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_373),
.B(n_321),
.Y(n_451)
);

OAI22xp33_ASAP7_75t_L g452 ( 
.A1(n_353),
.A2(n_270),
.B1(n_278),
.B2(n_269),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_365),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_355),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_393),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_366),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_389),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_391),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_398),
.B(n_260),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

INVx4_ASAP7_75t_SL g466 ( 
.A(n_395),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_383),
.A2(n_292),
.B1(n_285),
.B2(n_284),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_398),
.B(n_260),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_368),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_355),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_357),
.A2(n_281),
.B1(n_280),
.B2(n_279),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_357),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_360),
.B(n_275),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_410),
.B(n_2),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_360),
.Y(n_479)
);

NAND3x1_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_3),
.C(n_4),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_362),
.Y(n_481)
);

BUFx4f_ASAP7_75t_L g482 ( 
.A(n_372),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_362),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_367),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_367),
.B(n_229),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_448),
.B(n_230),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_231),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_447),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_425),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_434),
.A2(n_370),
.B1(n_406),
.B2(n_380),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_432),
.B(n_232),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_482),
.B(n_407),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_481),
.B(n_374),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_437),
.A2(n_234),
.B(n_233),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_412),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_413),
.B(n_374),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_432),
.B(n_235),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_434),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_437),
.A2(n_237),
.B(n_236),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

BUFx8_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_415),
.B(n_238),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_415),
.A2(n_403),
.B1(n_400),
.B2(n_399),
.Y(n_505)
);

O2A1O1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_445),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_482),
.B(n_220),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_453),
.B(n_239),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_6),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_482),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_466),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_453),
.B(n_248),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_453),
.B(n_252),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_447),
.B(n_254),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_466),
.B(n_376),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_417),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_447),
.B(n_255),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_455),
.B(n_220),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_455),
.B(n_261),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_L g522 ( 
.A(n_476),
.B(n_376),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_444),
.A2(n_403),
.B1(n_400),
.B2(n_399),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_455),
.B(n_262),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_466),
.B(n_390),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_456),
.B(n_264),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_444),
.A2(n_390),
.B1(n_260),
.B2(n_220),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_431),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_431),
.B(n_371),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_456),
.B(n_271),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_459),
.B(n_272),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_445),
.B(n_8),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_451),
.Y(n_534)
);

CKINVDCx6p67_ASAP7_75t_R g535 ( 
.A(n_481),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_421),
.A2(n_258),
.B(n_220),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_460),
.B(n_258),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_428),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_454),
.B(n_377),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_459),
.B(n_258),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_422),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_431),
.B(n_476),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_468),
.B(n_258),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_469),
.B(n_9),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_468),
.B(n_258),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_R g546 ( 
.A(n_476),
.B(n_377),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_446),
.A2(n_260),
.B1(n_258),
.B2(n_384),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_460),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_441),
.A2(n_384),
.B1(n_11),
.B2(n_12),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_419),
.B(n_10),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_419),
.B(n_10),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_446),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_426),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_441),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_414),
.B(n_15),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_423),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_423),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_418),
.B(n_16),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_458),
.B(n_16),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_469),
.B(n_17),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_460),
.B(n_17),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_460),
.B(n_18),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_469),
.B(n_19),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_438),
.B(n_479),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_440),
.B(n_19),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_485),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_442),
.B(n_20),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_430),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_457),
.B(n_21),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_477),
.B(n_22),
.C(n_23),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_430),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_510),
.A2(n_449),
.B(n_443),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_496),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_507),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_512),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_520),
.A2(n_424),
.B(n_411),
.Y(n_576)
);

BUFx8_ASAP7_75t_L g577 ( 
.A(n_529),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_499),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_542),
.B(n_479),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_499),
.B(n_449),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_494),
.B(n_431),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_497),
.B(n_436),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_490),
.Y(n_583)
);

NAND2x1p5_ASAP7_75t_L g584 ( 
.A(n_512),
.B(n_528),
.Y(n_584)
);

A2O1A1Ixp33_ASAP7_75t_L g585 ( 
.A1(n_532),
.A2(n_477),
.B(n_484),
.C(n_483),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_501),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_503),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_542),
.B(n_478),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_516),
.B(n_525),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_553),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_547),
.A2(n_441),
.B1(n_452),
.B2(n_478),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_511),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_516),
.B(n_485),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_532),
.A2(n_441),
.B1(n_480),
.B2(n_478),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_538),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_546),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_517),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_539),
.B(n_429),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_534),
.B(n_472),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_546),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_511),
.B(n_485),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_535),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_528),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_568),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_510),
.B(n_461),
.Y(n_605)
);

BUFx12f_ASAP7_75t_L g606 ( 
.A(n_502),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_548),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_489),
.B(n_462),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_547),
.A2(n_463),
.B1(n_470),
.B2(n_465),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_554),
.A2(n_480),
.B1(n_438),
.B2(n_420),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_489),
.B(n_474),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_502),
.B(n_428),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_525),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_534),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_494),
.B(n_529),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_571),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_494),
.Y(n_617)
);

NOR2x1_ASAP7_75t_L g618 ( 
.A(n_493),
.B(n_439),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_518),
.Y(n_619)
);

BUFx12f_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_491),
.B(n_485),
.Y(n_621)
);

BUFx4f_ASAP7_75t_SL g622 ( 
.A(n_493),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_533),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_SL g624 ( 
.A(n_570),
.B(n_486),
.C(n_475),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_492),
.B(n_438),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_504),
.A2(n_416),
.B1(n_433),
.B2(n_485),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_498),
.B(n_467),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_548),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_558),
.B(n_424),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_541),
.B(n_424),
.Y(n_630)
);

CKINVDCx6p67_ASAP7_75t_R g631 ( 
.A(n_565),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_556),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_557),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_566),
.B(n_474),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_522),
.B(n_411),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_567),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_491),
.B(n_464),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_576),
.A2(n_536),
.B(n_537),
.Y(n_638)
);

NOR2x1_ASAP7_75t_L g639 ( 
.A(n_603),
.B(n_564),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_580),
.B(n_555),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_625),
.A2(n_537),
.B(n_540),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_575),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_625),
.A2(n_545),
.B(n_543),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_583),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_595),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_572),
.A2(n_520),
.B(n_508),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_603),
.B(n_564),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_586),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_630),
.A2(n_551),
.B(n_550),
.Y(n_649)
);

OAI21x1_ASAP7_75t_SL g650 ( 
.A1(n_605),
.A2(n_554),
.B(n_569),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_589),
.B(n_505),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_572),
.A2(n_544),
.B(n_560),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_602),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_605),
.A2(n_508),
.B(n_515),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_630),
.A2(n_563),
.B(n_562),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_608),
.A2(n_629),
.B(n_601),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_627),
.A2(n_521),
.B(n_519),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_585),
.A2(n_524),
.B(n_544),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_581),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_580),
.B(n_527),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_614),
.A2(n_506),
.B(n_561),
.C(n_562),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_606),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_592),
.B(n_561),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_612),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_584),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_577),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_608),
.A2(n_474),
.B(n_495),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_581),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_587),
.A2(n_500),
.B(n_464),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_590),
.A2(n_513),
.B(n_509),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_610),
.A2(n_552),
.B(n_549),
.C(n_527),
.Y(n_671)
);

NAND2x1_ASAP7_75t_L g672 ( 
.A(n_611),
.B(n_427),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_593),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_610),
.A2(n_624),
.B(n_594),
.C(n_552),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_636),
.B(n_613),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_573),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_L g677 ( 
.A1(n_594),
.A2(n_523),
.B1(n_487),
.B2(n_488),
.Y(n_677)
);

OA21x2_ASAP7_75t_L g678 ( 
.A1(n_604),
.A2(n_514),
.B(n_526),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_574),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_584),
.Y(n_680)
);

OAI21x1_ASAP7_75t_L g681 ( 
.A1(n_616),
.A2(n_531),
.B(n_530),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_607),
.B(n_427),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_632),
.A2(n_450),
.B(n_427),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_599),
.B(n_598),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_597),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_591),
.A2(n_523),
.B1(n_23),
.B2(n_24),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_635),
.A2(n_471),
.B(n_22),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_619),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_578),
.B(n_471),
.Y(n_689)
);

NOR2x1_ASAP7_75t_SL g690 ( 
.A(n_581),
.B(n_471),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_623),
.A2(n_471),
.B(n_40),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_657),
.A2(n_635),
.B(n_579),
.Y(n_692)
);

AO32x2_ASAP7_75t_L g693 ( 
.A1(n_686),
.A2(n_617),
.A3(n_637),
.B1(n_621),
.B2(n_631),
.Y(n_693)
);

AOI21xp33_ASAP7_75t_L g694 ( 
.A1(n_677),
.A2(n_626),
.B(n_609),
.Y(n_694)
);

OA21x2_ASAP7_75t_L g695 ( 
.A1(n_658),
.A2(n_633),
.B(n_634),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_652),
.B(n_588),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_644),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_643),
.A2(n_634),
.B(n_618),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_677),
.A2(n_582),
.B(n_596),
.C(n_600),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_673),
.B(n_589),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_648),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_685),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_680),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_686),
.A2(n_620),
.B1(n_588),
.B2(n_577),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_688),
.Y(n_705)
);

OA21x2_ASAP7_75t_L g706 ( 
.A1(n_658),
.A2(n_593),
.B(n_611),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_651),
.A2(n_588),
.B1(n_615),
.B2(n_622),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_683),
.A2(n_611),
.B(n_607),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_649),
.A2(n_611),
.B(n_607),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_674),
.B(n_615),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_676),
.Y(n_711)
);

OA21x2_ASAP7_75t_L g712 ( 
.A1(n_652),
.A2(n_628),
.B(n_471),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_679),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_657),
.A2(n_628),
.B(n_615),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_655),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_684),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_645),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_667),
.A2(n_628),
.B(n_592),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_674),
.A2(n_592),
.B1(n_588),
.B2(n_27),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_659),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_673),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_640),
.B(n_471),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_670),
.A2(n_131),
.B(n_203),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_668),
.Y(n_724)
);

BUFx2_ASAP7_75t_R g725 ( 
.A(n_664),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_675),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_680),
.Y(n_727)
);

OA21x2_ASAP7_75t_L g728 ( 
.A1(n_681),
.A2(n_130),
.B(n_202),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_638),
.A2(n_128),
.B(n_200),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_672),
.Y(n_730)
);

BUFx2_ASAP7_75t_SL g731 ( 
.A(n_666),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_669),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_651),
.Y(n_733)
);

AO31x2_ASAP7_75t_L g734 ( 
.A1(n_646),
.A2(n_25),
.A3(n_26),
.B(n_28),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_656),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_653),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_640),
.A2(n_132),
.B(n_198),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_642),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_671),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_663),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_665),
.B(n_29),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_665),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_SL g743 ( 
.A1(n_660),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_696),
.A2(n_654),
.B(n_646),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_716),
.B(n_660),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_717),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_697),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_699),
.B(n_707),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_719),
.A2(n_671),
.B1(n_663),
.B2(n_687),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_733),
.B(n_662),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_701),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_702),
.Y(n_752)
);

CKINVDCx16_ASAP7_75t_R g753 ( 
.A(n_736),
.Y(n_753)
);

AOI21x1_ASAP7_75t_L g754 ( 
.A1(n_714),
.A2(n_654),
.B(n_678),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_694),
.A2(n_661),
.B(n_687),
.C(n_647),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_710),
.B(n_647),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_720),
.B(n_678),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_736),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_710),
.B(n_661),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_739),
.A2(n_650),
.B1(n_690),
.B2(n_689),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_704),
.A2(n_639),
.B1(n_642),
.B2(n_682),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_713),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_727),
.B(n_700),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_724),
.B(n_682),
.Y(n_764)
);

AO31x2_ASAP7_75t_L g765 ( 
.A1(n_732),
.A2(n_689),
.A3(n_641),
.B(n_691),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_721),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_766)
);

NAND3x1_ASAP7_75t_L g767 ( 
.A(n_726),
.B(n_34),
.C(n_35),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_725),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_740),
.B(n_36),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_713),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_770)
);

CKINVDCx11_ASAP7_75t_R g771 ( 
.A(n_703),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_727),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_705),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_703),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_731),
.B(n_37),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_696),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_700),
.B(n_50),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_711),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_741),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_742),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_700),
.B(n_56),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_743),
.A2(n_57),
.B1(n_61),
.B2(n_64),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_703),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_734),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_734),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_703),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_SL g787 ( 
.A1(n_693),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_734),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_721),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_695),
.A2(n_68),
.B(n_70),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_695),
.A2(n_73),
.B(n_77),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_734),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_734),
.Y(n_794)
);

AOI221xp5_ASAP7_75t_L g795 ( 
.A1(n_737),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_703),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_SL g797 ( 
.A(n_721),
.B(n_738),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_742),
.Y(n_798)
);

INVx1_ASAP7_75t_SL g799 ( 
.A(n_740),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_748),
.A2(n_692),
.B1(n_722),
.B2(n_706),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_759),
.B(n_706),
.Y(n_801)
);

OAI221xp5_ASAP7_75t_L g802 ( 
.A1(n_782),
.A2(n_728),
.B1(n_706),
.B2(n_738),
.C(n_732),
.Y(n_802)
);

OAI221xp5_ASAP7_75t_SL g803 ( 
.A1(n_759),
.A2(n_755),
.B1(n_749),
.B2(n_775),
.C(n_795),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_747),
.Y(n_804)
);

AOI222xp33_ASAP7_75t_L g805 ( 
.A1(n_766),
.A2(n_693),
.B1(n_723),
.B2(n_729),
.C1(n_698),
.C2(n_715),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_778),
.A2(n_693),
.B1(n_712),
.B2(n_695),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_784),
.B(n_785),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_795),
.A2(n_723),
.B(n_693),
.C(n_729),
.Y(n_808)
);

AOI221xp5_ASAP7_75t_L g809 ( 
.A1(n_787),
.A2(n_693),
.B1(n_715),
.B2(n_735),
.C(n_730),
.Y(n_809)
);

AO21x2_ASAP7_75t_L g810 ( 
.A1(n_788),
.A2(n_718),
.B(n_735),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_756),
.A2(n_712),
.B1(n_698),
.B2(n_728),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_766),
.A2(n_712),
.B1(n_728),
.B2(n_730),
.Y(n_812)
);

OAI33xp33_ASAP7_75t_L g813 ( 
.A1(n_769),
.A2(n_82),
.A3(n_84),
.B1(n_85),
.B2(n_86),
.B3(n_87),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_751),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_767),
.A2(n_730),
.B1(n_709),
.B2(n_718),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_752),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_773),
.Y(n_817)
);

AOI21xp33_ASAP7_75t_L g818 ( 
.A1(n_793),
.A2(n_709),
.B(n_708),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_761),
.A2(n_708),
.B1(n_93),
.B2(n_94),
.Y(n_819)
);

AOI221xp5_ASAP7_75t_L g820 ( 
.A1(n_794),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.C(n_98),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_757),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_745),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_754),
.A2(n_111),
.B(n_112),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_762),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_790),
.A2(n_117),
.B(n_120),
.C(n_121),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_765),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_746),
.B(n_122),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_772),
.Y(n_828)
);

OAI211xp5_ASAP7_75t_L g829 ( 
.A1(n_744),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_765),
.Y(n_830)
);

AO21x2_ASAP7_75t_L g831 ( 
.A1(n_790),
.A2(n_792),
.B(n_744),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_764),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_792),
.A2(n_133),
.B(n_136),
.C(n_139),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_765),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_780),
.B(n_141),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_799),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_760),
.A2(n_142),
.B1(n_145),
.B2(n_147),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_783),
.B(n_148),
.Y(n_838)
);

AOI221xp5_ASAP7_75t_L g839 ( 
.A1(n_779),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.C(n_155),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_799),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_796),
.Y(n_841)
);

AO21x2_ASAP7_75t_L g842 ( 
.A1(n_776),
.A2(n_157),
.B(n_161),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_798),
.B(n_162),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_758),
.B(n_163),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_760),
.A2(n_164),
.B1(n_168),
.B2(n_170),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_832),
.B(n_753),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_831),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_803),
.A2(n_791),
.B(n_781),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_826),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_801),
.B(n_769),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_801),
.B(n_750),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_807),
.B(n_841),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_830),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_836),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_807),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_830),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_828),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_804),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_840),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_834),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_814),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_834),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_816),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_810),
.B(n_786),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_842),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_817),
.B(n_774),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_810),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_810),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_806),
.B(n_763),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_831),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_824),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_815),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_809),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_831),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_818),
.Y(n_875)
);

BUFx5_ASAP7_75t_L g876 ( 
.A(n_808),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_805),
.B(n_763),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_812),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_808),
.B(n_771),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_843),
.B(n_789),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_823),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_879),
.B(n_843),
.Y(n_882)
);

NOR2x1_ASAP7_75t_L g883 ( 
.A(n_850),
.B(n_835),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_861),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_850),
.B(n_859),
.Y(n_885)
);

OAI22xp33_ASAP7_75t_L g886 ( 
.A1(n_873),
.A2(n_819),
.B1(n_802),
.B2(n_827),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_858),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_858),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_R g889 ( 
.A(n_879),
.B(n_768),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_854),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_866),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_866),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_SL g893 ( 
.A1(n_873),
.A2(n_845),
.B1(n_837),
.B2(n_821),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_872),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_852),
.Y(n_895)
);

AOI33xp33_ASAP7_75t_L g896 ( 
.A1(n_878),
.A2(n_844),
.A3(n_800),
.B1(n_770),
.B2(n_839),
.B3(n_822),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_857),
.B(n_855),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_863),
.Y(n_898)
);

AOI221xp5_ASAP7_75t_L g899 ( 
.A1(n_878),
.A2(n_813),
.B1(n_833),
.B2(n_825),
.C(n_820),
.Y(n_899)
);

AOI221xp5_ASAP7_75t_L g900 ( 
.A1(n_848),
.A2(n_833),
.B1(n_825),
.B2(n_844),
.C(n_829),
.Y(n_900)
);

AOI21xp33_ASAP7_75t_L g901 ( 
.A1(n_875),
.A2(n_842),
.B(n_838),
.Y(n_901)
);

CKINVDCx16_ASAP7_75t_R g902 ( 
.A(n_851),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_863),
.Y(n_903)
);

OAI211xp5_ASAP7_75t_L g904 ( 
.A1(n_865),
.A2(n_811),
.B(n_789),
.C(n_777),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_902),
.B(n_876),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_887),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_882),
.B(n_865),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_894),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_895),
.B(n_876),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_888),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_891),
.B(n_876),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_882),
.B(n_875),
.Y(n_912)
);

AND2x2_ASAP7_75t_SL g913 ( 
.A(n_891),
.B(n_865),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_882),
.B(n_864),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_892),
.B(n_897),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_890),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_892),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_885),
.B(n_876),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_885),
.B(n_876),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_898),
.Y(n_920)
);

NAND2x1_ASAP7_75t_SL g921 ( 
.A(n_905),
.B(n_883),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_908),
.B(n_884),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_907),
.A2(n_900),
.B1(n_886),
.B2(n_899),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_906),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_908),
.B(n_903),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_916),
.B(n_855),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_912),
.Y(n_927)
);

INVxp67_ASAP7_75t_SL g928 ( 
.A(n_916),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_906),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_905),
.B(n_851),
.Y(n_930)
);

NOR3xp33_ASAP7_75t_L g931 ( 
.A(n_923),
.B(n_900),
.C(n_893),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_928),
.B(n_912),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_927),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_930),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_922),
.B(n_910),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_924),
.B(n_918),
.Y(n_936)
);

NAND4xp25_ASAP7_75t_SL g937 ( 
.A(n_926),
.B(n_911),
.C(n_919),
.D(n_918),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_929),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_927),
.B(n_912),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_938),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_935),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_932),
.B(n_911),
.Y(n_942)
);

OAI222xp33_ASAP7_75t_L g943 ( 
.A1(n_934),
.A2(n_907),
.B1(n_865),
.B2(n_919),
.C1(n_912),
.C2(n_877),
.Y(n_943)
);

AOI221xp5_ASAP7_75t_L g944 ( 
.A1(n_940),
.A2(n_931),
.B1(n_901),
.B2(n_936),
.C(n_937),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_941),
.B(n_936),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_940),
.B(n_932),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_942),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_R g948 ( 
.A(n_946),
.B(n_889),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_944),
.A2(n_943),
.B(n_933),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_947),
.B(n_942),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_945),
.B(n_925),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_945),
.Y(n_952)
);

NAND4xp25_ASAP7_75t_L g953 ( 
.A(n_950),
.B(n_939),
.C(n_917),
.D(n_911),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_952),
.B(n_951),
.Y(n_954)
);

OAI321xp33_ASAP7_75t_L g955 ( 
.A1(n_949),
.A2(n_907),
.A3(n_904),
.B1(n_877),
.B2(n_867),
.C(n_876),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_948),
.B(n_917),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_952),
.B(n_917),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_SL g958 ( 
.A(n_949),
.B(n_896),
.C(n_915),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_950),
.B(n_915),
.Y(n_959)
);

NAND5xp2_ASAP7_75t_L g960 ( 
.A(n_949),
.B(n_880),
.C(n_901),
.D(n_913),
.E(n_909),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_951),
.Y(n_961)
);

AOI321xp33_ASAP7_75t_L g962 ( 
.A1(n_955),
.A2(n_864),
.A3(n_846),
.B1(n_914),
.B2(n_876),
.C(n_869),
.Y(n_962)
);

O2A1O1Ixp5_ASAP7_75t_L g963 ( 
.A1(n_956),
.A2(n_917),
.B(n_920),
.C(n_914),
.Y(n_963)
);

OAI211xp5_ASAP7_75t_SL g964 ( 
.A1(n_961),
.A2(n_910),
.B(n_870),
.C(n_874),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_L g965 ( 
.A(n_954),
.B(n_957),
.C(n_953),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_959),
.A2(n_907),
.B1(n_913),
.B2(n_914),
.Y(n_966)
);

NAND2x1_ASAP7_75t_SL g967 ( 
.A(n_958),
.B(n_914),
.Y(n_967)
);

AOI221xp5_ASAP7_75t_SL g968 ( 
.A1(n_960),
.A2(n_920),
.B1(n_847),
.B2(n_870),
.C(n_874),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_961),
.B(n_907),
.C(n_913),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_965),
.B(n_781),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_967),
.Y(n_971)
);

AOI211xp5_ASAP7_75t_L g972 ( 
.A1(n_969),
.A2(n_797),
.B(n_920),
.C(n_909),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_963),
.Y(n_973)
);

NAND2xp33_ASAP7_75t_R g974 ( 
.A(n_962),
.B(n_907),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_966),
.Y(n_975)
);

NAND3xp33_ASAP7_75t_SL g976 ( 
.A(n_968),
.B(n_909),
.C(n_921),
.Y(n_976)
);

OAI322xp33_ASAP7_75t_L g977 ( 
.A1(n_964),
.A2(n_847),
.A3(n_874),
.B1(n_870),
.B2(n_876),
.C1(n_881),
.C2(n_867),
.Y(n_977)
);

AOI221xp5_ASAP7_75t_L g978 ( 
.A1(n_968),
.A2(n_874),
.B1(n_847),
.B2(n_870),
.C(n_881),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_968),
.A2(n_876),
.B1(n_842),
.B2(n_847),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_973),
.B(n_852),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_971),
.Y(n_981)
);

NAND4xp75_ASAP7_75t_L g982 ( 
.A(n_979),
.B(n_838),
.C(n_869),
.D(n_871),
.Y(n_982)
);

AND3x4_ASAP7_75t_L g983 ( 
.A(n_970),
.B(n_975),
.C(n_972),
.Y(n_983)
);

NAND4xp25_ASAP7_75t_L g984 ( 
.A(n_974),
.B(n_881),
.C(n_864),
.D(n_852),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_976),
.B(n_977),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_SL g986 ( 
.A(n_978),
.B(n_868),
.C(n_871),
.Y(n_986)
);

AND3x4_ASAP7_75t_L g987 ( 
.A(n_970),
.B(n_864),
.C(n_852),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_971),
.A2(n_868),
.B1(n_862),
.B2(n_860),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_983),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_986),
.A2(n_868),
.B1(n_862),
.B2(n_860),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_981),
.B(n_862),
.C(n_860),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_985),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_980),
.A2(n_856),
.B(n_853),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_987),
.Y(n_994)
);

XNOR2xp5_ASAP7_75t_L g995 ( 
.A(n_984),
.B(n_171),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_989),
.B(n_982),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_992),
.Y(n_997)
);

NAND4xp25_ASAP7_75t_L g998 ( 
.A(n_994),
.B(n_988),
.C(n_175),
.D(n_176),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_995),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_997),
.B(n_991),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_996),
.A2(n_993),
.B(n_990),
.Y(n_1001)
);

OAI22x1_ASAP7_75t_L g1002 ( 
.A1(n_999),
.A2(n_856),
.B1(n_853),
.B2(n_849),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_1000),
.A2(n_996),
.B1(n_998),
.B2(n_856),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_1003),
.Y(n_1004)
);

OAI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_1004),
.A2(n_1001),
.B1(n_1002),
.B2(n_853),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_1005),
.A2(n_178),
.B(n_179),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_SL g1007 ( 
.A1(n_1006),
.A2(n_181),
.B1(n_183),
.B2(n_184),
.Y(n_1007)
);

OAI221xp5_ASAP7_75t_R g1008 ( 
.A1(n_1007),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.C(n_190),
.Y(n_1008)
);

AOI211xp5_ASAP7_75t_L g1009 ( 
.A1(n_1008),
.A2(n_191),
.B(n_192),
.C(n_193),
.Y(n_1009)
);


endmodule