module fake_jpeg_17897_n_275 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_54),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_34),
.C(n_31),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_16),
.B(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_24),
.B1(n_34),
.B2(n_31),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_64),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_5),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_100),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_72),
.A2(n_88),
.B(n_11),
.Y(n_141)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_78),
.B(n_83),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_22),
.B1(n_37),
.B2(n_24),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_59),
.B1(n_30),
.B2(n_26),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_19),
.Y(n_87)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_27),
.B1(n_37),
.B2(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_36),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_95),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_90),
.A2(n_13),
.B(n_68),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_18),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_18),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_101),
.Y(n_137)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_43),
.B(n_33),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_33),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_30),
.C(n_53),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_26),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_27),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_9),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_108),
.B(n_121),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_109),
.B(n_125),
.Y(n_171)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_131),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_80),
.B1(n_93),
.B2(n_94),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_118),
.B(n_136),
.Y(n_175)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_26),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_8),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_138),
.Y(n_163)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_124),
.A2(n_99),
.B1(n_91),
.B2(n_82),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_102),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_141),
.B(n_122),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_66),
.B(n_9),
.Y(n_132)
);

CKINVDCx12_ASAP7_75t_R g133 ( 
.A(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_135),
.Y(n_167)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_73),
.B(n_11),
.Y(n_138)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_11),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_67),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_132),
.C(n_140),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_145),
.B(n_142),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_74),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_98),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_107),
.B(n_77),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_152),
.B(n_164),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_136),
.A2(n_73),
.B(n_76),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_160),
.B(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_156),
.B(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_109),
.A2(n_91),
.B1(n_82),
.B2(n_76),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_161),
.B1(n_129),
.B2(n_116),
.Y(n_185)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_159),
.A2(n_116),
.B1(n_123),
.B2(n_111),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_80),
.B(n_99),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_93),
.B1(n_96),
.B2(n_118),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_173),
.B1(n_137),
.B2(n_129),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_121),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_117),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_108),
.B(n_115),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_134),
.B1(n_124),
.B2(n_127),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_178),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_185),
.A2(n_191),
.B1(n_153),
.B2(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_145),
.B(n_163),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_174),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_196),
.Y(n_203)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_112),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_170),
.Y(n_197)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_150),
.A2(n_110),
.B1(n_139),
.B2(n_135),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_198),
.A2(n_159),
.B1(n_168),
.B2(n_171),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_114),
.C(n_110),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_200),
.C(n_154),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_119),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_202),
.A2(n_213),
.B1(n_215),
.B2(n_183),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_207),
.C(n_211),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_154),
.C(n_149),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_166),
.C(n_169),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_152),
.B(n_159),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_146),
.Y(n_216)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_164),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_184),
.C(n_178),
.Y(n_238)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_208),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_230),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_195),
.B1(n_182),
.B2(n_177),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_224),
.A2(n_232),
.B1(n_233),
.B2(n_212),
.Y(n_245)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_183),
.B1(n_191),
.B2(n_182),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_221),
.B1(n_177),
.B2(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_196),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_236),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_184),
.C(n_199),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_215),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_204),
.C(n_207),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_202),
.B1(n_203),
.B2(n_211),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_245),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_229),
.C(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_243),
.C(n_241),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_218),
.B(n_212),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_248),
.B(n_227),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_163),
.B(n_209),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_226),
.B(n_242),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_249),
.B(n_227),
.Y(n_251)
);

OAI31xp33_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_253),
.A3(n_198),
.B(n_181),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_229),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_256),
.Y(n_264)
);

OA21x2_ASAP7_75t_SL g253 ( 
.A1(n_244),
.A2(n_238),
.B(n_237),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_258),
.C(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_235),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_156),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_224),
.C(n_228),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_262),
.C(n_256),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_265),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_263),
.A3(n_260),
.B1(n_223),
.B2(n_186),
.C1(n_228),
.C2(n_259),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_258),
.A2(n_242),
.B(n_226),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_268),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_214),
.A3(n_219),
.B1(n_179),
.B2(n_167),
.C1(n_119),
.C2(n_165),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_214),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_270),
.B(n_165),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_147),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_272),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_273),
.Y(n_275)
);


endmodule