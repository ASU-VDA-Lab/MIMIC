module real_aes_8831_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g519 ( .A1(n_0), .A2(n_166), .B(n_520), .C(n_523), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_1), .B(n_515), .Y(n_524) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g164 ( .A(n_3), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_4), .B(n_167), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_5), .A2(n_484), .B(n_559), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_6), .A2(n_768), .B1(n_771), .B2(n_772), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_6), .Y(n_772) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_7), .A2(n_174), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_8), .A2(n_37), .B1(n_154), .B2(n_202), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_9), .B(n_174), .Y(n_182) );
AND2x6_ASAP7_75t_L g169 ( .A(n_10), .B(n_170), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_11), .A2(n_169), .B(n_489), .C(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_12), .A2(n_41), .B1(n_769), .B2(n_770), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_12), .Y(n_769) );
INVx1_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_13), .B(n_38), .Y(n_464) );
INVx1_ASAP7_75t_L g148 ( .A(n_14), .Y(n_148) );
INVx1_ASAP7_75t_L g145 ( .A(n_15), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_16), .B(n_150), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_17), .B(n_167), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_18), .B(n_141), .Y(n_248) );
AO32x2_ASAP7_75t_L g218 ( .A1(n_19), .A2(n_140), .A3(n_174), .B1(n_193), .B2(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_20), .B(n_154), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_21), .B(n_141), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_22), .A2(n_57), .B1(n_154), .B2(n_202), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_23), .A2(n_85), .B1(n_150), .B2(n_154), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_24), .B(n_154), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_25), .A2(n_193), .B(n_489), .C(n_507), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_26), .A2(n_193), .B(n_489), .C(n_541), .Y(n_540) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_27), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_28), .B(n_195), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_29), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_29), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_30), .A2(n_484), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_31), .B(n_195), .Y(n_236) );
INVx2_ASAP7_75t_L g152 ( .A(n_32), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_33), .A2(n_487), .B(n_491), .C(n_497), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_34), .B(n_154), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_35), .B(n_195), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_36), .B(n_213), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_38), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_39), .B(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_40), .Y(n_536) );
INVx1_ASAP7_75t_L g770 ( .A(n_41), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_42), .B(n_167), .Y(n_553) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_43), .A2(n_452), .B1(n_455), .B2(n_456), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_43), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_44), .B(n_484), .Y(n_539) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_45), .A2(n_47), .B1(n_453), .B2(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_45), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g471 ( .A1(n_45), .A2(n_128), .B1(n_129), .B2(n_454), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_46), .A2(n_487), .B(n_497), .C(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_47), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_48), .B(n_154), .Y(n_177) );
INVx1_ASAP7_75t_L g521 ( .A(n_49), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_50), .A2(n_94), .B1(n_202), .B2(n_203), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_51), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_52), .B(n_154), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_53), .B(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g552 ( .A(n_54), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_55), .B(n_484), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_56), .B(n_162), .Y(n_181) );
AOI22xp33_ASAP7_75t_SL g246 ( .A1(n_58), .A2(n_62), .B1(n_150), .B2(n_154), .Y(n_246) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_59), .A2(n_69), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_59), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_60), .B(n_154), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_61), .B(n_154), .Y(n_210) );
INVx1_ASAP7_75t_L g170 ( .A(n_63), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_64), .B(n_484), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_65), .B(n_515), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_66), .A2(n_156), .B(n_162), .C(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_67), .B(n_154), .Y(n_165) );
INVx1_ASAP7_75t_L g144 ( .A(n_68), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_69), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_70), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_71), .B(n_167), .Y(n_495) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_72), .A2(n_174), .A3(n_193), .B1(n_200), .B2(n_205), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_73), .B(n_168), .Y(n_533) );
INVx1_ASAP7_75t_L g189 ( .A(n_74), .Y(n_189) );
INVx1_ASAP7_75t_L g231 ( .A(n_75), .Y(n_231) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_76), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_77), .B(n_494), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_78), .A2(n_489), .B(n_497), .C(n_586), .Y(n_585) );
AOI222xp33_ASAP7_75t_L g469 ( .A1(n_79), .A2(n_470), .B1(n_763), .B2(n_764), .C1(n_773), .C2(n_777), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_80), .B(n_150), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_81), .A2(n_106), .B1(n_115), .B2(n_782), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g560 ( .A(n_82), .Y(n_560) );
INVx1_ASAP7_75t_L g114 ( .A(n_83), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_84), .B(n_493), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_86), .B(n_202), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_87), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_88), .B(n_150), .Y(n_235) );
INVx2_ASAP7_75t_L g142 ( .A(n_89), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_90), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_91), .B(n_192), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_92), .B(n_150), .Y(n_178) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_93), .B(n_111), .C(n_112), .Y(n_110) );
OR2x2_ASAP7_75t_L g461 ( .A(n_93), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g474 ( .A(n_93), .B(n_463), .Y(n_474) );
INVx2_ASAP7_75t_L g762 ( .A(n_93), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_95), .A2(n_104), .B1(n_150), .B2(n_151), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_96), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g492 ( .A(n_97), .Y(n_492) );
INVxp67_ASAP7_75t_L g563 ( .A(n_98), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_99), .B(n_150), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_100), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g529 ( .A(n_101), .Y(n_529) );
INVx1_ASAP7_75t_L g587 ( .A(n_102), .Y(n_587) );
AND2x2_ASAP7_75t_L g554 ( .A(n_103), .B(n_195), .Y(n_554) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx4f_ASAP7_75t_SL g782 ( .A(n_107), .Y(n_782) );
OR2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g463 ( .A(n_111), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_468), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g781 ( .A(n_119), .Y(n_781) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_458), .B(n_465), .Y(n_121) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_126), .B1(n_127), .B2(n_457), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_123), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_124), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_129), .B1(n_450), .B2(n_451), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_416), .Y(n_129) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_320), .C(n_404), .Y(n_130) );
NAND4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_263), .C(n_285), .D(n_301), .Y(n_131) );
AOI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_196), .B1(n_222), .B2(n_241), .C(n_249), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_172), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_135), .B(n_241), .Y(n_275) );
NAND4xp25_ASAP7_75t_L g315 ( .A(n_135), .B(n_303), .C(n_316), .D(n_318), .Y(n_315) );
INVxp67_ASAP7_75t_L g432 ( .A(n_135), .Y(n_432) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g314 ( .A(n_136), .B(n_252), .Y(n_314) );
AND2x2_ASAP7_75t_L g338 ( .A(n_136), .B(n_172), .Y(n_338) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g305 ( .A(n_137), .B(n_240), .Y(n_305) );
AND2x2_ASAP7_75t_L g345 ( .A(n_137), .B(n_326), .Y(n_345) );
AND2x2_ASAP7_75t_L g362 ( .A(n_137), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_137), .B(n_173), .Y(n_386) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g239 ( .A(n_138), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g257 ( .A(n_138), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g269 ( .A(n_138), .B(n_173), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_138), .B(n_183), .Y(n_291) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_146), .B(n_171), .Y(n_138) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_139), .A2(n_184), .B(n_194), .Y(n_183) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_140), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_142), .B(n_143), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_160), .B(n_169), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_153), .C(n_156), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_149), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_149), .A2(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
INVx1_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
INVx3_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_154), .Y(n_589) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
AND2x6_ASAP7_75t_L g489 ( .A(n_155), .B(n_490), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g586 ( .A1(n_156), .A2(n_587), .B(n_588), .C(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_157), .A2(n_234), .B(n_235), .Y(n_233) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g494 ( .A(n_158), .Y(n_494) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g168 ( .A(n_159), .Y(n_168) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
INVx1_ASAP7_75t_L g213 ( .A(n_159), .Y(n_213) );
AND2x2_ASAP7_75t_L g485 ( .A(n_159), .B(n_163), .Y(n_485) );
INVx1_ASAP7_75t_L g490 ( .A(n_159), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_164), .B(n_165), .C(n_166), .Y(n_160) );
O2A1O1Ixp5_ASAP7_75t_L g188 ( .A1(n_161), .A2(n_189), .B(n_190), .C(n_191), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_161), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_166), .A2(n_180), .B(n_181), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_166), .A2(n_192), .B1(n_220), .B2(n_221), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_166), .A2(n_192), .B1(n_245), .B2(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_167), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_167), .A2(n_186), .B(n_187), .Y(n_185) );
O2A1O1Ixp5_ASAP7_75t_SL g229 ( .A1(n_167), .A2(n_230), .B(n_231), .C(n_232), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_167), .B(n_563), .Y(n_562) );
INVx5_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g200 ( .A1(n_168), .A2(n_192), .B1(n_201), .B2(n_204), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g175 ( .A1(n_169), .A2(n_176), .B(n_179), .Y(n_175) );
BUFx3_ASAP7_75t_L g193 ( .A(n_169), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_169), .A2(n_209), .B(n_214), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_169), .A2(n_229), .B(n_233), .Y(n_228) );
AND2x4_ASAP7_75t_L g484 ( .A(n_169), .B(n_485), .Y(n_484) );
INVx4_ASAP7_75t_SL g498 ( .A(n_169), .Y(n_498) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_169), .B(n_485), .Y(n_530) );
AND2x2_ASAP7_75t_L g272 ( .A(n_172), .B(n_273), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_172), .A2(n_322), .B1(n_325), .B2(n_327), .C(n_331), .Y(n_321) );
AND2x2_ASAP7_75t_L g380 ( .A(n_172), .B(n_345), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_172), .B(n_362), .Y(n_414) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_183), .Y(n_172) );
INVx3_ASAP7_75t_L g240 ( .A(n_173), .Y(n_240) );
AND2x2_ASAP7_75t_L g289 ( .A(n_173), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g343 ( .A(n_173), .B(n_258), .Y(n_343) );
AND2x2_ASAP7_75t_L g401 ( .A(n_173), .B(n_402), .Y(n_401) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_182), .Y(n_173) );
INVx4_ASAP7_75t_L g243 ( .A(n_174), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_174), .A2(n_539), .B(n_540), .Y(n_538) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_174), .Y(n_557) );
AND2x2_ASAP7_75t_L g241 ( .A(n_183), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g313 ( .A(n_183), .Y(n_313) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_183), .Y(n_319) );
AND2x2_ASAP7_75t_L g364 ( .A(n_183), .B(n_240), .Y(n_364) );
OR2x2_ASAP7_75t_L g403 ( .A(n_183), .B(n_242), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_188), .B(n_193), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_191), .A2(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx4_ASAP7_75t_L g522 ( .A(n_192), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g262 ( .A(n_193), .B(n_243), .C(n_244), .Y(n_262) );
INVx2_ASAP7_75t_L g205 ( .A(n_195), .Y(n_205) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_195), .A2(n_208), .B(n_217), .Y(n_207) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_195), .A2(n_228), .B(n_236), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_195), .A2(n_483), .B(n_486), .Y(n_482) );
INVx1_ASAP7_75t_L g512 ( .A(n_195), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_195), .A2(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_196), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_206), .Y(n_196) );
AND2x2_ASAP7_75t_L g399 ( .A(n_197), .B(n_396), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_197), .B(n_381), .Y(n_431) );
BUFx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g330 ( .A(n_198), .B(n_254), .Y(n_330) );
AND2x2_ASAP7_75t_L g379 ( .A(n_198), .B(n_225), .Y(n_379) );
INVx1_ASAP7_75t_L g425 ( .A(n_198), .Y(n_425) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_199), .Y(n_238) );
AND2x2_ASAP7_75t_L g280 ( .A(n_199), .B(n_254), .Y(n_280) );
INVx1_ASAP7_75t_L g297 ( .A(n_199), .Y(n_297) );
AND2x2_ASAP7_75t_L g303 ( .A(n_199), .B(n_218), .Y(n_303) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_203), .Y(n_496) );
INVx2_ASAP7_75t_L g523 ( .A(n_203), .Y(n_523) );
INVx1_ASAP7_75t_L g510 ( .A(n_205), .Y(n_510) );
AND2x2_ASAP7_75t_L g371 ( .A(n_206), .B(n_279), .Y(n_371) );
INVx2_ASAP7_75t_L g436 ( .A(n_206), .Y(n_436) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_218), .Y(n_206) );
AND2x2_ASAP7_75t_L g253 ( .A(n_207), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g266 ( .A(n_207), .B(n_226), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_207), .B(n_225), .Y(n_294) );
INVx1_ASAP7_75t_L g300 ( .A(n_207), .Y(n_300) );
INVx1_ASAP7_75t_L g317 ( .A(n_207), .Y(n_317) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_207), .Y(n_329) );
INVx2_ASAP7_75t_L g397 ( .A(n_207), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
BUFx2_ASAP7_75t_L g351 ( .A(n_218), .Y(n_351) );
AND2x2_ASAP7_75t_L g396 ( .A(n_218), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_224), .B(n_333), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_224), .A2(n_395), .B(n_409), .Y(n_419) );
AND2x2_ASAP7_75t_L g444 ( .A(n_224), .B(n_330), .Y(n_444) );
BUFx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g366 ( .A(n_226), .Y(n_366) );
AND2x2_ASAP7_75t_L g395 ( .A(n_226), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_227), .Y(n_279) );
INVx2_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_227), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g252 ( .A(n_238), .Y(n_252) );
OR2x2_ASAP7_75t_L g265 ( .A(n_238), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g333 ( .A(n_238), .B(n_329), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_238), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g434 ( .A(n_238), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_238), .B(n_371), .Y(n_446) );
AND2x2_ASAP7_75t_L g325 ( .A(n_239), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g348 ( .A(n_239), .B(n_241), .Y(n_348) );
INVx2_ASAP7_75t_L g260 ( .A(n_240), .Y(n_260) );
AND2x2_ASAP7_75t_L g288 ( .A(n_240), .B(n_261), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_240), .B(n_313), .Y(n_369) );
AND2x2_ASAP7_75t_L g283 ( .A(n_241), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g430 ( .A(n_241), .Y(n_430) );
AND2x2_ASAP7_75t_L g442 ( .A(n_241), .B(n_305), .Y(n_442) );
AND2x2_ASAP7_75t_L g268 ( .A(n_242), .B(n_258), .Y(n_268) );
INVx1_ASAP7_75t_L g363 ( .A(n_242), .Y(n_363) );
AO21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_247), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_243), .B(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g515 ( .A(n_243), .Y(n_515) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_243), .A2(n_528), .B(n_535), .Y(n_527) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_243), .A2(n_584), .B(n_591), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_243), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g261 ( .A(n_248), .B(n_262), .Y(n_261) );
INVxp67_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_255), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_252), .B(n_299), .Y(n_308) );
OR2x2_ASAP7_75t_L g440 ( .A(n_252), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g357 ( .A(n_253), .B(n_298), .Y(n_357) );
AND2x2_ASAP7_75t_L g365 ( .A(n_253), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g424 ( .A(n_253), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g448 ( .A(n_253), .B(n_295), .Y(n_448) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_254), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g435 ( .A(n_254), .B(n_298), .Y(n_435) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2x1p5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
AND2x2_ASAP7_75t_L g287 ( .A(n_257), .B(n_288), .Y(n_287) );
INVxp67_ASAP7_75t_L g449 ( .A(n_257), .Y(n_449) );
NOR2x1_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g284 ( .A(n_260), .Y(n_284) );
AND2x2_ASAP7_75t_L g335 ( .A(n_260), .B(n_268), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_260), .B(n_403), .Y(n_429) );
INVx2_ASAP7_75t_L g274 ( .A(n_261), .Y(n_274) );
INVx3_ASAP7_75t_L g326 ( .A(n_261), .Y(n_326) );
OR2x2_ASAP7_75t_L g354 ( .A(n_261), .B(n_355), .Y(n_354) );
AOI311xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .A3(n_269), .B(n_270), .C(n_281), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_264), .A2(n_302), .B(n_304), .C(n_306), .Y(n_301) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_SL g286 ( .A(n_266), .Y(n_286) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g304 ( .A(n_268), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_268), .B(n_284), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_268), .B(n_269), .Y(n_437) );
AND2x2_ASAP7_75t_L g359 ( .A(n_269), .B(n_273), .Y(n_359) );
AOI21xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_275), .B(n_276), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g417 ( .A(n_273), .B(n_305), .Y(n_417) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_274), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g311 ( .A(n_274), .Y(n_311) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
AND2x2_ASAP7_75t_L g302 ( .A(n_278), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g347 ( .A(n_280), .Y(n_347) );
AND2x4_ASAP7_75t_L g409 ( .A(n_280), .B(n_378), .Y(n_409) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AOI222xp33_ASAP7_75t_L g360 ( .A1(n_283), .A2(n_349), .B1(n_361), .B2(n_365), .C1(n_367), .C2(n_371), .Y(n_360) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_289), .C(n_292), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_286), .B(n_330), .Y(n_353) );
INVx1_ASAP7_75t_L g375 ( .A(n_288), .Y(n_375) );
INVx1_ASAP7_75t_L g309 ( .A(n_290), .Y(n_309) );
OR2x2_ASAP7_75t_L g374 ( .A(n_291), .B(n_375), .Y(n_374) );
OAI21xp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_299), .Y(n_292) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_293), .B(n_311), .C(n_312), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_293), .A2(n_330), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_297), .Y(n_350) );
AND2x2_ASAP7_75t_SL g316 ( .A(n_298), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g407 ( .A(n_298), .Y(n_407) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_298), .Y(n_423) );
INVx2_ASAP7_75t_L g381 ( .A(n_299), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_303), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g355 ( .A(n_305), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B1(n_310), .B2(n_314), .C(n_315), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_309), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g443 ( .A(n_309), .Y(n_443) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g324 ( .A(n_316), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_316), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g382 ( .A(n_316), .B(n_330), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_316), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g415 ( .A(n_316), .B(n_350), .Y(n_415) );
BUFx3_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND5xp2_ASAP7_75t_L g320 ( .A(n_321), .B(n_339), .C(n_360), .D(n_372), .E(n_387), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI32xp33_ASAP7_75t_L g412 ( .A1(n_324), .A2(n_351), .A3(n_367), .B1(n_413), .B2(n_415), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_326), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g336 ( .A(n_330), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B1(n_336), .B2(n_337), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_346), .B1(n_348), .B2(n_349), .C(n_352), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g411 ( .A(n_343), .B(n_362), .Y(n_411) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_348), .A2(n_409), .B1(n_427), .B2(n_432), .C(n_433), .Y(n_426) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx2_ASAP7_75t_L g392 ( .A(n_351), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_356), .B2(n_358), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g370 ( .A(n_362), .Y(n_370) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_376), .B1(n_380), .B2(n_381), .C1(n_382), .C2(n_383), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_381), .A2(n_428), .B1(n_430), .B2(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B(n_393), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_398), .B(n_400), .Y(n_393) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g441 ( .A(n_396), .Y(n_441) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_408), .B(n_410), .C(n_412), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B(n_420), .C(n_445), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_417), .Y(n_421) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI211xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B(n_426), .C(n_438), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B(n_437), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_452), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_461), .Y(n_467) );
NOR2x2_ASAP7_75t_L g779 ( .A(n_462), .B(n_762), .Y(n_779) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g761 ( .A(n_463), .B(n_762), .Y(n_761) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_465), .B(n_469), .C(n_780), .Y(n_468) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_472), .B1(n_475), .B2(n_761), .Y(n_470) );
INVx1_ASAP7_75t_L g774 ( .A(n_471), .Y(n_774) );
OAI22x1_ASAP7_75t_SL g773 ( .A1(n_472), .A2(n_476), .B1(n_774), .B2(n_775), .Y(n_773) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR3x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_675), .C(n_718), .Y(n_476) );
NAND5xp2_ASAP7_75t_L g477 ( .A(n_478), .B(n_602), .C(n_632), .D(n_649), .E(n_664), .Y(n_477) );
AOI221xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_525), .B1(n_565), .B2(n_571), .C(n_575), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_501), .Y(n_479) );
OR2x2_ASAP7_75t_L g580 ( .A(n_480), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g619 ( .A(n_480), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g637 ( .A(n_480), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_480), .B(n_573), .Y(n_654) );
OR2x2_ASAP7_75t_L g666 ( .A(n_480), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_480), .B(n_625), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_480), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_480), .B(n_603), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_480), .B(n_611), .Y(n_717) );
AND2x2_ASAP7_75t_L g749 ( .A(n_480), .B(n_513), .Y(n_749) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_480), .Y(n_757) );
INVx5_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_481), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g577 ( .A(n_481), .B(n_555), .Y(n_577) );
BUFx2_ASAP7_75t_L g599 ( .A(n_481), .Y(n_599) );
AND2x2_ASAP7_75t_L g628 ( .A(n_481), .B(n_502), .Y(n_628) );
AND2x2_ASAP7_75t_L g683 ( .A(n_481), .B(n_581), .Y(n_683) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_499), .Y(n_481) );
BUFx2_ASAP7_75t_L g505 ( .A(n_484), .Y(n_505) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g517 ( .A1(n_488), .A2(n_498), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g559 ( .A1(n_488), .A2(n_498), .B(n_560), .C(n_561), .Y(n_559) );
INVx5_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_495), .C(n_496), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_493), .A2(n_496), .B(n_552), .C(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_501), .B(n_637), .Y(n_646) );
OAI32xp33_ASAP7_75t_L g660 ( .A1(n_501), .A2(n_596), .A3(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_501), .B(n_662), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_501), .B(n_580), .Y(n_703) );
INVx1_ASAP7_75t_SL g732 ( .A(n_501), .Y(n_732) );
NAND4xp25_ASAP7_75t_L g741 ( .A(n_501), .B(n_527), .C(n_683), .D(n_742), .Y(n_741) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_513), .Y(n_501) );
INVx5_ASAP7_75t_L g574 ( .A(n_502), .Y(n_574) );
AND2x2_ASAP7_75t_L g603 ( .A(n_502), .B(n_514), .Y(n_603) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_502), .Y(n_682) );
AND2x2_ASAP7_75t_L g752 ( .A(n_502), .B(n_699), .Y(n_752) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_511), .Y(n_502) );
AOI21xp5_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_506), .B(n_510), .Y(n_503) );
AND2x4_ASAP7_75t_L g625 ( .A(n_513), .B(n_574), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_513), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g659 ( .A(n_513), .B(n_581), .Y(n_659) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g573 ( .A(n_514), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g611 ( .A(n_514), .B(n_583), .Y(n_611) );
AND2x2_ASAP7_75t_L g620 ( .A(n_514), .B(n_582), .Y(n_620) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_524), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g688 ( .A1(n_525), .A2(n_689), .B1(n_691), .B2(n_693), .C1(n_696), .C2(n_697), .Y(n_688) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_544), .Y(n_525) );
AND2x2_ASAP7_75t_L g621 ( .A(n_526), .B(n_622), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_526), .B(n_599), .C(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
INVx5_ASAP7_75t_SL g570 ( .A(n_527), .Y(n_570) );
OAI322xp33_ASAP7_75t_L g575 ( .A1(n_527), .A2(n_576), .A3(n_578), .B1(n_579), .B2(n_593), .C1(n_596), .C2(n_598), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_527), .B(n_568), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_527), .B(n_556), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_531), .Y(n_528) );
INVx2_ASAP7_75t_L g568 ( .A(n_537), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_537), .B(n_546), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_544), .B(n_606), .Y(n_661) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g640 ( .A(n_545), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_555), .Y(n_545) );
OR2x2_ASAP7_75t_L g569 ( .A(n_546), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_546), .B(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g608 ( .A(n_546), .B(n_556), .Y(n_608) );
AND2x2_ASAP7_75t_L g631 ( .A(n_546), .B(n_568), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_546), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g647 ( .A(n_546), .B(n_606), .Y(n_647) );
AND2x2_ASAP7_75t_L g655 ( .A(n_546), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_546), .B(n_615), .Y(n_705) );
INVx5_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g595 ( .A(n_547), .B(n_570), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_547), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g622 ( .A(n_547), .B(n_556), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_547), .B(n_669), .Y(n_710) );
OR2x2_ASAP7_75t_L g726 ( .A(n_547), .B(n_670), .Y(n_726) );
AND2x2_ASAP7_75t_SL g733 ( .A(n_547), .B(n_687), .Y(n_733) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_547), .Y(n_740) );
OR2x6_ASAP7_75t_L g547 ( .A(n_548), .B(n_554), .Y(n_547) );
AND2x2_ASAP7_75t_L g594 ( .A(n_555), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g644 ( .A(n_555), .B(n_568), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_555), .B(n_570), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_555), .B(n_606), .Y(n_728) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_556), .B(n_570), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_556), .B(n_568), .Y(n_616) );
OR2x2_ASAP7_75t_L g670 ( .A(n_556), .B(n_568), .Y(n_670) );
AND2x2_ASAP7_75t_L g687 ( .A(n_556), .B(n_567), .Y(n_687) );
INVxp67_ASAP7_75t_L g709 ( .A(n_556), .Y(n_709) );
AND2x2_ASAP7_75t_L g736 ( .A(n_556), .B(n_606), .Y(n_736) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_556), .Y(n_743) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B(n_564), .Y(n_556) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_567), .B(n_617), .Y(n_690) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g606 ( .A(n_568), .B(n_570), .Y(n_606) );
OR2x2_ASAP7_75t_L g673 ( .A(n_568), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g617 ( .A(n_569), .Y(n_617) );
OR2x2_ASAP7_75t_L g678 ( .A(n_569), .B(n_670), .Y(n_678) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g578 ( .A(n_573), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_573), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g579 ( .A(n_574), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_574), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_574), .B(n_581), .Y(n_613) );
INVx2_ASAP7_75t_L g658 ( .A(n_574), .Y(n_658) );
AND2x2_ASAP7_75t_L g671 ( .A(n_574), .B(n_611), .Y(n_671) );
AND2x2_ASAP7_75t_L g696 ( .A(n_574), .B(n_620), .Y(n_696) );
INVx1_ASAP7_75t_L g648 ( .A(n_579), .Y(n_648) );
INVx2_ASAP7_75t_SL g635 ( .A(n_580), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_581), .Y(n_638) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_582), .Y(n_601) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
BUFx2_ASAP7_75t_L g699 ( .A(n_583), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g668 ( .A(n_595), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g674 ( .A(n_595), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_595), .A2(n_677), .B1(n_679), .B2(n_684), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_595), .B(n_687), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_596), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g630 ( .A(n_597), .Y(n_630) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
OR2x2_ASAP7_75t_L g612 ( .A(n_599), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_599), .B(n_603), .Y(n_663) );
AND2x2_ASAP7_75t_L g686 ( .A(n_599), .B(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g662 ( .A(n_601), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_609), .C(n_623), .Y(n_602) );
INVx1_ASAP7_75t_L g626 ( .A(n_603), .Y(n_626) );
OAI221xp5_ASAP7_75t_SL g734 ( .A1(n_603), .A2(n_735), .B1(n_737), .B2(n_738), .C(n_741), .Y(n_734) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g753 ( .A(n_606), .Y(n_753) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g702 ( .A(n_608), .B(n_641), .Y(n_702) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B(n_614), .C(n_618), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OAI32xp33_ASAP7_75t_L g727 ( .A1(n_616), .A2(n_617), .A3(n_680), .B1(n_717), .B2(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
AND2x2_ASAP7_75t_L g759 ( .A(n_619), .B(n_658), .Y(n_759) );
AND2x2_ASAP7_75t_L g706 ( .A(n_620), .B(n_658), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_620), .B(n_628), .Y(n_724) );
AOI31xp33_ASAP7_75t_SL g623 ( .A1(n_624), .A2(n_626), .A3(n_627), .B(n_629), .Y(n_623) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_625), .B(n_637), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_625), .B(n_635), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_625), .A2(n_655), .B1(n_745), .B2(n_748), .C(n_750), .Y(n_744) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g650 ( .A(n_630), .B(n_651), .Y(n_650) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_639), .B1(n_642), .B2(n_645), .C1(n_647), .C2(n_648), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g715 ( .A(n_634), .Y(n_715) );
INVx1_ASAP7_75t_L g737 ( .A(n_637), .Y(n_737) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_640), .A2(n_751), .B1(n_753), .B2(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g656 ( .A(n_641), .Y(n_656) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B1(n_655), .B2(n_657), .C(n_660), .Y(n_649) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g694 ( .A(n_652), .B(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g746 ( .A(n_652), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g721 ( .A(n_657), .Y(n_721) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g685 ( .A(n_658), .Y(n_685) );
INVx1_ASAP7_75t_L g667 ( .A(n_659), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_662), .B(n_749), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B1(n_671), .B2(n_672), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g758 ( .A(n_671), .Y(n_758) );
INVxp33_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_673), .B(n_717), .Y(n_716) );
OAI32xp33_ASAP7_75t_L g707 ( .A1(n_674), .A2(n_708), .A3(n_709), .B1(n_710), .B2(n_711), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_688), .C(n_700), .D(n_712), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_683), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g693 ( .A(n_694), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_697), .A2(n_713), .B1(n_730), .B2(n_733), .C(n_734), .Y(n_729) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g748 ( .A(n_699), .B(n_749), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B1(n_704), .B2(n_706), .C(n_707), .Y(n_700) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_709), .B(n_740), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g718 ( .A(n_719), .B(n_729), .C(n_744), .D(n_755), .Y(n_718) );
O2A1O1Ixp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_723), .B(n_725), .C(n_727), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g760 ( .A(n_747), .Y(n_760) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_759), .B(n_760), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g776 ( .A(n_761), .Y(n_776) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
CKINVDCx14_ASAP7_75t_R g771 ( .A(n_768), .Y(n_771) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
endmodule