module fake_netlist_6_940_n_1695 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1695);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1695;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_55),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_25),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_3),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_121),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_39),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_40),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_23),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_34),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_86),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_18),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_52),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_29),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_18),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_26),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_60),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_54),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_47),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_15),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_103),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_26),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_65),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_88),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_10),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_124),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_119),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_24),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_29),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_72),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_81),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_74),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_142),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_78),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_44),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_120),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_42),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_24),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_38),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_129),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_21),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_38),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_66),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_113),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_27),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_92),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_53),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_117),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_25),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_111),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_22),
.Y(n_210)
);

INVxp33_ASAP7_75t_SL g211 ( 
.A(n_36),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_57),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_56),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_67),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_62),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_73),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_118),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_47),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_48),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_48),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_80),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_99),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_58),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_90),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_45),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_17),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_136),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_131),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_35),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_35),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_114),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_8),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_97),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_32),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_63),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_16),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_115),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_83),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_46),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_12),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_112),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_0),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_27),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_37),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_31),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_68),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_50),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_122),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_140),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_23),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_108),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_42),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_98),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_102),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_19),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_39),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_84),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_100),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_107),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_137),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_9),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_17),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_30),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_40),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_4),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_70),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_64),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_44),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_11),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_87),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_85),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_4),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_59),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_75),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_34),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_93),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_6),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_51),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_12),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_134),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_49),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_77),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_32),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_43),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_89),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_45),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_1),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_2),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_138),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_36),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_188),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_151),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_151),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_147),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_166),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_194),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_166),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_210),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_148),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_289),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_149),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_198),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_226),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_230),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_230),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_231),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_231),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_152),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_242),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_242),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_243),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_243),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_246),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_246),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_153),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_159),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_262),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_149),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_154),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_161),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_167),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_171),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_154),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_176),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_163),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_162),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_177),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_150),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_188),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_162),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_168),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_262),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_269),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_269),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_273),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_281),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_281),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_181),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_192),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_192),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_264),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_207),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_207),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_209),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_184),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_248),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_182),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_183),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_168),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_303),
.B(n_305),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_321),
.B(n_280),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_320),
.A2(n_180),
.B(n_174),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_303),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_302),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_309),
.B(n_214),
.Y(n_381)
);

NOR3xp33_ASAP7_75t_L g382 ( 
.A(n_319),
.B(n_196),
.C(n_195),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_316),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_229),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_304),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_304),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_306),
.B(n_214),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_306),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_320),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_338),
.A2(n_202),
.B(n_173),
.Y(n_390)
);

CKINVDCx6p67_ASAP7_75t_R g391 ( 
.A(n_346),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_308),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_339),
.B(n_185),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_344),
.B(n_187),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_311),
.A2(n_203),
.B1(n_282),
.B2(n_294),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_328),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_155),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_371),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_335),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_315),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

NOR2x1_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_173),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_307),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_340),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_342),
.B(n_211),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_351),
.A2(n_352),
.B(n_310),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_361),
.B(n_202),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_343),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_366),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_361),
.B(n_224),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_362),
.B(n_224),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_324),
.Y(n_423)
);

OA21x2_ASAP7_75t_L g424 ( 
.A1(n_307),
.A2(n_180),
.B(n_174),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_310),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_312),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_312),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_364),
.B(n_189),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_364),
.B(n_251),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_324),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_348),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_313),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_313),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_325),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_426),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_426),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

AND3x2_ASAP7_75t_L g441 ( 
.A(n_382),
.B(n_317),
.C(n_259),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_386),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_345),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_426),
.Y(n_446)
);

AOI22x1_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_365),
.B1(n_251),
.B2(n_259),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_420),
.B(n_369),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_372),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_381),
.B(n_341),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_420),
.B(n_172),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_402),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_420),
.Y(n_453)
);

AND3x2_ASAP7_75t_L g454 ( 
.A(n_382),
.B(n_208),
.C(n_186),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_412),
.B(n_330),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_420),
.B(n_284),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_290),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_389),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_389),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_420),
.Y(n_461)
);

OAI22xp33_ASAP7_75t_L g462 ( 
.A1(n_398),
.A2(n_287),
.B1(n_199),
.B2(n_300),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_SL g463 ( 
.A(n_376),
.B(n_233),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_SL g465 ( 
.A(n_395),
.B(n_257),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_379),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_401),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_402),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_428),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_379),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_428),
.B(n_365),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_401),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_373),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_384),
.B(n_190),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_384),
.B(n_191),
.Y(n_476)
);

BUFx10_ASAP7_75t_L g477 ( 
.A(n_383),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_403),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_402),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_411),
.B(n_193),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_373),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_372),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_394),
.B(n_360),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_378),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_374),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_208),
.C(n_186),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_394),
.B(n_197),
.Y(n_490)
);

OR2x6_ASAP7_75t_L g491 ( 
.A(n_404),
.B(n_429),
.Y(n_491)
);

BUFx4f_ASAP7_75t_L g492 ( 
.A(n_424),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_418),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_378),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_374),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_379),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_377),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_377),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_378),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_378),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_378),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_379),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_380),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_416),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_397),
.B(n_200),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_380),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_385),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_429),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_397),
.B(n_201),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_415),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_385),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_375),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_375),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_432),
.Y(n_516)
);

OAI21xp33_ASAP7_75t_SL g517 ( 
.A1(n_390),
.A2(n_327),
.B(n_326),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_400),
.B(n_363),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_391),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_398),
.B(n_204),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_386),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_417),
.B(n_367),
.Y(n_522)
);

BUFx16f_ASAP7_75t_R g523 ( 
.A(n_391),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_375),
.B(n_415),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_386),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_375),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_416),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_396),
.A2(n_165),
.B1(n_164),
.B2(n_298),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_417),
.B(n_314),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_396),
.B(n_156),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_416),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_424),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_417),
.B(n_421),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_386),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_415),
.B(n_205),
.Y(n_536)
);

BUFx4f_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

CKINVDCx11_ASAP7_75t_R g538 ( 
.A(n_391),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_405),
.B(n_157),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_415),
.B(n_206),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_421),
.B(n_367),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_415),
.B(n_212),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_386),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_415),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_386),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_421),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_388),
.Y(n_547)
);

BUFx6f_ASAP7_75t_SL g548 ( 
.A(n_421),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_388),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_422),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_390),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_405),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_406),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_408),
.B(n_270),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_422),
.B(n_215),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_388),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_388),
.B(n_217),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_407),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_422),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_388),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_422),
.B(n_221),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_390),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_424),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_407),
.B(n_158),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_409),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_409),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_388),
.B(n_222),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_413),
.B(n_160),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_410),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_410),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_410),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_413),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_410),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_414),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_433),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_430),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_414),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_433),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_419),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_433),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_430),
.B(n_368),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_419),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_423),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_577),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_455),
.B(n_236),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_510),
.B(n_430),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_449),
.B(n_408),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_449),
.B(n_433),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_485),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_485),
.B(n_430),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_554),
.B(n_245),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_486),
.A2(n_258),
.B1(n_299),
.B2(n_295),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_530),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_450),
.B(n_169),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_533),
.B(n_387),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_546),
.A2(n_267),
.B1(n_253),
.B2(n_260),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_469),
.B(n_170),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_539),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_533),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_565),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_522),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_505),
.B(n_387),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_505),
.B(n_213),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_546),
.B(n_252),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_522),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_550),
.A2(n_263),
.B1(n_279),
.B2(n_283),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_458),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_477),
.B(n_293),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_550),
.B(n_286),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_560),
.B(n_288),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_506),
.B(n_527),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_490),
.B(n_175),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_507),
.B(n_178),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_506),
.B(n_213),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_529),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_458),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_527),
.A2(n_238),
.B1(n_275),
.B2(n_274),
.Y(n_618)
);

O2A1O1Ixp5_ASAP7_75t_L g619 ( 
.A1(n_492),
.A2(n_436),
.B(n_423),
.C(n_434),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_529),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_531),
.B(n_216),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_459),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_459),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_560),
.B(n_291),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_472),
.Y(n_625)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_462),
.A2(n_327),
.B1(n_326),
.B2(n_329),
.C(n_331),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_475),
.B(n_179),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_511),
.B(n_218),
.Y(n_628)
);

AO22x2_ASAP7_75t_L g629 ( 
.A1(n_520),
.A2(n_531),
.B1(n_535),
.B2(n_489),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_552),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_535),
.B(n_216),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_464),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_476),
.B(n_179),
.Y(n_633)
);

BUFx6f_ASAP7_75t_SL g634 ( 
.A(n_477),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_552),
.B(n_553),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_495),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_456),
.B(n_179),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_464),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_553),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_569),
.B(n_179),
.Y(n_640)
);

INVxp33_ASAP7_75t_L g641 ( 
.A(n_472),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_451),
.B(n_179),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_541),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_557),
.B(n_223),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_457),
.B(n_431),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_557),
.B(n_219),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_518),
.B(n_431),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_559),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_495),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_477),
.B(n_434),
.Y(n_650)
);

OR2x2_ASAP7_75t_SL g651 ( 
.A(n_463),
.B(n_223),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_516),
.B(n_436),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_491),
.A2(n_232),
.B1(n_225),
.B2(n_228),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_566),
.Y(n_654)
);

INVx8_ASAP7_75t_L g655 ( 
.A(n_491),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_489),
.A2(n_232),
.B1(n_254),
.B2(n_256),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_566),
.B(n_225),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_567),
.B(n_228),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_477),
.B(n_478),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_482),
.B(n_220),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_491),
.A2(n_548),
.B1(n_448),
.B2(n_555),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_567),
.B(n_235),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_541),
.B(n_368),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_573),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_573),
.B(n_235),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_SL g666 ( 
.A(n_548),
.B(n_227),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_467),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_491),
.A2(n_274),
.B1(n_240),
.B2(n_241),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_575),
.B(n_238),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_478),
.B(n_240),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_575),
.B(n_241),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_512),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_578),
.Y(n_673)
);

BUFx5_ASAP7_75t_L g674 ( 
.A(n_495),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_578),
.B(n_234),
.Y(n_675)
);

INVx8_ASAP7_75t_L g676 ( 
.A(n_491),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_580),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_582),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_478),
.B(n_250),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_478),
.B(n_250),
.Y(n_680)
);

AND2x4_ASAP7_75t_SL g681 ( 
.A(n_480),
.B(n_494),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_580),
.B(n_254),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_583),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_583),
.B(n_256),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_480),
.B(n_266),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_444),
.B(n_266),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_584),
.B(n_275),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_L g688 ( 
.A(n_532),
.B(n_292),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_584),
.B(n_237),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_582),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_487),
.B(n_292),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_467),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_528),
.B(n_331),
.C(n_329),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_487),
.B(n_500),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_480),
.B(n_239),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_562),
.B(n_244),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_514),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_465),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_514),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_515),
.Y(n_700)
);

BUFx6f_ASAP7_75t_SL g701 ( 
.A(n_480),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_551),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_538),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_500),
.B(n_425),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_501),
.B(n_425),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_515),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_526),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_474),
.B(n_332),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_470),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_519),
.B(n_392),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_526),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_474),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_551),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_470),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_548),
.B(n_247),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_501),
.B(n_425),
.Y(n_716)
);

AND2x6_ASAP7_75t_SL g717 ( 
.A(n_523),
.B(n_332),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_473),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_484),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_492),
.A2(n_393),
.B1(n_392),
.B2(n_427),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_502),
.B(n_427),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_532),
.B(n_249),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_502),
.B(n_427),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_473),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_564),
.B(n_435),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_492),
.A2(n_393),
.B1(n_435),
.B2(n_255),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_484),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_564),
.B(n_435),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_537),
.A2(n_359),
.B1(n_358),
.B2(n_357),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_488),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_519),
.B(n_95),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_551),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_570),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_570),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_494),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_494),
.B(n_272),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_537),
.A2(n_333),
.B(n_358),
.C(n_357),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_441),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_571),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_494),
.B(n_261),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_571),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_488),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_516),
.B(n_261),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_572),
.B(n_359),
.Y(n_744)
);

BUFx5_ASAP7_75t_L g745 ( 
.A(n_438),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_572),
.B(n_268),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_537),
.B(n_271),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_572),
.B(n_496),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_572),
.B(n_356),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_496),
.B(n_276),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_574),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_498),
.B(n_356),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_536),
.A2(n_277),
.B1(n_278),
.B2(n_285),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_600),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_595),
.A2(n_542),
.B1(n_540),
.B2(n_568),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_702),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_694),
.A2(n_563),
.B(n_461),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_674),
.B(n_574),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_674),
.B(n_576),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_594),
.B(n_499),
.Y(n_760)
);

OAI21xp33_ASAP7_75t_L g761 ( 
.A1(n_595),
.A2(n_517),
.B(n_354),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_733),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_589),
.A2(n_453),
.B(n_461),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_609),
.A2(n_499),
.B1(n_513),
.B2(n_509),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_625),
.B(n_454),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_748),
.A2(n_453),
.B(n_558),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_712),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_594),
.B(n_504),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_681),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_734),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_735),
.B(n_517),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_618),
.A2(n_656),
.B1(n_729),
.B2(n_629),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_599),
.A2(n_504),
.B1(n_513),
.B2(n_509),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_739),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_618),
.A2(n_656),
.B1(n_729),
.B2(n_629),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_741),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_719),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_727),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_599),
.B(n_508),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_601),
.B(n_576),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_751),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_730),
.Y(n_782)
);

AND3x2_ASAP7_75t_SL g783 ( 
.A(n_651),
.B(n_523),
.C(n_265),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_674),
.B(n_579),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_601),
.B(n_508),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_674),
.B(n_579),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_585),
.B(n_333),
.Y(n_787)
);

BUFx12f_ASAP7_75t_SL g788 ( 
.A(n_740),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_613),
.B(n_581),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_590),
.B(n_265),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_643),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_590),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_SL g793 ( 
.A(n_634),
.B(n_581),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_743),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_613),
.B(n_438),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_643),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_629),
.A2(n_447),
.B1(n_355),
.B2(n_354),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_702),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_614),
.B(n_452),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_652),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_603),
.A2(n_447),
.B1(n_337),
.B2(n_355),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_614),
.A2(n_544),
.B1(n_481),
.B2(n_468),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_742),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_636),
.B(n_503),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_636),
.A2(n_524),
.B1(n_452),
.B2(n_460),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_628),
.B(n_460),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_634),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_674),
.B(n_468),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_674),
.B(n_481),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_708),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_628),
.A2(n_334),
.B1(n_337),
.B2(n_353),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_697),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_708),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_702),
.B(n_483),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_SL g815 ( 
.A(n_626),
.B(n_334),
.C(n_353),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_713),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_602),
.B(n_503),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_691),
.A2(n_437),
.B1(n_445),
.B2(n_442),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_713),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_596),
.B(n_503),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_588),
.B(n_503),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_630),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_R g823 ( 
.A(n_703),
.B(n_466),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_604),
.A2(n_446),
.B1(n_445),
.B2(n_442),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_591),
.B(n_649),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_639),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_649),
.B(n_466),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_648),
.B(n_466),
.Y(n_828)
);

INVx5_ASAP7_75t_L g829 ( 
.A(n_713),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_701),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_698),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_699),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_L g833 ( 
.A(n_732),
.B(n_483),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_654),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_698),
.B(n_544),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_626),
.A2(n_314),
.B(n_437),
.C(n_439),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_701),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_664),
.B(n_497),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_732),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_615),
.A2(n_631),
.B1(n_621),
.B2(n_693),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_641),
.B(n_606),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_663),
.Y(n_842)
);

INVx5_ASAP7_75t_L g843 ( 
.A(n_732),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_746),
.B(n_439),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_726),
.A2(n_471),
.B1(n_493),
.B2(n_497),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_673),
.B(n_497),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_663),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_693),
.A2(n_440),
.B1(n_446),
.B2(n_549),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_SL g849 ( 
.A(n_598),
.B(n_0),
.C(n_1),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_677),
.B(n_471),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_616),
.Y(n_851)
);

XOR2xp5_ASAP7_75t_L g852 ( 
.A(n_661),
.B(n_94),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_620),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_655),
.Y(n_854)
);

AO22x1_ASAP7_75t_L g855 ( 
.A1(n_696),
.A2(n_440),
.B1(n_556),
.B2(n_549),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_612),
.B(n_561),
.Y(n_856)
);

NOR2x2_ASAP7_75t_L g857 ( 
.A(n_717),
.B(n_561),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_683),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_678),
.B(n_690),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_700),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_672),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_587),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_746),
.B(n_512),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_738),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_725),
.A2(n_443),
.B(n_534),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_647),
.B(n_471),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_644),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_598),
.Y(n_868)
);

BUFx8_ASAP7_75t_L g869 ( 
.A(n_706),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_710),
.B(n_493),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_731),
.B(n_493),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_635),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_659),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_704),
.Y(n_874)
);

NOR2x2_ASAP7_75t_L g875 ( 
.A(n_653),
.B(n_556),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_707),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_711),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_655),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_722),
.B(n_521),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_752),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_586),
.B(n_521),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_646),
.B(n_547),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_608),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_617),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_622),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_688),
.A2(n_545),
.B1(n_543),
.B2(n_547),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_722),
.B(n_521),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_646),
.B(n_545),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_672),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_744),
.B(n_749),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_657),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_675),
.B(n_543),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_650),
.B(n_534),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_623),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_632),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_593),
.Y(n_896)
);

CKINVDCx11_ASAP7_75t_R g897 ( 
.A(n_655),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_638),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_745),
.B(n_747),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_675),
.B(n_483),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_676),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_705),
.A2(n_512),
.B1(n_483),
.B2(n_534),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_689),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_676),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_667),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_692),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_689),
.B(n_483),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_676),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_709),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_658),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_670),
.B(n_679),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_750),
.B(n_512),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_662),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_680),
.B(n_534),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_750),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_666),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_728),
.B(n_512),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_665),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_669),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_685),
.B(n_443),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_714),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_645),
.B(n_443),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_716),
.A2(n_443),
.B1(n_479),
.B2(n_525),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_696),
.B(n_2),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_592),
.B(n_5),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_671),
.B(n_479),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_718),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_682),
.B(n_479),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_724),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_745),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_684),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_687),
.B(n_479),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_660),
.B(n_479),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_745),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_721),
.B(n_479),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_723),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_715),
.Y(n_937)
);

OR2x6_ASAP7_75t_L g938 ( 
.A(n_695),
.B(n_5),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_745),
.B(n_525),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_899),
.A2(n_637),
.B(n_737),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_896),
.A2(n_624),
.B1(n_605),
.B2(n_611),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_792),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_872),
.B(n_668),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_903),
.B(n_736),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_868),
.B(n_597),
.Y(n_945)
);

OAI21xp33_ASAP7_75t_L g946 ( 
.A1(n_800),
.A2(n_753),
.B(n_607),
.Y(n_946)
);

AOI221xp5_ASAP7_75t_L g947 ( 
.A1(n_903),
.A2(n_610),
.B1(n_640),
.B2(n_627),
.C(n_633),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_924),
.A2(n_619),
.B(n_720),
.C(n_686),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_794),
.B(n_619),
.Y(n_949)
);

AO22x2_ASAP7_75t_L g950 ( 
.A1(n_852),
.A2(n_642),
.B1(n_7),
.B2(n_9),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_822),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_899),
.A2(n_525),
.B(n_745),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_826),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_812),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_915),
.A2(n_525),
.B(n_7),
.C(n_10),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_872),
.B(n_6),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_925),
.A2(n_525),
.B(n_14),
.C(n_16),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_874),
.B(n_13),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_874),
.B(n_14),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_925),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_832),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_862),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_829),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_760),
.A2(n_20),
.B(n_22),
.C(n_28),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_788),
.B(n_82),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_930),
.A2(n_525),
.B(n_91),
.Y(n_966)
);

O2A1O1Ixp5_ASAP7_75t_L g967 ( 
.A1(n_863),
.A2(n_79),
.B(n_143),
.C(n_139),
.Y(n_967)
);

OA21x2_ASAP7_75t_L g968 ( 
.A1(n_879),
.A2(n_887),
.B(n_761),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_768),
.B(n_28),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_930),
.A2(n_61),
.B(n_106),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_834),
.Y(n_971)
);

OAI21xp33_ASAP7_75t_SL g972 ( 
.A1(n_772),
.A2(n_30),
.B(n_31),
.Y(n_972)
);

O2A1O1Ixp5_ASAP7_75t_SL g973 ( 
.A1(n_844),
.A2(n_33),
.B(n_41),
.C(n_43),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_862),
.B(n_33),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_816),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_876),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_SL g977 ( 
.A(n_873),
.B(n_937),
.C(n_830),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_863),
.A2(n_101),
.B(n_104),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_757),
.A2(n_105),
.B(n_144),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_779),
.A2(n_785),
.B(n_815),
.C(n_791),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_890),
.A2(n_41),
.B(n_46),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_912),
.A2(n_825),
.B(n_900),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_829),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_775),
.A2(n_811),
.B1(n_902),
.B2(n_840),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_R g985 ( 
.A(n_807),
.B(n_837),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_911),
.A2(n_847),
.B1(n_842),
.B2(n_771),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_907),
.A2(n_833),
.B(n_814),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_867),
.B(n_891),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_855),
.A2(n_844),
.B(n_892),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_775),
.A2(n_811),
.B1(n_902),
.B2(n_840),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_831),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_917),
.A2(n_820),
.B(n_766),
.Y(n_992)
);

NAND2x1p5_ASAP7_75t_L g993 ( 
.A(n_829),
.B(n_839),
.Y(n_993)
);

NOR2xp67_ASAP7_75t_L g994 ( 
.A(n_864),
.B(n_841),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_795),
.A2(n_806),
.B(n_799),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_933),
.A2(n_789),
.B(n_827),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_816),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_790),
.B(n_859),
.Y(n_998)
);

BUFx12f_ASAP7_75t_L g999 ( 
.A(n_897),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_SL g1000 ( 
.A(n_829),
.B(n_839),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_913),
.B(n_918),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_815),
.A2(n_797),
.B1(n_836),
.B2(n_931),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_841),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_797),
.A2(n_836),
.B1(n_858),
.B2(n_853),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_880),
.A2(n_919),
.B(n_910),
.C(n_881),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_823),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_754),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_816),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_839),
.B(n_843),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_851),
.A2(n_853),
.B1(n_936),
.B2(n_923),
.Y(n_1010)
);

AND2x6_ASAP7_75t_SL g1011 ( 
.A(n_938),
.B(n_765),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_810),
.A2(n_813),
.B1(n_916),
.B2(n_910),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_839),
.B(n_843),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_767),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_865),
.A2(n_821),
.B(n_786),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_851),
.B(n_780),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_823),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_791),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_758),
.A2(n_784),
.B(n_786),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_869),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_843),
.B(n_816),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_796),
.B(n_765),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_893),
.A2(n_920),
.B1(n_914),
.B2(n_835),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_877),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_843),
.B(n_861),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_936),
.A2(n_923),
.B1(n_801),
.B2(n_796),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_936),
.B(n_817),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_861),
.B(n_764),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_787),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_758),
.A2(n_784),
.B(n_759),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_882),
.B(n_888),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_787),
.B(n_878),
.Y(n_1032)
);

BUFx4f_ASAP7_75t_L g1033 ( 
.A(n_938),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_861),
.B(n_764),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_861),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_817),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_869),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_773),
.A2(n_938),
.B(n_849),
.C(n_803),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_SL g1039 ( 
.A(n_783),
.B(n_857),
.C(n_773),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_854),
.B(n_901),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_793),
.B(n_756),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_759),
.A2(n_939),
.B(n_808),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_756),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_936),
.B(n_778),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_849),
.A2(n_782),
.B(n_777),
.C(n_860),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_854),
.Y(n_1046)
);

CKINVDCx14_ASAP7_75t_R g1047 ( 
.A(n_769),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_883),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_808),
.A2(n_809),
.B(n_935),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_769),
.Y(n_1050)
);

AOI33xp33_ASAP7_75t_L g1051 ( 
.A1(n_801),
.A2(n_848),
.A3(n_885),
.B1(n_929),
.B2(n_884),
.B3(n_895),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_809),
.A2(n_763),
.B(n_922),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_875),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_894),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_934),
.A2(n_848),
.B1(n_909),
.B2(n_798),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_798),
.B(n_819),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_926),
.A2(n_932),
.B(n_928),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_755),
.A2(n_881),
.B(n_871),
.Y(n_1058)
);

AOI221x1_ASAP7_75t_L g1059 ( 
.A1(n_805),
.A2(n_845),
.B1(n_866),
.B2(n_846),
.C(n_850),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_866),
.A2(n_838),
.B(n_828),
.C(n_906),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_893),
.A2(n_920),
.B1(n_914),
.B2(n_870),
.Y(n_1061)
);

O2A1O1Ixp5_ASAP7_75t_L g1062 ( 
.A1(n_871),
.A2(n_870),
.B(n_819),
.C(n_927),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_889),
.A2(n_804),
.B(n_824),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_818),
.A2(n_824),
.B(n_802),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_889),
.A2(n_804),
.B(n_818),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_894),
.B(n_905),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_901),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_898),
.A2(n_921),
.B(n_770),
.C(n_774),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_SL g1069 ( 
.A(n_904),
.B(n_908),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_904),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_908),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_909),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_762),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_776),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_909),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_909),
.A2(n_886),
.B(n_781),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_886),
.B(n_783),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_856),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_856),
.A2(n_649),
.B(n_636),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_856),
.B(n_872),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_856),
.B(n_1015),
.Y(n_1081)
);

CKINVDCx11_ASAP7_75t_R g1082 ( 
.A(n_999),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1040),
.B(n_856),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1042),
.A2(n_1030),
.B(n_1019),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_995),
.A2(n_982),
.B(n_996),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_998),
.B(n_1029),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_1020),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1031),
.B(n_944),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1003),
.B(n_1053),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_991),
.B(n_994),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_984),
.B(n_990),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_953),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_R g1093 ( 
.A(n_977),
.B(n_1017),
.Y(n_1093)
);

AOI21xp33_ASAP7_75t_L g1094 ( 
.A1(n_984),
.A2(n_990),
.B(n_1002),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_992),
.A2(n_1058),
.B(n_987),
.Y(n_1095)
);

NOR4xp25_ASAP7_75t_L g1096 ( 
.A(n_960),
.B(n_964),
.C(n_957),
.D(n_1038),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1052),
.A2(n_952),
.B(n_1049),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_943),
.B(n_988),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_945),
.B(n_956),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_980),
.B(n_1027),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1057),
.A2(n_1034),
.B(n_1028),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1063),
.A2(n_1065),
.B(n_940),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1064),
.A2(n_968),
.B(n_948),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1046),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_971),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_941),
.B(n_1007),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1064),
.A2(n_968),
.B(n_1076),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1014),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_946),
.A2(n_979),
.B(n_1045),
.C(n_1005),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1060),
.A2(n_979),
.B(n_1055),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1002),
.A2(n_1061),
.B1(n_1023),
.B2(n_1026),
.Y(n_1111)
);

XNOR2xp5_ASAP7_75t_L g1112 ( 
.A(n_1006),
.B(n_1039),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1059),
.A2(n_989),
.B(n_1004),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_974),
.B(n_1018),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_969),
.B(n_958),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_991),
.B(n_1018),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1055),
.A2(n_1010),
.B(n_963),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1062),
.A2(n_1078),
.B(n_1010),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1051),
.B(n_1044),
.Y(n_1119)
);

AOI21x1_ASAP7_75t_SL g1120 ( 
.A1(n_959),
.A2(n_1080),
.B(n_1077),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_942),
.B(n_1022),
.Y(n_1121)
);

NOR2xp67_ASAP7_75t_L g1122 ( 
.A(n_1070),
.B(n_1035),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_966),
.A2(n_978),
.B(n_1004),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1036),
.B(n_962),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_973),
.A2(n_1026),
.B(n_967),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_986),
.A2(n_947),
.B(n_1012),
.C(n_972),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1001),
.B(n_1074),
.Y(n_1127)
);

BUFx8_ASAP7_75t_L g1128 ( 
.A(n_1037),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_955),
.A2(n_981),
.A3(n_1066),
.B(n_1016),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1046),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_949),
.B(n_976),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_1056),
.A2(n_970),
.A3(n_1048),
.B(n_961),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_954),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1075),
.A2(n_993),
.B(n_1070),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_950),
.B(n_1032),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_SL g1136 ( 
.A1(n_1041),
.A2(n_1021),
.B(n_1073),
.C(n_1008),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_963),
.A2(n_983),
.B(n_993),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_985),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1024),
.B(n_1054),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_SL g1140 ( 
.A(n_1046),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1075),
.A2(n_1025),
.B(n_1013),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1068),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_983),
.A2(n_1009),
.B(n_1069),
.Y(n_1143)
);

BUFx4_ASAP7_75t_SL g1144 ( 
.A(n_1011),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1072),
.A2(n_1035),
.B(n_975),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1067),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1033),
.B(n_1047),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_1071),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_1072),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_950),
.B(n_1071),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1072),
.A2(n_975),
.B(n_997),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_1071),
.B(n_1050),
.C(n_1043),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_965),
.B(n_975),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_997),
.A2(n_1079),
.B(n_1015),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_1043),
.A2(n_595),
.B1(n_462),
.B2(n_455),
.C(n_450),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_989),
.A2(n_855),
.B(n_863),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1079),
.A2(n_1015),
.B(n_1042),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1059),
.A2(n_984),
.A3(n_990),
.B(n_948),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1079),
.A2(n_1015),
.B(n_1042),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1031),
.B(n_872),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_951),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_SL g1162 ( 
.A1(n_941),
.A2(n_595),
.B(n_868),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1059),
.A2(n_996),
.B(n_982),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1059),
.A2(n_984),
.A3(n_990),
.B(n_948),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_984),
.A2(n_990),
.B(n_979),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1079),
.A2(n_1015),
.B(n_1042),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1079),
.A2(n_1015),
.B(n_1042),
.Y(n_1167)
);

O2A1O1Ixp5_ASAP7_75t_SL g1168 ( 
.A1(n_979),
.A2(n_640),
.B(n_1078),
.C(n_647),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1031),
.B(n_872),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_1005),
.A2(n_990),
.B(n_984),
.C(n_957),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1031),
.B(n_872),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1003),
.B(n_868),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_1046),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1059),
.A2(n_984),
.A3(n_990),
.B(n_948),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1077),
.A2(n_595),
.B1(n_924),
.B2(n_925),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_998),
.B(n_868),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1079),
.A2(n_1015),
.B(n_1042),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1031),
.B(n_872),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_995),
.A2(n_982),
.B(n_948),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1035),
.Y(n_1180)
);

BUFx2_ASAP7_75t_SL g1181 ( 
.A(n_1046),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_1046),
.Y(n_1182)
);

AO31x2_ASAP7_75t_L g1183 ( 
.A1(n_1059),
.A2(n_984),
.A3(n_990),
.B(n_948),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1059),
.A2(n_984),
.A3(n_990),
.B(n_948),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_998),
.B(n_868),
.Y(n_1185)
);

O2A1O1Ixp5_ASAP7_75t_L g1186 ( 
.A1(n_979),
.A2(n_595),
.B(n_990),
.C(n_984),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1046),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_998),
.B(n_868),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1046),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1079),
.A2(n_1015),
.B(n_1042),
.Y(n_1190)
);

O2A1O1Ixp5_ASAP7_75t_SL g1191 ( 
.A1(n_979),
.A2(n_640),
.B(n_1078),
.C(n_647),
.Y(n_1191)
);

INVxp67_ASAP7_75t_SL g1192 ( 
.A(n_1000),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_944),
.A2(n_903),
.B(n_924),
.C(n_595),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1079),
.A2(n_1015),
.B(n_1042),
.Y(n_1194)
);

AO21x2_ASAP7_75t_L g1195 ( 
.A1(n_996),
.A2(n_995),
.B(n_992),
.Y(n_1195)
);

AOI221xp5_ASAP7_75t_SL g1196 ( 
.A1(n_984),
.A2(n_990),
.B1(n_960),
.B2(n_1002),
.C(n_1038),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1003),
.B(n_868),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_942),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1059),
.A2(n_984),
.A3(n_990),
.B(n_948),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_1059),
.A2(n_996),
.B(n_982),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1031),
.B(n_872),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_999),
.B(n_904),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_951),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1059),
.A2(n_984),
.A3(n_990),
.B(n_948),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1079),
.A2(n_1015),
.B(n_1042),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_951),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1003),
.B(n_868),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1018),
.B(n_516),
.Y(n_1208)
);

INVx5_ASAP7_75t_L g1209 ( 
.A(n_963),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_995),
.A2(n_982),
.B(n_996),
.Y(n_1210)
);

AOI21x1_ASAP7_75t_L g1211 ( 
.A1(n_989),
.A2(n_855),
.B(n_863),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_951),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_995),
.A2(n_982),
.B(n_996),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_998),
.B(n_868),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_942),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_995),
.A2(n_982),
.B(n_948),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_SL g1217 ( 
.A1(n_1038),
.A2(n_1045),
.B(n_979),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_995),
.A2(n_982),
.B(n_948),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1083),
.B(n_1108),
.Y(n_1219)
);

INVx4_ASAP7_75t_L g1220 ( 
.A(n_1140),
.Y(n_1220)
);

AO21x2_ASAP7_75t_L g1221 ( 
.A1(n_1179),
.A2(n_1218),
.B(n_1216),
.Y(n_1221)
);

CKINVDCx6p67_ASAP7_75t_R g1222 ( 
.A(n_1140),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1203),
.Y(n_1223)
);

OAI211xp5_ASAP7_75t_SL g1224 ( 
.A1(n_1162),
.A2(n_1155),
.B(n_1175),
.C(n_1193),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1188),
.B(n_1214),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1148),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1111),
.Y(n_1227)
);

AO21x2_ASAP7_75t_L g1228 ( 
.A1(n_1179),
.A2(n_1218),
.B(n_1216),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1162),
.B(n_1088),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1092),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1099),
.B(n_1106),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1208),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1186),
.A2(n_1109),
.B(n_1126),
.C(n_1217),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1111),
.Y(n_1234)
);

NOR2x1_ASAP7_75t_SL g1235 ( 
.A(n_1209),
.B(n_1100),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1215),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1105),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1104),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1149),
.B(n_1133),
.Y(n_1240)
);

CKINVDCx8_ASAP7_75t_R g1241 ( 
.A(n_1181),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1104),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1118),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1098),
.B(n_1160),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1209),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1115),
.A2(n_1101),
.B(n_1096),
.Y(n_1246)
);

NAND3xp33_ASAP7_75t_L g1247 ( 
.A(n_1196),
.B(n_1096),
.C(n_1172),
.Y(n_1247)
);

OAI22x1_ASAP7_75t_L g1248 ( 
.A1(n_1150),
.A2(n_1135),
.B1(n_1112),
.B2(n_1185),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1091),
.A2(n_1094),
.B1(n_1113),
.B2(n_1171),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1091),
.A2(n_1094),
.B1(n_1113),
.B2(n_1171),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1089),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1161),
.B(n_1206),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1169),
.B(n_1178),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1196),
.B(n_1201),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1104),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1197),
.A2(n_1207),
.B1(n_1121),
.B2(n_1176),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_SL g1257 ( 
.A1(n_1103),
.A2(n_1114),
.B1(n_1086),
.B2(n_1125),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1117),
.A2(n_1125),
.B(n_1213),
.C(n_1085),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1159),
.A2(n_1177),
.B(n_1194),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1212),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1166),
.A2(n_1167),
.B(n_1190),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1139),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1210),
.A2(n_1095),
.B(n_1097),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1119),
.A2(n_1123),
.B(n_1131),
.C(n_1170),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1131),
.Y(n_1265)
);

BUFx8_ASAP7_75t_L g1266 ( 
.A(n_1087),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1130),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1119),
.A2(n_1084),
.B(n_1143),
.C(n_1142),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1205),
.A2(n_1156),
.B(n_1211),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1168),
.A2(n_1191),
.A3(n_1120),
.B(n_1200),
.Y(n_1270)
);

AOI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1163),
.A2(n_1200),
.B(n_1137),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1129),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1136),
.A2(n_1134),
.B(n_1141),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1124),
.B(n_1198),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1153),
.B(n_1116),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1151),
.A2(n_1145),
.B(n_1180),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1132),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1195),
.A2(n_1122),
.B(n_1192),
.Y(n_1278)
);

OR2x2_ASAP7_75t_L g1279 ( 
.A(n_1127),
.B(n_1146),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1180),
.A2(n_1152),
.B(n_1090),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1130),
.Y(n_1281)
);

OAI222xp33_ASAP7_75t_L g1282 ( 
.A1(n_1202),
.A2(n_1147),
.B1(n_1138),
.B2(n_1164),
.C1(n_1158),
.C2(n_1174),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1202),
.A2(n_1093),
.B1(n_1152),
.B2(n_1189),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1130),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1132),
.A2(n_1183),
.B(n_1204),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1209),
.A2(n_1184),
.B(n_1204),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1158),
.A2(n_1183),
.B(n_1204),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1132),
.A2(n_1174),
.B(n_1184),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_1173),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1129),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1129),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1158),
.A2(n_1183),
.B(n_1184),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1164),
.A2(n_1174),
.A3(n_1199),
.B(n_1144),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1173),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1173),
.Y(n_1295)
);

INVx4_ASAP7_75t_SL g1296 ( 
.A(n_1182),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1164),
.A2(n_1199),
.B(n_1182),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1187),
.A2(n_1189),
.B(n_1128),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1187),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1189),
.B(n_1128),
.Y(n_1300)
);

OAI222xp33_ASAP7_75t_L g1301 ( 
.A1(n_1082),
.A2(n_1091),
.B1(n_1175),
.B2(n_938),
.C1(n_1111),
.C2(n_852),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1111),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1088),
.B(n_1171),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1215),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1154),
.A2(n_1081),
.B(n_1095),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1188),
.B(n_1214),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1186),
.A2(n_990),
.B(n_984),
.C(n_1094),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1108),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1175),
.A2(n_1162),
.B1(n_868),
.B2(n_896),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1188),
.B(n_1214),
.Y(n_1310)
);

NOR2x1_ASAP7_75t_SL g1311 ( 
.A(n_1209),
.B(n_984),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1088),
.B(n_1171),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1154),
.A2(n_1081),
.B(n_1095),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1186),
.A2(n_990),
.B(n_984),
.C(n_1094),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1188),
.B(n_1214),
.Y(n_1315)
);

AOI22x1_ASAP7_75t_L g1316 ( 
.A1(n_1217),
.A2(n_924),
.B1(n_594),
.B2(n_601),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1154),
.A2(n_1081),
.B(n_1095),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1081),
.A2(n_1154),
.B(n_1157),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1165),
.A2(n_1110),
.A3(n_1102),
.B(n_1107),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1081),
.A2(n_1154),
.B(n_1157),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1186),
.A2(n_990),
.B(n_984),
.C(n_1094),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1148),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1140),
.Y(n_1323)
);

AO21x2_ASAP7_75t_L g1324 ( 
.A1(n_1179),
.A2(n_1218),
.B(n_1216),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1110),
.A2(n_1113),
.B(n_1216),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1165),
.A2(n_1094),
.B1(n_1175),
.B2(n_950),
.Y(n_1326)
);

AOI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1156),
.A2(n_1211),
.B(n_989),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1104),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1154),
.A2(n_1081),
.B(n_1095),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1188),
.B(n_1214),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1186),
.A2(n_990),
.B(n_984),
.C(n_1094),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1188),
.B(n_1214),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1108),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1154),
.A2(n_1081),
.B(n_1095),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1108),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1162),
.B(n_903),
.Y(n_1336)
);

AOI21xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1112),
.A2(n_519),
.B(n_595),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1188),
.B(n_1214),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1217),
.A2(n_1038),
.B(n_1045),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1188),
.B(n_1214),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1081),
.A2(n_1154),
.B(n_1157),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1156),
.A2(n_1211),
.B(n_989),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1110),
.A2(n_1113),
.B(n_1216),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1108),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1081),
.A2(n_1154),
.B(n_1157),
.Y(n_1345)
);

O2A1O1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1162),
.A2(n_1193),
.B(n_595),
.C(n_1186),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1110),
.A2(n_1113),
.B(n_1216),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1179),
.A2(n_1218),
.B(n_1216),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1081),
.A2(n_1154),
.B(n_1157),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1231),
.B(n_1303),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_SL g1351 ( 
.A1(n_1346),
.A2(n_1246),
.B(n_1224),
.C(n_1336),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1233),
.A2(n_1235),
.B(n_1307),
.Y(n_1352)
);

BUFx8_ASAP7_75t_SL g1353 ( 
.A(n_1300),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1326),
.A2(n_1247),
.B1(n_1229),
.B2(n_1309),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_SL g1355 ( 
.A(n_1241),
.B(n_1220),
.Y(n_1355)
);

INVx3_ASAP7_75t_SL g1356 ( 
.A(n_1222),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1301),
.A2(n_1314),
.B(n_1331),
.C(n_1307),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1225),
.B(n_1306),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1326),
.A2(n_1229),
.B1(n_1336),
.B2(n_1256),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1314),
.A2(n_1321),
.B(n_1331),
.C(n_1339),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1258),
.A2(n_1269),
.B(n_1285),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1297),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1272),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1231),
.B(n_1312),
.Y(n_1364)
);

O2A1O1Ixp5_ASAP7_75t_L g1365 ( 
.A1(n_1254),
.A2(n_1264),
.B(n_1268),
.C(n_1282),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1232),
.B(n_1279),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1266),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1244),
.B(n_1253),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1221),
.A2(n_1324),
.B(n_1348),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1310),
.B(n_1315),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1330),
.B(n_1332),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1338),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1277),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1340),
.B(n_1265),
.Y(n_1374)
);

NAND2xp33_ASAP7_75t_SL g1375 ( 
.A(n_1220),
.B(n_1323),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1298),
.Y(n_1376)
);

AND2x2_ASAP7_75t_SL g1377 ( 
.A(n_1325),
.B(n_1343),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1266),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1243),
.A2(n_1275),
.B(n_1240),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1265),
.B(n_1262),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1240),
.A2(n_1274),
.B(n_1252),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_SL g1382 ( 
.A1(n_1240),
.A2(n_1252),
.B(n_1239),
.Y(n_1382)
);

OA22x2_ASAP7_75t_L g1383 ( 
.A1(n_1248),
.A2(n_1251),
.B1(n_1219),
.B2(n_1252),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1293),
.B(n_1227),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1230),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1266),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1242),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1245),
.A2(n_1323),
.B(n_1311),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1249),
.A2(n_1250),
.B(n_1257),
.C(n_1227),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_SL g1390 ( 
.A1(n_1234),
.A2(n_1302),
.B(n_1316),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1337),
.A2(n_1283),
.B(n_1264),
.C(n_1268),
.Y(n_1391)
);

AOI221x1_ASAP7_75t_SL g1392 ( 
.A1(n_1283),
.A2(n_1237),
.B1(n_1260),
.B2(n_1344),
.C(n_1333),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1304),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1236),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1249),
.A2(n_1250),
.B1(n_1257),
.B2(n_1322),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1335),
.B(n_1223),
.Y(n_1396)
);

AOI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1234),
.A2(n_1302),
.B1(n_1290),
.B2(n_1228),
.C(n_1348),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1308),
.B(n_1293),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1245),
.A2(n_1325),
.B(n_1347),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1242),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1293),
.B(n_1295),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1238),
.B(n_1294),
.Y(n_1402)
);

AOI221xp5_ASAP7_75t_L g1403 ( 
.A1(n_1286),
.A2(n_1291),
.B1(n_1278),
.B2(n_1226),
.C(n_1267),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1285),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1238),
.B(n_1294),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1325),
.A2(n_1347),
.B(n_1343),
.C(n_1328),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1328),
.A2(n_1284),
.B1(n_1289),
.B2(n_1255),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1288),
.A2(n_1292),
.B(n_1280),
.C(n_1319),
.Y(n_1408)
);

NOR2xp67_ASAP7_75t_L g1409 ( 
.A(n_1255),
.B(n_1299),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1280),
.B(n_1276),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1255),
.B(n_1299),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1255),
.B(n_1299),
.Y(n_1412)
);

AOI21x1_ASAP7_75t_SL g1413 ( 
.A1(n_1270),
.A2(n_1296),
.B(n_1273),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1281),
.B(n_1296),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1281),
.B(n_1287),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1327),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1342),
.B(n_1271),
.Y(n_1417)
);

INVxp33_ASAP7_75t_L g1418 ( 
.A(n_1263),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1270),
.A2(n_1334),
.B(n_1329),
.C(n_1317),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1305),
.A2(n_1313),
.B(n_1320),
.C(n_1341),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1318),
.B(n_1320),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1259),
.B(n_1261),
.Y(n_1422)
);

BUFx8_ASAP7_75t_L g1423 ( 
.A(n_1345),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1349),
.B(n_1225),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1231),
.B(n_1303),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1326),
.A2(n_1175),
.B1(n_1247),
.B2(n_1162),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1231),
.B(n_1303),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1242),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1258),
.A2(n_1110),
.B(n_1113),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1225),
.B(n_1306),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1225),
.B(n_1306),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1301),
.A2(n_1162),
.B(n_1193),
.C(n_1346),
.Y(n_1432)
);

OR2x2_ASAP7_75t_SL g1433 ( 
.A(n_1247),
.B(n_1279),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1304),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1373),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1408),
.A2(n_1365),
.B(n_1369),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1377),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1410),
.B(n_1421),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1404),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1359),
.B(n_1354),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1380),
.B(n_1350),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1410),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1393),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1424),
.B(n_1422),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1429),
.B(n_1415),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1423),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1417),
.A2(n_1389),
.B(n_1399),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1429),
.B(n_1398),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1423),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1384),
.B(n_1363),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1361),
.B(n_1406),
.Y(n_1451)
);

NOR2x1_ASAP7_75t_L g1452 ( 
.A(n_1352),
.B(n_1389),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1364),
.B(n_1425),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1427),
.B(n_1368),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1397),
.A2(n_1362),
.B(n_1403),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1401),
.B(n_1418),
.Y(n_1456)
);

AOI322xp5_ASAP7_75t_L g1457 ( 
.A1(n_1358),
.A2(n_1431),
.A3(n_1430),
.B1(n_1370),
.B2(n_1371),
.C1(n_1372),
.C2(n_1357),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1385),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1418),
.B(n_1383),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1419),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1420),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1396),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1351),
.A2(n_1426),
.B(n_1360),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1351),
.B(n_1374),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1432),
.A2(n_1391),
.B(n_1413),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1416),
.Y(n_1466)
);

OAI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1395),
.A2(n_1394),
.B(n_1366),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1433),
.B(n_1376),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1392),
.B(n_1416),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1402),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1405),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1435),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1456),
.B(n_1434),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1445),
.B(n_1412),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1445),
.B(n_1411),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1442),
.B(n_1387),
.Y(n_1476)
);

AOI222xp33_ASAP7_75t_L g1477 ( 
.A1(n_1440),
.A2(n_1386),
.B1(n_1378),
.B2(n_1367),
.C1(n_1356),
.C2(n_1355),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1437),
.B(n_1400),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1452),
.A2(n_1386),
.B1(n_1367),
.B2(n_1378),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1438),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1458),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1445),
.B(n_1414),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1443),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1440),
.A2(n_1375),
.B1(n_1388),
.B2(n_1407),
.C(n_1356),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1456),
.B(n_1387),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1452),
.A2(n_1375),
.B1(n_1353),
.B2(n_1428),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1448),
.B(n_1409),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1439),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1448),
.B(n_1379),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1450),
.B(n_1390),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1448),
.B(n_1381),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1456),
.B(n_1353),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1448),
.B(n_1382),
.Y(n_1493)
);

AOI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1479),
.A2(n_1467),
.B1(n_1463),
.B2(n_1464),
.C(n_1469),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1488),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1488),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1482),
.B(n_1444),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1481),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1481),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1487),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1473),
.B(n_1437),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1472),
.Y(n_1502)
);

OAI211xp5_ASAP7_75t_L g1503 ( 
.A1(n_1477),
.A2(n_1467),
.B(n_1457),
.C(n_1464),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1483),
.Y(n_1504)
);

OAI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1484),
.A2(n_1469),
.B1(n_1466),
.B2(n_1457),
.C(n_1468),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1476),
.Y(n_1506)
);

OAI221xp5_ASAP7_75t_L g1507 ( 
.A1(n_1484),
.A2(n_1466),
.B1(n_1457),
.B2(n_1468),
.C(n_1454),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_R g1508 ( 
.A(n_1492),
.B(n_1466),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1477),
.A2(n_1463),
.B1(n_1465),
.B2(n_1447),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1485),
.B(n_1471),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1486),
.A2(n_1468),
.B(n_1449),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_R g1512 ( 
.A(n_1492),
.B(n_1443),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1478),
.B(n_1471),
.Y(n_1513)
);

OAI211xp5_ASAP7_75t_L g1514 ( 
.A1(n_1490),
.A2(n_1436),
.B(n_1441),
.C(n_1455),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1480),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1480),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1474),
.B(n_1470),
.Y(n_1517)
);

OAI31xp33_ASAP7_75t_L g1518 ( 
.A1(n_1491),
.A2(n_1463),
.A3(n_1453),
.B(n_1454),
.Y(n_1518)
);

AOI33xp33_ASAP7_75t_L g1519 ( 
.A1(n_1489),
.A2(n_1460),
.A3(n_1459),
.B1(n_1462),
.B2(n_1461),
.B3(n_1451),
.Y(n_1519)
);

NOR3xp33_ASAP7_75t_L g1520 ( 
.A(n_1503),
.B(n_1453),
.C(n_1460),
.Y(n_1520)
);

INVx4_ASAP7_75t_SL g1521 ( 
.A(n_1504),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1502),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1495),
.Y(n_1523)
);

INVx4_ASAP7_75t_SL g1524 ( 
.A(n_1504),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_L g1525 ( 
.A(n_1514),
.B(n_1463),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1495),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1496),
.B(n_1490),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1494),
.A2(n_1455),
.B(n_1490),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1500),
.B(n_1480),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1497),
.B(n_1493),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1504),
.Y(n_1531)
);

NOR3xp33_ASAP7_75t_SL g1532 ( 
.A(n_1508),
.B(n_1505),
.C(n_1511),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1498),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1516),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1518),
.B(n_1474),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1498),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1499),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1497),
.B(n_1487),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1506),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1506),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1522),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1521),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1520),
.B(n_1519),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1527),
.B(n_1501),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1520),
.B(n_1510),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1531),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1530),
.B(n_1538),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1539),
.B(n_1506),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1540),
.B(n_1521),
.Y(n_1550)
);

NOR2xp67_ASAP7_75t_L g1551 ( 
.A(n_1535),
.B(n_1516),
.Y(n_1551)
);

OR2x6_ASAP7_75t_L g1552 ( 
.A(n_1528),
.B(n_1511),
.Y(n_1552)
);

NAND4xp25_ASAP7_75t_L g1553 ( 
.A(n_1528),
.B(n_1509),
.C(n_1441),
.D(n_1461),
.Y(n_1553)
);

NOR3xp33_ASAP7_75t_SL g1554 ( 
.A(n_1535),
.B(n_1513),
.C(n_1461),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1537),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1521),
.B(n_1515),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1532),
.B(n_1517),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1522),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1537),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1533),
.Y(n_1560)
);

NAND2xp33_ASAP7_75t_L g1561 ( 
.A(n_1532),
.B(n_1512),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1525),
.A2(n_1465),
.B(n_1447),
.Y(n_1562)
);

INVxp67_ASAP7_75t_SL g1563 ( 
.A(n_1525),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1521),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1524),
.B(n_1475),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1524),
.B(n_1475),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1533),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1546),
.Y(n_1568)
);

NAND2x1_ASAP7_75t_SL g1569 ( 
.A(n_1542),
.B(n_1534),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1560),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1560),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1546),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1565),
.B(n_1524),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1567),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1546),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1567),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1566),
.B(n_1524),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1555),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1555),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1543),
.B(n_1523),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1548),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1541),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1559),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1561),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1566),
.B(n_1524),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1541),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1559),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1545),
.B(n_1526),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1541),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1550),
.B(n_1529),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1550),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1542),
.B(n_1547),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_SL g1594 ( 
.A(n_1542),
.B(n_1446),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1558),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1542),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1557),
.B(n_1536),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1558),
.Y(n_1598)
);

CKINVDCx16_ASAP7_75t_R g1599 ( 
.A(n_1594),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1570),
.B(n_1564),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1571),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1571),
.Y(n_1602)
);

INVx4_ASAP7_75t_L g1603 ( 
.A(n_1596),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1568),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1564),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1574),
.B(n_1547),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1597),
.B(n_1544),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1568),
.Y(n_1608)
);

CKINVDCx16_ASAP7_75t_R g1609 ( 
.A(n_1594),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1568),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1574),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1578),
.B(n_1549),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1582),
.A2(n_1552),
.B1(n_1553),
.B2(n_1562),
.Y(n_1613)
);

INVx4_ASAP7_75t_L g1614 ( 
.A(n_1596),
.Y(n_1614)
);

CKINVDCx16_ASAP7_75t_R g1615 ( 
.A(n_1578),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_SL g1616 ( 
.A1(n_1585),
.A2(n_1553),
.B(n_1563),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1573),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1573),
.B(n_1554),
.Y(n_1618)
);

OR2x6_ASAP7_75t_L g1619 ( 
.A(n_1573),
.B(n_1552),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1551),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_SL g1621 ( 
.A(n_1576),
.B(n_1552),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1586),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1586),
.B(n_1549),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1604),
.Y(n_1624)
);

AOI32xp33_ASAP7_75t_L g1625 ( 
.A1(n_1621),
.A2(n_1593),
.A3(n_1581),
.B1(n_1592),
.B2(n_1597),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1604),
.Y(n_1626)
);

NOR3xp33_ASAP7_75t_SL g1627 ( 
.A(n_1615),
.B(n_1581),
.C(n_1580),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1621),
.A2(n_1552),
.B1(n_1593),
.B2(n_1592),
.Y(n_1628)
);

O2A1O1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1616),
.A2(n_1552),
.B(n_1589),
.C(n_1576),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1615),
.B(n_1611),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1604),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1608),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1612),
.B(n_1591),
.Y(n_1633)
);

AOI222xp33_ASAP7_75t_L g1634 ( 
.A1(n_1616),
.A2(n_1551),
.B1(n_1589),
.B2(n_1588),
.C1(n_1584),
.C2(n_1580),
.Y(n_1634)
);

AOI322xp5_ASAP7_75t_L g1635 ( 
.A1(n_1613),
.A2(n_1591),
.A3(n_1579),
.B1(n_1588),
.B2(n_1584),
.C1(n_1577),
.C2(n_1572),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1612),
.B(n_1596),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1608),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1608),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1622),
.B(n_1596),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1610),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1603),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1623),
.B(n_1556),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1631),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1636),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1625),
.B(n_1599),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1633),
.B(n_1623),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1630),
.B(n_1599),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1631),
.Y(n_1648)
);

AOI221x1_ASAP7_75t_SL g1649 ( 
.A1(n_1639),
.A2(n_1618),
.B1(n_1600),
.B2(n_1620),
.C(n_1579),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1642),
.B(n_1605),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1624),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1626),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1636),
.B(n_1605),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1650),
.B(n_1627),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1645),
.A2(n_1629),
.B(n_1634),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1647),
.A2(n_1627),
.B(n_1619),
.C(n_1641),
.Y(n_1656)
);

AOI211xp5_ASAP7_75t_L g1657 ( 
.A1(n_1653),
.A2(n_1628),
.B(n_1600),
.C(n_1641),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1644),
.A2(n_1635),
.B(n_1619),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1643),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1643),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_SL g1661 ( 
.A(n_1650),
.B(n_1646),
.C(n_1648),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1642),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1648),
.A2(n_1609),
.B1(n_1600),
.B2(n_1619),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1651),
.Y(n_1664)
);

AOI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1655),
.A2(n_1652),
.B(n_1649),
.C(n_1637),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1663),
.A2(n_1600),
.B(n_1606),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1658),
.A2(n_1619),
.B1(n_1569),
.B2(n_1607),
.C(n_1610),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1656),
.A2(n_1609),
.B1(n_1638),
.B2(n_1640),
.C(n_1632),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1662),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1669),
.B(n_1657),
.Y(n_1670)
);

NOR2xp67_ASAP7_75t_L g1671 ( 
.A(n_1666),
.B(n_1661),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1665),
.Y(n_1672)
);

OAI31xp33_ASAP7_75t_L g1673 ( 
.A1(n_1667),
.A2(n_1654),
.A3(n_1660),
.B(n_1659),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1668),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1669),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1671),
.B(n_1664),
.Y(n_1676)
);

OAI21xp33_ASAP7_75t_L g1677 ( 
.A1(n_1674),
.A2(n_1619),
.B(n_1617),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1672),
.A2(n_1610),
.B1(n_1617),
.B2(n_1569),
.C(n_1603),
.Y(n_1678)
);

AOI21xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1670),
.A2(n_1617),
.B(n_1607),
.Y(n_1679)
);

NAND4xp75_ASAP7_75t_L g1680 ( 
.A(n_1673),
.B(n_1601),
.C(n_1602),
.D(n_1606),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1679),
.B(n_1670),
.Y(n_1681)
);

OAI32xp33_ASAP7_75t_L g1682 ( 
.A1(n_1676),
.A2(n_1675),
.A3(n_1614),
.B1(n_1603),
.B2(n_1601),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1677),
.A2(n_1614),
.B(n_1603),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1681),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1682),
.B1(n_1678),
.B2(n_1683),
.C(n_1614),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1685),
.B(n_1684),
.Y(n_1686)
);

OA22x2_ASAP7_75t_L g1687 ( 
.A1(n_1686),
.A2(n_1614),
.B1(n_1680),
.B2(n_1602),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1687),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1684),
.B(n_1587),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1689),
.B(n_1583),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1690),
.A2(n_1587),
.B(n_1583),
.Y(n_1691)
);

XNOR2xp5_ASAP7_75t_L g1692 ( 
.A(n_1691),
.B(n_1572),
.Y(n_1692)
);

AOI22x1_ASAP7_75t_L g1693 ( 
.A1(n_1691),
.A2(n_1583),
.B1(n_1587),
.B2(n_1598),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1692),
.A2(n_1575),
.B1(n_1577),
.B2(n_1590),
.C(n_1595),
.Y(n_1694)
);

AOI211xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1693),
.B(n_1590),
.C(n_1595),
.Y(n_1695)
);


endmodule