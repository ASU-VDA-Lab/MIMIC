module fake_jpeg_8124_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_0),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_13),
.B(n_15),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_11),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_20),
.B(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_19),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AO221x1_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_8),
.B1(n_7),
.B2(n_13),
.C(n_20),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_16),
.C(n_12),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.C(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AOI322xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.A3(n_33),
.B1(n_25),
.B2(n_29),
.C1(n_5),
.C2(n_3),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_21),
.C(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_32),
.Y(n_36)
);


endmodule