module real_jpeg_14733_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_2),
.A2(n_36),
.B1(n_40),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_2),
.Y(n_83)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_3),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_44),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_3),
.B(n_89),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_5),
.A2(n_29),
.B1(n_33),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_5),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_5),
.A2(n_36),
.B1(n_40),
.B2(n_65),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_29),
.B1(n_33),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_8),
.A2(n_36),
.B1(n_40),
.B2(n_72),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_10),
.A2(n_36),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_11),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_60)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_13),
.A2(n_36),
.B1(n_40),
.B2(n_57),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_92),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_86),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_18),
.B(n_86),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_61),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_47),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_21),
.B(n_34),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_24),
.B(n_27),
.C(n_32),
.Y(n_21)
);

OA22x2_ASAP7_75t_SL g68 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_22),
.A2(n_23),
.B1(n_29),
.B2(n_33),
.Y(n_69)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_25),
.C(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_25),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_24),
.B(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_28),
.A2(n_64),
.B1(n_67),
.B2(n_89),
.Y(n_88)
);

HAxp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_31),
.CON(n_28),
.SN(n_28)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_29),
.A2(n_33),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_31),
.B(n_40),
.C(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_31),
.B(n_44),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_31),
.B(n_54),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_41),
.B(n_43),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_35),
.B(n_42),
.Y(n_126)
);

CKINVDCx6p67_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_40),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_41),
.B(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_41),
.A2(n_42),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_82),
.B(n_84),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_44),
.A2(n_107),
.B1(n_115),
.B2(n_116),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_55),
.B(n_58),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_56),
.B1(n_59),
.B2(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_59),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_49),
.A2(n_59),
.B1(n_91),
.B2(n_102),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_73),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_81),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.C(n_90),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_90),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_133),
.B(n_137),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_122),
.B(n_132),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_110),
.B(n_121),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_105),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_103),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_116),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_117),
.B(n_120),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_119),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_124),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_128),
.C(n_131),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_136),
.Y(n_137)
);


endmodule