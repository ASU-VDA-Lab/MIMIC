module fake_jpeg_21271_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_SL g65 ( 
.A(n_6),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_89),
.Y(n_98)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_46),
.B1(n_61),
.B2(n_50),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_48),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_46),
.B1(n_49),
.B2(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_54),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_68),
.B1(n_59),
.B2(n_49),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_60),
.B1(n_72),
.B2(n_69),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_62),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_102),
.C(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_54),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_71),
.A3(n_63),
.B1(n_54),
.B2(n_60),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_106),
.B1(n_107),
.B2(n_69),
.Y(n_126)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_57),
.B1(n_71),
.B2(n_65),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_94),
.B1(n_76),
.B2(n_74),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_111),
.B1(n_3),
.B2(n_8),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_106),
.A2(n_58),
.B1(n_53),
.B2(n_57),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_55),
.Y(n_128)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_120),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_73),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_72),
.B1(n_66),
.B2(n_52),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_51),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_126),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_128),
.B(n_130),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_123),
.C(n_116),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_12),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_119),
.B1(n_118),
.B2(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_136),
.B1(n_13),
.B2(n_14),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_141),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_144),
.B(n_146),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_35),
.B1(n_44),
.B2(n_21),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_SL g151 ( 
.A(n_148),
.B(n_129),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_152)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_128),
.B1(n_132),
.B2(n_147),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_131),
.C(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_138),
.Y(n_157)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_127),
.B(n_14),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_127),
.B(n_13),
.Y(n_159)
);

OAI21x1_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_22),
.B(n_23),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_31),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_163)
);


endmodule