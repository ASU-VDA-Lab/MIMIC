module fake_jpeg_21625_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx4f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_19),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_18),
.A2(n_2),
.B(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_5),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_30),
.B1(n_29),
.B2(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_9),
.Y(n_30)
);

NAND2x1p5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_22),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

NOR3xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_13),
.C(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_25),
.C(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_41),
.C(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_33),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.C(n_40),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_33),
.C(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_39),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_43),
.Y(n_51)
);

XNOR2x2_ASAP7_75t_SL g52 ( 
.A(n_51),
.B(n_45),
.Y(n_52)
);


endmodule