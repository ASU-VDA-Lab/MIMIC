module fake_jpeg_233_n_497 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_497);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_497;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_41),
.B(n_49),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_42),
.B(n_43),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_47),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_48),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_13),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_51),
.B(n_64),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_13),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_53),
.B(n_62),
.Y(n_115)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_13),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g121 ( 
.A(n_65),
.Y(n_121)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_30),
.B(n_13),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_80),
.Y(n_119)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_82),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_23),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_12),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_11),
.Y(n_132)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_87),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_95),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_33),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_65),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_105),
.B(n_132),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_35),
.B1(n_23),
.B2(n_20),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_110),
.A2(n_123),
.B1(n_56),
.B2(n_81),
.Y(n_176)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_28),
.C(n_34),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_145),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_35),
.B1(n_15),
.B2(n_31),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_45),
.A2(n_34),
.B1(n_33),
.B2(n_31),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_126),
.A2(n_83),
.B1(n_39),
.B2(n_14),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_84),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_48),
.A2(n_33),
.B(n_31),
.C(n_15),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_136),
.A2(n_87),
.B1(n_59),
.B2(n_78),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_46),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_15),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_55),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_63),
.B(n_24),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_153),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_63),
.B(n_24),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_126),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_76),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_162),
.Y(n_218)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_104),
.A2(n_96),
.B1(n_92),
.B2(n_86),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_161),
.B(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_0),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_101),
.B(n_0),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_178),
.Y(n_222)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_110),
.A2(n_60),
.B1(n_66),
.B2(n_74),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_169),
.A2(n_187),
.B(n_189),
.C(n_124),
.Y(n_230)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_180),
.B1(n_188),
.B2(n_194),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_95),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_0),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_116),
.B(n_89),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_127),
.C(n_122),
.Y(n_217)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_89),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_185),
.Y(n_199)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_192),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_123),
.A2(n_73),
.B1(n_67),
.B2(n_57),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_117),
.A2(n_52),
.B1(n_68),
.B2(n_50),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_141),
.A2(n_24),
.B1(n_79),
.B2(n_70),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_99),
.B1(n_142),
.B2(n_139),
.Y(n_210)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_195),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_120),
.A2(n_84),
.B1(n_79),
.B2(n_70),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_12),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_196),
.Y(n_204)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_111),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_198),
.Y(n_224)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_149),
.B1(n_137),
.B2(n_103),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_187),
.B1(n_169),
.B2(n_190),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_225),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_227),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_228),
.B(n_220),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_159),
.B(n_158),
.Y(n_225)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_170),
.A2(n_106),
.B1(n_114),
.B2(n_122),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_118),
.C(n_146),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_182),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_166),
.B(n_137),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_175),
.Y(n_257)
);

BUFx4f_ASAP7_75t_SL g252 ( 
.A(n_230),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_232),
.B(n_234),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_201),
.B(n_162),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_233),
.B(n_235),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_222),
.B(n_167),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_242),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_237),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_243),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_207),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_247),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_191),
.B1(n_172),
.B2(n_178),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_246),
.A2(n_258),
.B1(n_202),
.B2(n_208),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_222),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_253),
.B(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_251),
.A2(n_209),
.B1(n_221),
.B2(n_165),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_161),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_182),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_254),
.A2(n_229),
.B(n_210),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_199),
.B(n_181),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_220),
.A2(n_103),
.B1(n_149),
.B2(n_150),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_236),
.B1(n_227),
.B2(n_258),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_208),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_205),
.A2(n_171),
.B1(n_160),
.B2(n_164),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_217),
.B(n_219),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_262),
.A2(n_265),
.B(n_279),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_218),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_267),
.C(n_281),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_244),
.A2(n_230),
.B(n_210),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_250),
.B(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_268),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_244),
.A2(n_230),
.B1(n_204),
.B2(n_210),
.Y(n_270)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_278),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_246),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_253),
.A2(n_230),
.B1(n_221),
.B2(n_196),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_214),
.B(n_163),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_214),
.B(n_124),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_238),
.B(n_234),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_192),
.C(n_197),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_283),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_272),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_285),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_288),
.A2(n_295),
.B(n_283),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_272),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_297),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_284),
.Y(n_290)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_232),
.Y(n_291)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_269),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_284),
.Y(n_297)
);

OA22x2_ASAP7_75t_L g298 ( 
.A1(n_273),
.A2(n_236),
.B1(n_254),
.B2(n_252),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_SL g326 ( 
.A1(n_298),
.A2(n_265),
.B(n_254),
.C(n_252),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_279),
.Y(n_299)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_255),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_302),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_239),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_264),
.B(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_274),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_306),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_260),
.B(n_247),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_248),
.Y(n_307)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_307),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_257),
.Y(n_308)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_308),
.Y(n_335)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_251),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_245),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_242),
.Y(n_311)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_311),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_297),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_314),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_286),
.A2(n_278),
.B1(n_256),
.B2(n_252),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_313),
.A2(n_309),
.B1(n_301),
.B2(n_306),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_302),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_262),
.B(n_280),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_323),
.B(n_326),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_259),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_320),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_285),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_333),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_259),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_300),
.A2(n_277),
.B(n_276),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_328),
.A2(n_288),
.B(n_299),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_332),
.B(n_336),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_289),
.Y(n_333)
);

AO21x2_ASAP7_75t_L g334 ( 
.A1(n_287),
.A2(n_252),
.B(n_258),
.Y(n_334)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_294),
.B(n_267),
.CI(n_263),
.CON(n_336),
.SN(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_267),
.C(n_281),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_320),
.C(n_316),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_329),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_345),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_328),
.Y(n_378)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_321),
.A2(n_287),
.B1(n_290),
.B2(n_304),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_346),
.A2(n_349),
.B1(n_361),
.B2(n_350),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_293),
.B(n_300),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_348),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_329),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_321),
.A2(n_295),
.B1(n_303),
.B2(n_305),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_339),
.Y(n_350)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_288),
.C(n_292),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_342),
.C(n_359),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_325),
.A2(n_303),
.B1(n_252),
.B2(n_307),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_355),
.A2(n_358),
.B1(n_366),
.B2(n_317),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_331),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_363),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_341),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_325),
.A2(n_311),
.B1(n_286),
.B2(n_291),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_308),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_360),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_335),
.B(n_264),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_339),
.A2(n_293),
.B1(n_298),
.B2(n_311),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_362),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_235),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_330),
.Y(n_364)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_364),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_293),
.B(n_286),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_365),
.B(n_334),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_368),
.A2(n_375),
.B(n_374),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_369),
.A2(n_344),
.B(n_327),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_345),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_371),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_322),
.Y(n_373)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_373),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_233),
.Y(n_377)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_377),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_378),
.B(n_381),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_298),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_380),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_298),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_383),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_317),
.C(n_335),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_385),
.C(n_386),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_330),
.C(n_282),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_352),
.B(n_298),
.C(n_336),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_387),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_352),
.B(n_298),
.C(n_336),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_392),
.Y(n_404)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_390),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_353),
.B(n_296),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_391),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_326),
.Y(n_392)
);

BUFx12_ASAP7_75t_L g395 ( 
.A(n_379),
.Y(n_395)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_395),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_388),
.A2(n_390),
.B1(n_373),
.B2(n_370),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_397),
.A2(n_399),
.B1(n_409),
.B2(n_415),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_382),
.A2(n_344),
.B1(n_355),
.B2(n_334),
.Y(n_399)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_403),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_406),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_SL g406 ( 
.A(n_386),
.B(n_361),
.C(n_347),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_368),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_407),
.B(n_396),
.Y(n_430)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_408),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_353),
.B1(n_334),
.B2(n_365),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_384),
.A2(n_346),
.B(n_349),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_413),
.B(n_392),
.Y(n_429)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_414),
.B(n_381),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_418),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_378),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_410),
.B(n_360),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_423),
.Y(n_446)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_398),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_434),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_400),
.B(n_296),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_380),
.C(n_389),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_432),
.C(n_395),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_271),
.Y(n_425)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_415),
.Y(n_426)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_429),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_430),
.A2(n_402),
.B1(n_405),
.B2(n_394),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_413),
.A2(n_376),
.B(n_326),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_431),
.A2(n_402),
.B1(n_411),
.B2(n_326),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_376),
.C(n_362),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_334),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_399),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_401),
.B(n_310),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_419),
.Y(n_435)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

NAND2x1_ASAP7_75t_SL g453 ( 
.A(n_436),
.B(n_429),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_394),
.C(n_408),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_447),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_404),
.Y(n_439)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_441),
.A2(n_443),
.B1(n_427),
.B2(n_420),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_139),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_428),
.A2(n_327),
.B1(n_401),
.B2(n_406),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_203),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_395),
.C(n_275),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_275),
.C(n_240),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_448),
.B(n_179),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_452),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_455),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_432),
.C(n_433),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_446),
.A2(n_403),
.B(n_241),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_456),
.A2(n_457),
.B(n_459),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_439),
.A2(n_211),
.B(n_215),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_447),
.B(n_211),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_458),
.B(n_448),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_445),
.A2(n_183),
.B(n_193),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_463),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_464),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_440),
.A2(n_152),
.B1(n_129),
.B2(n_108),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_462),
.B(n_449),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_467),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_SL g468 ( 
.A1(n_454),
.A2(n_436),
.B1(n_437),
.B2(n_450),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_468),
.A2(n_144),
.B(n_152),
.Y(n_479)
);

INVx11_ASAP7_75t_L g469 ( 
.A(n_451),
.Y(n_469)
);

AOI31xp33_ASAP7_75t_L g482 ( 
.A1(n_469),
.A2(n_173),
.A3(n_100),
.B(n_144),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_453),
.A2(n_435),
.B(n_203),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_470),
.A2(n_97),
.B(n_150),
.Y(n_478)
);

AOI221xp5_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_202),
.B1(n_198),
.B2(n_124),
.C(n_168),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_471),
.A2(n_114),
.B1(n_185),
.B2(n_97),
.Y(n_477)
);

O2A1O1Ixp33_ASAP7_75t_SL g476 ( 
.A1(n_466),
.A2(n_461),
.B(n_464),
.C(n_186),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_476),
.A2(n_478),
.B(n_479),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_477),
.B(n_481),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_473),
.A2(n_129),
.B(n_108),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_SL g488 ( 
.A1(n_482),
.A2(n_483),
.B(n_12),
.C(n_10),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_39),
.C(n_113),
.Y(n_483)
);

AOI322xp5_ASAP7_75t_L g484 ( 
.A1(n_480),
.A2(n_472),
.A3(n_474),
.B1(n_475),
.B2(n_471),
.C1(n_39),
.C2(n_113),
.Y(n_484)
);

OAI311xp33_ASAP7_75t_L g492 ( 
.A1(n_484),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.C1(n_4),
.Y(n_492)
);

OAI221xp5_ASAP7_75t_L g487 ( 
.A1(n_477),
.A2(n_113),
.B1(n_12),
.B2(n_11),
.C(n_10),
.Y(n_487)
);

NOR3xp33_ASAP7_75t_L g491 ( 
.A(n_487),
.B(n_488),
.C(n_489),
.Y(n_491)
);

OAI331xp33_ASAP7_75t_L g489 ( 
.A1(n_480),
.A2(n_10),
.A3(n_9),
.B1(n_2),
.B2(n_3),
.B3(n_0),
.C1(n_5),
.Y(n_489)
);

AOI21x1_ASAP7_75t_L g490 ( 
.A1(n_486),
.A2(n_1),
.B(n_2),
.Y(n_490)
);

NOR3xp33_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_485),
.C(n_491),
.Y(n_493)
);

O2A1O1Ixp33_ASAP7_75t_SL g494 ( 
.A1(n_492),
.A2(n_5),
.B(n_1),
.C(n_4),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_493),
.A2(n_494),
.B(n_4),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_495),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_496),
.B(n_5),
.Y(n_497)
);


endmodule