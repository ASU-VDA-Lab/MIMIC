module fake_ariane_2546_n_1883 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1883);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1883;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g180 ( 
.A(n_12),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_18),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_106),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_7),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_74),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_56),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_43),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_41),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_103),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_78),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_29),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_12),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_137),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_51),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_14),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_50),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_58),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_87),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_66),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_27),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_95),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_16),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_99),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_81),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_76),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_92),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_63),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_46),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_174),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_56),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_128),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_39),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_8),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_48),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_110),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_97),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_104),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_79),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_154),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_88),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_86),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_123),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_80),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_2),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_47),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_126),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_127),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_35),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_131),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_161),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_146),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_120),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_54),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_11),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_133),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_165),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_33),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_19),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_144),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_61),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_7),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_89),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_54),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_148),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_27),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_130),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_72),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_57),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_141),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_16),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_132),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_17),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_41),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_107),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_31),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_136),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_39),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_85),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_26),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_11),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_34),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_57),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_28),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_37),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_67),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_176),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_18),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_142),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_14),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_102),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_162),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_159),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_153),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_167),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_117),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_114),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_82),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_172),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_94),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_6),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_101),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_48),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_145),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_118),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_108),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_36),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_17),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_24),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_29),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_52),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_15),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_45),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_60),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_5),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_175),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_98),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_19),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_71),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_77),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_112),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_63),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_38),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_179),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_53),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_46),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_96),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_8),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_21),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_138),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_36),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_49),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_49),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_134),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_42),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_155),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_1),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_22),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_35),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_171),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_70),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_121),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_119),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_60),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_170),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_23),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_3),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_31),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_166),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_152),
.Y(n_350)
);

BUFx8_ASAP7_75t_SL g351 ( 
.A(n_25),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_158),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_169),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_75),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_34),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_50),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_149),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_24),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_30),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_3),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_190),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_194),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_211),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_211),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_190),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_199),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_257),
.B(n_0),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_199),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_200),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_351),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_200),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_204),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_184),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_208),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_204),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_255),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_266),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_276),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_206),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_306),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_316),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_322),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_206),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_224),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_343),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_224),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_181),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_231),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_231),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_322),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_183),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_232),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_257),
.B(n_0),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_277),
.B(n_1),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_210),
.B(n_4),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_254),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_232),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_186),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_301),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_233),
.B(n_4),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_185),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_241),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_253),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_187),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_188),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_233),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_239),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_239),
.B(n_9),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_337),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_243),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_194),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_243),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_191),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_249),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_249),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_193),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_197),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_252),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_322),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_252),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_256),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_205),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_207),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_256),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_220),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_294),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_202),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_277),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_209),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_294),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_300),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_227),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_216),
.B(n_10),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_309),
.B(n_10),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_322),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_300),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_228),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_322),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_321),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_321),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_244),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_245),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_248),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_202),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_335),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_202),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_323),
.B(n_13),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_180),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_251),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_324),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_324),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_258),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_336),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_383),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_336),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_R g459 ( 
.A(n_388),
.B(n_182),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_361),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_392),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_361),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_405),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_374),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_377),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_366),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_366),
.B(n_348),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_367),
.B(n_342),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_402),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_403),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_367),
.B(n_348),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_381),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_404),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_369),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_411),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_R g479 ( 
.A(n_399),
.B(n_189),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_386),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_369),
.B(n_202),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_431),
.B(n_342),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_370),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_375),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_370),
.B(n_349),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_372),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_378),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_362),
.B(n_278),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_379),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_372),
.B(n_349),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_373),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_382),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_437),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_371),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_406),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_415),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_362),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_373),
.B(n_278),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_418),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_376),
.B(n_278),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_437),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_376),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_440),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_380),
.B(n_323),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_380),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_447),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_419),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_384),
.B(n_265),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_447),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_384),
.B(n_357),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_385),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_385),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_387),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_387),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_389),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_389),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_390),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_424),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_393),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_393),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_398),
.B(n_278),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_398),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_408),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_409),
.A2(n_357),
.B(n_246),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_499),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_460),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_521),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_481),
.B(n_436),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_456),
.B(n_363),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_482),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_L g541 ( 
.A(n_521),
.B(n_459),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_488),
.A2(n_435),
.B1(n_396),
.B2(n_450),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_521),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_460),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_456),
.B(n_364),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_461),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_481),
.B(n_500),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_521),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_463),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_482),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_529),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g553 ( 
.A(n_481),
.B(n_436),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_500),
.A2(n_443),
.B1(n_444),
.B2(n_439),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_470),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_482),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_458),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_500),
.A2(n_451),
.B1(n_454),
.B2(n_445),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_534),
.A2(n_414),
.B1(n_416),
.B2(n_412),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_467),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_521),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_521),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_488),
.B(n_407),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_467),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_502),
.B(n_412),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_502),
.B(n_414),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_458),
.B(n_416),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_477),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_508),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_505),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_505),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_477),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_484),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_417),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_527),
.B(n_417),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_462),
.Y(n_577)
);

NAND2x1p5_ASAP7_75t_L g578 ( 
.A(n_527),
.B(n_394),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_471),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_484),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_519),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_527),
.B(n_420),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_469),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_508),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_487),
.B(n_420),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_487),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_493),
.B(n_504),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_493),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_512),
.B(n_215),
.Y(n_589)
);

INVx4_ASAP7_75t_L g590 ( 
.A(n_508),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_479),
.B(n_504),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_529),
.B(n_430),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_508),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_468),
.B(n_394),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_509),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_534),
.A2(n_455),
.B1(n_453),
.B2(n_452),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_507),
.B(n_430),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_507),
.B(n_429),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_490),
.A2(n_410),
.B1(n_401),
.B2(n_395),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_469),
.A2(n_395),
.B1(n_449),
.B2(n_368),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_515),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_516),
.B(n_422),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_468),
.B(n_423),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_462),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_516),
.B(n_423),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_464),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_464),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_462),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_497),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_498),
.A2(n_223),
.B1(n_282),
.B2(n_260),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_501),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_511),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_534),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_517),
.B(n_215),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_468),
.B(n_426),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_462),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_525),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_462),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_517),
.B(n_426),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_525),
.B(n_446),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_518),
.B(n_246),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_518),
.B(n_428),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_465),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_464),
.Y(n_627)
);

BUFx8_ASAP7_75t_SL g628 ( 
.A(n_496),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_520),
.B(n_523),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_520),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_523),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_524),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_522),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_466),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_528),
.B(n_448),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_528),
.A2(n_284),
.B1(n_310),
.B2(n_329),
.Y(n_636)
);

INVx4_ASAP7_75t_SL g637 ( 
.A(n_462),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_524),
.B(n_428),
.Y(n_638)
);

AO22x2_ASAP7_75t_L g639 ( 
.A1(n_486),
.A2(n_441),
.B1(n_453),
.B2(n_452),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_526),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_473),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_472),
.B(n_365),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_475),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_530),
.Y(n_644)
);

BUFx4f_ASAP7_75t_L g645 ( 
.A(n_534),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_475),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_L g647 ( 
.A(n_457),
.B(n_433),
.C(n_432),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_530),
.B(n_433),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_476),
.B(n_438),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_532),
.B(n_438),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_532),
.B(n_533),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_512),
.B(n_274),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_533),
.B(n_335),
.Y(n_653)
);

BUFx6f_ASAP7_75t_SL g654 ( 
.A(n_512),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_519),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_519),
.B(n_441),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_480),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_534),
.A2(n_455),
.B1(n_442),
.B2(n_180),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_476),
.B(n_442),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_531),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_475),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_462),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_531),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_531),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_512),
.Y(n_665)
);

INVx6_ASAP7_75t_L g666 ( 
.A(n_472),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_472),
.Y(n_667)
);

AND2x6_ASAP7_75t_L g668 ( 
.A(n_486),
.B(n_274),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_492),
.B(n_285),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_475),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_485),
.B(n_196),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_492),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_514),
.A2(n_219),
.B1(n_226),
.B2(n_214),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_503),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_514),
.A2(n_219),
.B1(n_226),
.B2(n_214),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_489),
.B(n_341),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_503),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_457),
.B(n_483),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_503),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_503),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_483),
.B(n_295),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_510),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_494),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_510),
.B(n_299),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_510),
.B(n_495),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_540),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_592),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_540),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_553),
.B(n_309),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_626),
.B(n_491),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_660),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_551),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_SL g693 ( 
.A(n_626),
.B(n_268),
.C(n_261),
.Y(n_693)
);

BUFx6f_ASAP7_75t_SL g694 ( 
.A(n_641),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_583),
.B(n_510),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_628),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_576),
.B(n_582),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_663),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_619),
.B(n_474),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_551),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_576),
.B(n_196),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_582),
.B(n_198),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_553),
.B(n_555),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_666),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_678),
.B(n_198),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_664),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_557),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_L g708 ( 
.A(n_543),
.B(n_203),
.C(n_201),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_559),
.B(n_309),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_672),
.B(n_201),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_571),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_548),
.B(n_566),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_567),
.B(n_203),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_641),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_549),
.B(n_335),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_666),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_574),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_591),
.B(n_478),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_575),
.B(n_213),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_681),
.B(n_213),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_558),
.B(n_240),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_558),
.B(n_240),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_581),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_543),
.A2(n_264),
.B1(n_288),
.B2(n_286),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_552),
.B(n_270),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_556),
.B(n_263),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_587),
.A2(n_506),
.B(n_495),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_591),
.B(n_272),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_574),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_604),
.B(n_263),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_581),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_604),
.B(n_280),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_604),
.B(n_280),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_617),
.B(n_287),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_617),
.B(n_287),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_611),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_666),
.B(n_273),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_655),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_614),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_617),
.B(n_312),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_570),
.B(n_312),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_594),
.A2(n_341),
.B1(n_335),
.B2(n_265),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_538),
.B(n_275),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_549),
.B(n_335),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_655),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_570),
.B(n_279),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_584),
.B(n_313),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_676),
.B(n_341),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_538),
.B(n_281),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_584),
.B(n_313),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_571),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_572),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_590),
.B(n_326),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_578),
.B(n_332),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_613),
.B(n_633),
.C(n_657),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_649),
.B(n_332),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_578),
.B(n_283),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_593),
.B(n_289),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_593),
.B(n_339),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_671),
.B(n_292),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_568),
.B(n_339),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_SL g762 ( 
.A(n_536),
.B(n_347),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_568),
.B(n_347),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_634),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_649),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_612),
.B(n_307),
.C(n_360),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_594),
.B(n_303),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_594),
.B(n_308),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_545),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_572),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_564),
.B(n_314),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_550),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_554),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_561),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_601),
.B(n_315),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_565),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_601),
.B(n_318),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_537),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_603),
.B(n_325),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_634),
.B(n_600),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_603),
.B(n_328),
.Y(n_781)
);

OAI221xp5_ASAP7_75t_L g782 ( 
.A1(n_673),
.A2(n_331),
.B1(n_359),
.B2(n_358),
.C(n_356),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_589),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_639),
.A2(n_341),
.B1(n_335),
.B2(n_265),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_639),
.A2(n_355),
.B1(n_265),
.B2(n_238),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_634),
.B(n_333),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_649),
.B(n_338),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_621),
.B(n_344),
.Y(n_788)
);

AOI221xp5_ASAP7_75t_L g789 ( 
.A1(n_673),
.A2(n_346),
.B1(n_355),
.B2(n_265),
.C(n_302),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_642),
.B(n_192),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_638),
.B(n_195),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_607),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_659),
.B(n_13),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_607),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_598),
.B(n_212),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_638),
.B(n_217),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_665),
.B(n_218),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_650),
.B(n_221),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_667),
.B(n_355),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_608),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_650),
.B(n_222),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_665),
.B(n_225),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_539),
.B(n_229),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_636),
.A2(n_355),
.B1(n_238),
.B2(n_209),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_539),
.B(n_546),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_546),
.B(n_651),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_651),
.B(n_230),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_639),
.B(n_355),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_599),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_659),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_569),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_573),
.Y(n_812)
);

OAI22x1_ASAP7_75t_SL g813 ( 
.A1(n_683),
.A2(n_340),
.B1(n_259),
.B2(n_250),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_647),
.B(n_235),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_580),
.B(n_236),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_586),
.B(n_237),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_659),
.B(n_242),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_628),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_588),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_585),
.B(n_247),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_595),
.B(n_262),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_606),
.B(n_625),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_596),
.B(n_267),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_648),
.B(n_269),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_535),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_549),
.B(n_234),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_675),
.B(n_319),
.C(n_271),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_675),
.B(n_290),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_602),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_645),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_630),
.B(n_631),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_632),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_645),
.A2(n_296),
.B1(n_334),
.B2(n_285),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_654),
.B(n_291),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_589),
.A2(n_327),
.B1(n_293),
.B2(n_304),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_640),
.B(n_297),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_644),
.B(n_298),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_683),
.B(n_305),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_560),
.B(n_317),
.Y(n_839)
);

CKINVDCx11_ASAP7_75t_R g840 ( 
.A(n_579),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_608),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_560),
.B(n_320),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_629),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_547),
.B(n_15),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_597),
.B(n_350),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_597),
.B(n_352),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_622),
.B(n_345),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_654),
.B(n_330),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_697),
.A2(n_541),
.B(n_537),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_806),
.A2(n_541),
.B(n_563),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_805),
.B(n_589),
.Y(n_851)
);

CKINVDCx6p67_ASAP7_75t_R g852 ( 
.A(n_694),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_783),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_727),
.A2(n_680),
.B(n_623),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_714),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_703),
.A2(n_658),
.B1(n_668),
.B2(n_669),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_769),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_712),
.A2(n_615),
.B(n_685),
.Y(n_858)
);

NOR3xp33_ASAP7_75t_L g859 ( 
.A(n_699),
.B(n_635),
.C(n_656),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_783),
.Y(n_860)
);

CKINVDCx10_ASAP7_75t_R g861 ( 
.A(n_694),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_843),
.B(n_615),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_686),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_843),
.A2(n_841),
.B(n_800),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_704),
.B(n_670),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_687),
.B(n_579),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_803),
.B(n_589),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_704),
.B(n_679),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_779),
.B(n_781),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_830),
.B(n_549),
.Y(n_870)
);

O2A1O1Ixp5_ASAP7_75t_L g871 ( 
.A1(n_762),
.A2(n_822),
.B(n_702),
.C(n_701),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_788),
.B(n_705),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_785),
.A2(n_658),
.B1(n_668),
.B2(n_669),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_765),
.B(n_652),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_771),
.B(n_754),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_760),
.B(n_679),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_754),
.B(n_652),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_695),
.A2(n_563),
.B(n_562),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_769),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_716),
.B(n_684),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_831),
.A2(n_562),
.B(n_544),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_686),
.Y(n_882)
);

OAI321xp33_ASAP7_75t_L g883 ( 
.A1(n_724),
.A2(n_804),
.A3(n_782),
.B1(n_789),
.B2(n_784),
.C(n_777),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_688),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_762),
.A2(n_616),
.B(n_623),
.C(n_677),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_688),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_SL g887 ( 
.A1(n_780),
.A2(n_616),
.B(n_302),
.C(n_353),
.Y(n_887)
);

OAI321xp33_ASAP7_75t_L g888 ( 
.A1(n_775),
.A2(n_761),
.A3(n_763),
.B1(n_809),
.B2(n_728),
.C(n_720),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_689),
.B(n_609),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_717),
.A2(n_682),
.B1(n_677),
.B2(n_674),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_810),
.B(n_637),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_783),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_810),
.B(n_624),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_748),
.B(n_624),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_708),
.A2(n_682),
.B(n_674),
.C(n_661),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_723),
.A2(n_542),
.B(n_627),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_772),
.B(n_668),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_717),
.B(n_542),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_718),
.B(n_627),
.Y(n_899)
);

AOI21x1_ASAP7_75t_L g900 ( 
.A1(n_839),
.A2(n_661),
.B(n_646),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_772),
.B(n_669),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_717),
.A2(n_643),
.B1(n_646),
.B2(n_542),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_731),
.A2(n_643),
.B(n_662),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_773),
.B(n_669),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_736),
.B(n_653),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_800),
.A2(n_610),
.B(n_653),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_773),
.B(n_577),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_731),
.A2(n_662),
.B(n_577),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_774),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_692),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_774),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_776),
.B(n_811),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_729),
.A2(n_662),
.B1(n_620),
.B2(n_618),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_738),
.A2(n_662),
.B(n_577),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_714),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_726),
.B(n_20),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_776),
.A2(n_353),
.B(n_296),
.C(n_334),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_755),
.B(n_577),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_807),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_738),
.A2(n_620),
.B(n_618),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_790),
.A2(n_749),
.B1(n_743),
.B2(n_757),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_729),
.A2(n_620),
.B1(n_618),
.B2(n_605),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_791),
.A2(n_23),
.B(n_26),
.C(n_28),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_745),
.A2(n_620),
.B(n_618),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_690),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_842),
.A2(n_637),
.B(n_605),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_811),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_700),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_812),
.B(n_605),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_737),
.A2(n_605),
.B1(n_354),
.B2(n_637),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_707),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_812),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_739),
.B(n_495),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_745),
.A2(n_610),
.B(n_234),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_819),
.B(n_829),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_819),
.B(n_513),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_829),
.Y(n_937)
);

OAI321xp33_ASAP7_75t_L g938 ( 
.A1(n_827),
.A2(n_513),
.A3(n_506),
.B1(n_495),
.B2(n_234),
.C(n_42),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_778),
.A2(n_506),
.B(n_495),
.Y(n_939)
);

AND2x2_ASAP7_75t_SL g940 ( 
.A(n_808),
.B(n_513),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_691),
.A2(n_706),
.B(n_698),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_729),
.A2(n_506),
.B1(n_495),
.B2(n_513),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_832),
.B(n_513),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_832),
.A2(n_706),
.B(n_698),
.C(n_801),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_799),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_766),
.A2(n_513),
.B1(n_32),
.B2(n_33),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_799),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_796),
.A2(n_30),
.B(n_40),
.C(n_43),
.Y(n_948)
);

O2A1O1Ixp5_ASAP7_75t_L g949 ( 
.A1(n_710),
.A2(n_40),
.B(n_44),
.C(n_45),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_764),
.Y(n_950)
);

O2A1O1Ixp5_ASAP7_75t_L g951 ( 
.A1(n_845),
.A2(n_52),
.B(n_53),
.C(n_55),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_793),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_707),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_798),
.A2(n_100),
.B(n_157),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_815),
.A2(n_93),
.B(n_151),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_795),
.B(n_55),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_793),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_721),
.B(n_58),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_SL g959 ( 
.A(n_696),
.B(n_59),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_817),
.A2(n_59),
.B1(n_62),
.B2(n_64),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_722),
.B(n_62),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_741),
.A2(n_64),
.B(n_65),
.C(n_68),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_726),
.B(n_65),
.Y(n_963)
);

NOR2x1_ASAP7_75t_L g964 ( 
.A(n_764),
.B(n_69),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_711),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_816),
.A2(n_73),
.B(n_83),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_747),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_750),
.A2(n_84),
.B1(n_90),
.B2(n_91),
.Y(n_968)
);

OA22x2_ASAP7_75t_L g969 ( 
.A1(n_847),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_828),
.A2(n_116),
.B1(n_124),
.B2(n_125),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_840),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_835),
.B(n_129),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_821),
.A2(n_140),
.B(n_143),
.Y(n_973)
);

AO22x1_ASAP7_75t_L g974 ( 
.A1(n_696),
.A2(n_147),
.B1(n_177),
.B2(n_818),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_709),
.A2(n_725),
.B1(n_768),
.B2(n_767),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_711),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_753),
.A2(n_759),
.B(n_719),
.C(n_713),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_730),
.B(n_734),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_751),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_756),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_751),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_840),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_732),
.A2(n_740),
.B(n_733),
.C(n_735),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_834),
.B(n_848),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_823),
.A2(n_837),
.B(n_836),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_825),
.B(n_814),
.C(n_787),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_797),
.A2(n_802),
.B(n_824),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_756),
.B(n_787),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_752),
.A2(n_794),
.B(n_792),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_820),
.A2(n_758),
.B(n_746),
.Y(n_990)
);

O2A1O1Ixp5_ASAP7_75t_L g991 ( 
.A1(n_846),
.A2(n_794),
.B(n_770),
.C(n_792),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_770),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_808),
.A2(n_833),
.B1(n_742),
.B2(n_693),
.Y(n_993)
);

OA22x2_ASAP7_75t_L g994 ( 
.A1(n_838),
.A2(n_786),
.B1(n_813),
.B2(n_818),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_826),
.A2(n_715),
.B(n_744),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_844),
.B(n_694),
.Y(n_996)
);

OAI321xp33_ASAP7_75t_L g997 ( 
.A1(n_844),
.A2(n_543),
.A3(n_805),
.B1(n_601),
.B2(n_724),
.C(n_600),
.Y(n_997)
);

OA21x2_ASAP7_75t_L g998 ( 
.A1(n_727),
.A2(n_698),
.B(n_691),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_697),
.A2(n_806),
.B(n_712),
.Y(n_999)
);

OA21x2_ASAP7_75t_L g1000 ( 
.A1(n_727),
.A2(n_698),
.B(n_691),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_697),
.A2(n_806),
.B(n_712),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_769),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_697),
.A2(n_806),
.B(n_712),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_687),
.B(n_556),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_783),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_697),
.A2(n_806),
.B(n_712),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_825),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_687),
.B(n_592),
.Y(n_1008)
);

O2A1O1Ixp5_ASAP7_75t_L g1009 ( 
.A1(n_697),
.A2(n_762),
.B(n_822),
.C(n_806),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_805),
.B(n_697),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_697),
.A2(n_806),
.B(n_712),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_805),
.B(n_697),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_697),
.A2(n_806),
.B(n_712),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_805),
.A2(n_703),
.B1(n_785),
.B2(n_553),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_697),
.A2(n_806),
.B(n_712),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_697),
.B(n_703),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_697),
.B(n_830),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_SL g1018 ( 
.A1(n_697),
.A2(n_806),
.B(n_780),
.C(n_702),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_697),
.A2(n_806),
.B(n_712),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_840),
.Y(n_1020)
);

INVxp67_ASAP7_75t_SL g1021 ( 
.A(n_912),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_1016),
.B(n_921),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_991),
.A2(n_926),
.B(n_900),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1016),
.B(n_875),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_872),
.B(n_1006),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_991),
.A2(n_989),
.B(n_854),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1014),
.A2(n_859),
.B1(n_1008),
.B2(n_866),
.Y(n_1028)
);

AO31x2_ASAP7_75t_L g1029 ( 
.A1(n_944),
.A2(n_862),
.A3(n_941),
.B(n_1011),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_908),
.A2(n_920),
.B(n_914),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_1013),
.B(n_1015),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_1019),
.A2(n_1018),
.B(n_985),
.Y(n_1032)
);

OAI22x1_ASAP7_75t_L g1033 ( 
.A1(n_963),
.A2(n_956),
.B1(n_925),
.B2(n_952),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_924),
.A2(n_903),
.B(n_864),
.Y(n_1034)
);

BUFx2_ASAP7_75t_L g1035 ( 
.A(n_1007),
.Y(n_1035)
);

OR2x6_ASAP7_75t_L g1036 ( 
.A(n_925),
.B(n_980),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_869),
.B(n_984),
.Y(n_1037)
);

INVxp67_ASAP7_75t_L g1038 ( 
.A(n_1004),
.Y(n_1038)
);

AOI21x1_ASAP7_75t_L g1039 ( 
.A1(n_1017),
.A2(n_972),
.B(n_995),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_978),
.B(n_967),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1014),
.A2(n_859),
.B1(n_988),
.B2(n_956),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_899),
.B(n_876),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_952),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_855),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1018),
.A2(n_850),
.B(n_858),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_939),
.A2(n_896),
.B(n_849),
.Y(n_1046)
);

AO31x2_ASAP7_75t_L g1047 ( 
.A1(n_862),
.A2(n_901),
.A3(n_904),
.B(n_897),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_R g1048 ( 
.A(n_861),
.B(n_1020),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_957),
.B(n_916),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_899),
.B(n_935),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1009),
.A2(n_977),
.B(n_851),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_934),
.A2(n_913),
.B(n_922),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1009),
.A2(n_871),
.B(n_885),
.Y(n_1053)
);

AOI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_997),
.A2(n_888),
.B(n_883),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_871),
.A2(n_960),
.B(n_983),
.C(n_949),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_857),
.B(n_879),
.Y(n_1056)
);

BUFx12f_ASAP7_75t_L g1057 ( 
.A(n_915),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_867),
.A2(n_929),
.B(n_907),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_891),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_906),
.A2(n_936),
.B(n_943),
.Y(n_1060)
);

AND2x6_ASAP7_75t_L g1061 ( 
.A(n_853),
.B(n_860),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_957),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_909),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_949),
.A2(n_946),
.B(n_919),
.C(n_948),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_891),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_905),
.B(n_994),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_870),
.A2(n_1000),
.B(n_998),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_994),
.B(n_996),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_852),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_998),
.A2(n_1000),
.B(n_878),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_853),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_950),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_863),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_998),
.A2(n_1000),
.B(n_890),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_881),
.A2(n_898),
.B(n_987),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_911),
.A2(n_927),
.B1(n_932),
.B2(n_1002),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_880),
.B(n_986),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_937),
.B(n_945),
.Y(n_1078)
);

AOI21x1_ASAP7_75t_L g1079 ( 
.A1(n_958),
.A2(n_961),
.B(n_990),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_882),
.Y(n_1080)
);

AO31x2_ASAP7_75t_L g1081 ( 
.A1(n_917),
.A2(n_889),
.A3(n_947),
.B(n_979),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_971),
.Y(n_1082)
);

OAI22x1_ASAP7_75t_L g1083 ( 
.A1(n_975),
.A2(n_982),
.B1(n_894),
.B2(n_893),
.Y(n_1083)
);

AOI221xp5_ASAP7_75t_L g1084 ( 
.A1(n_993),
.A2(n_938),
.B1(n_923),
.B2(n_959),
.C(n_951),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_993),
.A2(n_873),
.B1(n_940),
.B2(n_865),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_942),
.A2(n_902),
.B(n_895),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_SL g1087 ( 
.A(n_940),
.B(n_874),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_884),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_954),
.A2(n_973),
.B(n_966),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_877),
.B(n_894),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_886),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_873),
.A2(n_865),
.B1(n_868),
.B2(n_856),
.Y(n_1092)
);

AOI21x1_ASAP7_75t_SL g1093 ( 
.A1(n_951),
.A2(n_933),
.B(n_969),
.Y(n_1093)
);

NAND2x1p5_ASAP7_75t_L g1094 ( 
.A(n_853),
.B(n_1005),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_893),
.B(n_874),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_868),
.A2(n_955),
.B(n_887),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_953),
.B(n_965),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_887),
.A2(n_918),
.B(n_889),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_SL g1099 ( 
.A1(n_964),
.A2(n_856),
.B(n_970),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_853),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_962),
.A2(n_968),
.B(n_953),
.C(n_930),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_860),
.B(n_1005),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_910),
.A2(n_931),
.A3(n_992),
.B(n_928),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_860),
.B(n_892),
.Y(n_1104)
);

AOI221x1_ASAP7_75t_L g1105 ( 
.A1(n_981),
.A2(n_976),
.B1(n_969),
.B2(n_892),
.C(n_1005),
.Y(n_1105)
);

NOR2x1_ASAP7_75t_SL g1106 ( 
.A(n_892),
.B(n_1005),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_981),
.B(n_974),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_981),
.A2(n_1001),
.B(n_999),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_981),
.A2(n_1001),
.B(n_999),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_988),
.B(n_1008),
.Y(n_1110)
);

AND3x4_ASAP7_75t_L g1111 ( 
.A(n_859),
.B(n_714),
.C(n_755),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1010),
.A2(n_1012),
.B(n_1016),
.C(n_805),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_853),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1010),
.A2(n_1012),
.B(n_1009),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1016),
.B(n_921),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_855),
.B(n_915),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_857),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_857),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_857),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_891),
.Y(n_1125)
);

AO31x2_ASAP7_75t_L g1126 ( 
.A1(n_944),
.A2(n_862),
.A3(n_941),
.B(n_1016),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_991),
.A2(n_871),
.B(n_1009),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_891),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_SL g1129 ( 
.A1(n_941),
.A2(n_935),
.B(n_912),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_999),
.A2(n_1003),
.B(n_1001),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_L g1131 ( 
.A(n_1010),
.B(n_1012),
.C(n_997),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1010),
.A2(n_1012),
.B1(n_697),
.B2(n_921),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_863),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_SL g1137 ( 
.A1(n_1010),
.A2(n_1012),
.B(n_869),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_855),
.B(n_915),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1010),
.A2(n_1012),
.B(n_1009),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_891),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_853),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_853),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_857),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_SL g1144 ( 
.A(n_1020),
.B(n_714),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_900),
.A2(n_926),
.B(n_989),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_991),
.A2(n_926),
.B(n_900),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_855),
.Y(n_1148)
);

AND2x2_ASAP7_75t_SL g1149 ( 
.A(n_940),
.B(n_748),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_853),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_L g1151 ( 
.A(n_921),
.B(n_1012),
.C(n_1010),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_991),
.A2(n_926),
.B(n_900),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_991),
.A2(n_926),
.B(n_900),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_991),
.A2(n_926),
.B(n_900),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_988),
.B(n_1008),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_857),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1010),
.A2(n_1012),
.B(n_1016),
.C(n_805),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_991),
.A2(n_926),
.B(n_900),
.Y(n_1159)
);

AOI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_921),
.A2(n_803),
.B(n_760),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_999),
.A2(n_1003),
.B(n_1001),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_991),
.A2(n_926),
.B(n_900),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1163)
);

AOI21xp33_ASAP7_75t_L g1164 ( 
.A1(n_921),
.A2(n_803),
.B(n_760),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_863),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_863),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1010),
.A2(n_1012),
.B1(n_697),
.B2(n_921),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1063),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1057),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1119),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_1035),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1024),
.B(n_1120),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_1048),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1112),
.A2(n_1158),
.B1(n_1168),
.B2(n_1133),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1059),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1110),
.B(n_1155),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_SL g1178 ( 
.A1(n_1053),
.A2(n_1164),
.B(n_1160),
.C(n_1139),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1043),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1024),
.B(n_1120),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1131),
.A2(n_1054),
.B1(n_1149),
.B2(n_1041),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1048),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_1061),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1036),
.B(n_1059),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1065),
.B(n_1125),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1065),
.B(n_1125),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1128),
.B(n_1140),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1112),
.A2(n_1158),
.B(n_1115),
.Y(n_1188)
);

INVx3_ASAP7_75t_L g1189 ( 
.A(n_1113),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1131),
.B(n_1147),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_SL g1191 ( 
.A1(n_1151),
.A2(n_1111),
.B1(n_1028),
.B2(n_1147),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1073),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1128),
.B(n_1140),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1116),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1116),
.B(n_1138),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1113),
.Y(n_1196)
);

CKINVDCx6p67_ASAP7_75t_R g1197 ( 
.A(n_1069),
.Y(n_1197)
);

BUFx4_ASAP7_75t_SL g1198 ( 
.A(n_1036),
.Y(n_1198)
);

NAND2x1_ASAP7_75t_L g1199 ( 
.A(n_1061),
.B(n_1071),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1138),
.B(n_1036),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1123),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1095),
.B(n_1148),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1113),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1044),
.B(n_1043),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1066),
.B(n_1124),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1143),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1117),
.B(n_1118),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_1072),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1026),
.A2(n_1031),
.B(n_1130),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1049),
.B(n_1062),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1037),
.A2(n_1084),
.B(n_1022),
.C(n_1115),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1025),
.B(n_1050),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1157),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1022),
.A2(n_1122),
.B(n_1166),
.C(n_1163),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1080),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1121),
.A2(n_1135),
.B1(n_1132),
.B2(n_1156),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1136),
.B(n_1040),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1038),
.B(n_1042),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1038),
.B(n_1021),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1082),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1021),
.B(n_1077),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1056),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1068),
.B(n_1077),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1033),
.B(n_1078),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1083),
.B(n_1149),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_1061),
.Y(n_1226)
);

BUFx8_ASAP7_75t_SL g1227 ( 
.A(n_1113),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1111),
.Y(n_1228)
);

NAND3xp33_ASAP7_75t_L g1229 ( 
.A(n_1055),
.B(n_1064),
.C(n_1114),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1027),
.A2(n_1023),
.B(n_1152),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_1090),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1106),
.B(n_1100),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1141),
.Y(n_1233)
);

AOI21xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1076),
.A2(n_1107),
.B(n_1144),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1055),
.B(n_1064),
.C(n_1032),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1088),
.B(n_1107),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1091),
.B(n_1134),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1165),
.B(n_1167),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1087),
.B(n_1085),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_SL g1240 ( 
.A1(n_1101),
.A2(n_1102),
.B(n_1092),
.C(n_1051),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1161),
.A2(n_1108),
.B(n_1109),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1141),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1126),
.B(n_1097),
.Y(n_1243)
);

INVx6_ASAP7_75t_SL g1244 ( 
.A(n_1105),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_1141),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1100),
.B(n_1150),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1141),
.B(n_1142),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1142),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1126),
.B(n_1103),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1061),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1103),
.B(n_1061),
.Y(n_1251)
);

INVx5_ASAP7_75t_L g1252 ( 
.A(n_1142),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1129),
.B(n_1029),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1081),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1101),
.A2(n_1098),
.B1(n_1058),
.B2(n_1096),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1142),
.Y(n_1256)
);

OAI21xp33_ASAP7_75t_L g1257 ( 
.A1(n_1079),
.A2(n_1096),
.B(n_1098),
.Y(n_1257)
);

AO32x1_ASAP7_75t_L g1258 ( 
.A1(n_1137),
.A2(n_1127),
.A3(n_1067),
.B1(n_1093),
.B2(n_1039),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1150),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_1150),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1058),
.A2(n_1094),
.B1(n_1104),
.B2(n_1075),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1094),
.A2(n_1104),
.B1(n_1075),
.B2(n_1127),
.Y(n_1262)
);

INVx5_ASAP7_75t_L g1263 ( 
.A(n_1093),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1137),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1081),
.B(n_1029),
.Y(n_1265)
);

NAND2xp33_ASAP7_75t_L g1266 ( 
.A(n_1029),
.B(n_1099),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1034),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1029),
.B(n_1047),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1047),
.B(n_1074),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1047),
.B(n_1086),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1047),
.B(n_1060),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_SL g1272 ( 
.A1(n_1052),
.A2(n_1089),
.B(n_1046),
.C(n_1030),
.Y(n_1272)
);

OR2x2_ASAP7_75t_SL g1273 ( 
.A(n_1145),
.B(n_1146),
.Y(n_1273)
);

CKINVDCx6p67_ASAP7_75t_R g1274 ( 
.A(n_1153),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1154),
.B(n_1159),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1162),
.B(n_1110),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1160),
.A2(n_1164),
.B(n_1168),
.C(n_1133),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1112),
.B(n_1158),
.Y(n_1278)
);

BUFx12f_ASAP7_75t_L g1279 ( 
.A(n_1057),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1059),
.B(n_1065),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1024),
.B(n_1120),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1059),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1063),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1160),
.A2(n_1164),
.B(n_921),
.C(n_1012),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1057),
.Y(n_1285)
);

OR2x6_ASAP7_75t_SL g1286 ( 
.A(n_1151),
.B(n_696),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1110),
.B(n_1155),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1035),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1041),
.A2(n_921),
.B1(n_1012),
.B2(n_1010),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1053),
.A2(n_1045),
.B(n_1070),
.Y(n_1290)
);

BUFx4_ASAP7_75t_SL g1291 ( 
.A(n_1069),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1063),
.Y(n_1292)
);

INVx3_ASAP7_75t_SL g1293 ( 
.A(n_1069),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1110),
.B(n_1155),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1057),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1057),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1021),
.A2(n_1050),
.B(n_1112),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1059),
.B(n_1065),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1057),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1024),
.B(n_1120),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1131),
.A2(n_413),
.B1(n_375),
.B2(n_379),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1035),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1026),
.A2(n_1001),
.B(n_999),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1059),
.B(n_1065),
.Y(n_1304)
);

OAI21xp33_ASAP7_75t_L g1305 ( 
.A1(n_1160),
.A2(n_1164),
.B(n_1012),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1035),
.Y(n_1306)
);

AOI21xp33_ASAP7_75t_L g1307 ( 
.A1(n_1054),
.A2(n_1164),
.B(n_1160),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1063),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1026),
.A2(n_1001),
.B(n_999),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1035),
.Y(n_1310)
);

NOR2xp67_ASAP7_75t_L g1311 ( 
.A(n_1038),
.B(n_613),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1026),
.A2(n_1001),
.B(n_999),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1110),
.B(n_1155),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1160),
.B(n_921),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1024),
.B(n_1120),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1041),
.A2(n_748),
.B1(n_921),
.B2(n_676),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1026),
.A2(n_1001),
.B(n_999),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1057),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1048),
.Y(n_1319)
);

BUFx2_ASAP7_75t_SL g1320 ( 
.A(n_1069),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1169),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1171),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1174),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1191),
.A2(n_1301),
.B1(n_1181),
.B2(n_1316),
.Y(n_1324)
);

INVx6_ASAP7_75t_SL g1325 ( 
.A(n_1184),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1191),
.A2(n_1316),
.B1(n_1190),
.B2(n_1180),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1249),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1225),
.A2(n_1190),
.B1(n_1315),
.B2(n_1175),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1201),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1195),
.Y(n_1330)
);

BUFx10_ASAP7_75t_L g1331 ( 
.A(n_1182),
.Y(n_1331)
);

BUFx8_ASAP7_75t_L g1332 ( 
.A(n_1279),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1243),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_1183),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1277),
.A2(n_1284),
.B(n_1314),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1289),
.A2(n_1305),
.B1(n_1307),
.B2(n_1239),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1206),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1213),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1175),
.A2(n_1228),
.B1(n_1224),
.B2(n_1223),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1283),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1292),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1308),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_SL g1343 ( 
.A(n_1319),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1226),
.B(n_1250),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1305),
.A2(n_1307),
.B1(n_1205),
.B2(n_1236),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1173),
.B(n_1281),
.Y(n_1346)
);

INVx4_ASAP7_75t_SL g1347 ( 
.A(n_1265),
.Y(n_1347)
);

AOI222xp33_ASAP7_75t_L g1348 ( 
.A1(n_1300),
.A2(n_1216),
.B1(n_1207),
.B2(n_1212),
.C1(n_1188),
.C2(n_1211),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1205),
.A2(n_1231),
.B1(n_1221),
.B2(n_1216),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1219),
.B(n_1268),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1192),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1215),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1195),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1237),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1188),
.A2(n_1278),
.B1(n_1231),
.B2(n_1229),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1177),
.A2(n_1287),
.B1(n_1294),
.B2(n_1313),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1209),
.A2(n_1269),
.B(n_1241),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1217),
.B(n_1212),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1238),
.Y(n_1359)
);

BUFx10_ASAP7_75t_L g1360 ( 
.A(n_1204),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1214),
.A2(n_1253),
.B(n_1251),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1260),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1179),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1276),
.B(n_1222),
.Y(n_1364)
);

INVxp67_ASAP7_75t_SL g1365 ( 
.A(n_1253),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1264),
.A2(n_1263),
.B1(n_1235),
.B2(n_1266),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1218),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1210),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1286),
.A2(n_1202),
.B1(n_1311),
.B2(n_1263),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1265),
.B(n_1254),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1204),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1270),
.B(n_1271),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1227),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1273),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1260),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1247),
.B(n_1202),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1189),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1189),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1302),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1196),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1196),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1285),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1233),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1291),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1233),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1244),
.A2(n_1220),
.B1(n_1200),
.B2(n_1194),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1288),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1197),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1257),
.A2(n_1235),
.B(n_1230),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1184),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1267),
.Y(n_1391)
);

CKINVDCx6p67_ASAP7_75t_R g1392 ( 
.A(n_1293),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1263),
.A2(n_1208),
.B1(n_1193),
.B2(n_1185),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1285),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1234),
.A2(n_1255),
.B(n_1282),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1242),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1172),
.A2(n_1306),
.B1(n_1310),
.B2(n_1282),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1245),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1320),
.A2(n_1295),
.B1(n_1170),
.B2(n_1299),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1226),
.A2(n_1255),
.B1(n_1193),
.B2(n_1185),
.Y(n_1400)
);

AOI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1303),
.A2(n_1309),
.B(n_1317),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1203),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1186),
.A2(n_1187),
.B1(n_1285),
.B2(n_1296),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1203),
.Y(n_1404)
);

AOI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1312),
.A2(n_1275),
.B(n_1261),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1187),
.B(n_1304),
.Y(n_1406)
);

AO21x1_ASAP7_75t_L g1407 ( 
.A1(n_1262),
.A2(n_1178),
.B(n_1199),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1274),
.Y(n_1408)
);

BUFx8_ASAP7_75t_SL g1409 ( 
.A(n_1296),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1296),
.A2(n_1318),
.B1(n_1304),
.B2(n_1298),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1203),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1290),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1248),
.Y(n_1413)
);

INVx3_ASAP7_75t_SL g1414 ( 
.A(n_1318),
.Y(n_1414)
);

BUFx2_ASAP7_75t_SL g1415 ( 
.A(n_1318),
.Y(n_1415)
);

BUFx8_ASAP7_75t_L g1416 ( 
.A(n_1176),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1272),
.A2(n_1258),
.B(n_1240),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1248),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1248),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1259),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1256),
.B(n_1259),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1280),
.B(n_1298),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1252),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1198),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1246),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1258),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1232),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1232),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1258),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1280),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1176),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1176),
.B(n_1297),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1169),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1267),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1267),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1173),
.A2(n_921),
.B1(n_748),
.B2(n_1041),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1191),
.A2(n_1131),
.B1(n_1301),
.B2(n_1164),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1169),
.Y(n_1438)
);

INVx5_ASAP7_75t_L g1439 ( 
.A(n_1183),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1169),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1173),
.A2(n_921),
.B1(n_748),
.B2(n_1041),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1267),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1179),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1173),
.A2(n_921),
.B1(n_748),
.B2(n_1041),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1169),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1169),
.Y(n_1446)
);

CKINVDCx6p67_ASAP7_75t_R g1447 ( 
.A(n_1293),
.Y(n_1447)
);

BUFx3_ASAP7_75t_L g1448 ( 
.A(n_1195),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1260),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1387),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1363),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1346),
.B(n_1384),
.Y(n_1452)
);

INVx5_ASAP7_75t_SL g1453 ( 
.A(n_1432),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1364),
.B(n_1333),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1443),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1364),
.B(n_1333),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1379),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1350),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1335),
.A2(n_1437),
.B(n_1326),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1360),
.Y(n_1460)
);

AND2x4_ASAP7_75t_SL g1461 ( 
.A(n_1432),
.B(n_1360),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1401),
.A2(n_1412),
.B(n_1426),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1334),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1334),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1372),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1372),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1365),
.Y(n_1467)
);

CKINVDCx11_ASAP7_75t_R g1468 ( 
.A(n_1323),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1426),
.A2(n_1429),
.B(n_1405),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1370),
.B(n_1327),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1374),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1348),
.B(n_1355),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1408),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1327),
.B(n_1321),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1349),
.B(n_1328),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1322),
.B(n_1329),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1337),
.B(n_1338),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1340),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1341),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1342),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1433),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1438),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1440),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1360),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1446),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1391),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1434),
.B(n_1435),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1421),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1408),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1407),
.A2(n_1417),
.B(n_1389),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1347),
.B(n_1442),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1370),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1371),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1357),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1442),
.B(n_1347),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1432),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1368),
.B(n_1429),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1361),
.B(n_1345),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1376),
.B(n_1389),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1432),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1389),
.B(n_1356),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1357),
.B(n_1336),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1436),
.A2(n_1441),
.B(n_1444),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1367),
.B(n_1358),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1324),
.A2(n_1339),
.B1(n_1386),
.B2(n_1351),
.Y(n_1505)
);

AO21x1_ASAP7_75t_SL g1506 ( 
.A1(n_1377),
.A2(n_1385),
.B(n_1378),
.Y(n_1506)
);

BUFx12f_ASAP7_75t_L g1507 ( 
.A(n_1384),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1395),
.B(n_1366),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1417),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1417),
.B(n_1380),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1397),
.B(n_1421),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1354),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1381),
.B(n_1383),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1352),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1359),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1369),
.A2(n_1403),
.B1(n_1410),
.B2(n_1330),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1323),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1390),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1407),
.A2(n_1427),
.B(n_1428),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_SL g1520 ( 
.A(n_1416),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1396),
.B(n_1398),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1362),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1402),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1325),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1404),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1425),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1430),
.B(n_1418),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1411),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1413),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1419),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1420),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1431),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1468),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1499),
.B(n_1501),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1400),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1465),
.B(n_1396),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1465),
.B(n_1398),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1490),
.A2(n_1406),
.B(n_1422),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1472),
.B(n_1508),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1510),
.B(n_1392),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1510),
.B(n_1447),
.Y(n_1541)
);

INVx4_ASAP7_75t_L g1542 ( 
.A(n_1491),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1502),
.B(n_1447),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1466),
.B(n_1424),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1509),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1459),
.A2(n_1448),
.B1(n_1353),
.B2(n_1394),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1480),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1480),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1454),
.B(n_1456),
.Y(n_1549)
);

A2O1A1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1459),
.A2(n_1344),
.B(n_1393),
.C(n_1375),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1454),
.B(n_1373),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1458),
.B(n_1423),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1482),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1482),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1469),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1483),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1497),
.B(n_1414),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_L g1558 ( 
.A(n_1473),
.B(n_1375),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1483),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1472),
.A2(n_1448),
.B1(n_1353),
.B2(n_1449),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1509),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1474),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1469),
.Y(n_1563)
);

AND2x2_ASAP7_75t_SL g1564 ( 
.A(n_1498),
.B(n_1439),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1469),
.B(n_1414),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1462),
.B(n_1449),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1462),
.B(n_1449),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1451),
.Y(n_1568)
);

AND2x4_ASAP7_75t_SL g1569 ( 
.A(n_1463),
.B(n_1331),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_R g1570 ( 
.A(n_1517),
.B(n_1388),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1489),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1508),
.B(n_1362),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1474),
.Y(n_1573)
);

OAI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1503),
.A2(n_1399),
.B1(n_1415),
.B2(n_1362),
.C(n_1388),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1494),
.B(n_1331),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1494),
.B(n_1331),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1494),
.B(n_1394),
.Y(n_1577)
);

OAI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1539),
.A2(n_1475),
.B1(n_1498),
.B2(n_1503),
.C(n_1574),
.Y(n_1578)
);

OR2x6_ASAP7_75t_SL g1579 ( 
.A(n_1544),
.B(n_1511),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1568),
.B(n_1455),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1568),
.B(n_1457),
.Y(n_1581)
);

OAI221xp5_ASAP7_75t_SL g1582 ( 
.A1(n_1539),
.A2(n_1475),
.B1(n_1505),
.B2(n_1511),
.C(n_1516),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1574),
.A2(n_1516),
.B1(n_1452),
.B2(n_1520),
.Y(n_1583)
);

OAI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1550),
.A2(n_1471),
.B1(n_1504),
.B2(n_1515),
.C(n_1512),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1549),
.B(n_1450),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_R g1586 ( 
.A(n_1533),
.B(n_1332),
.Y(n_1586)
);

AOI221x1_ASAP7_75t_SL g1587 ( 
.A1(n_1547),
.A2(n_1521),
.B1(n_1492),
.B2(n_1529),
.C(n_1512),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1549),
.B(n_1478),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1557),
.A2(n_1496),
.B1(n_1500),
.B2(n_1522),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1550),
.A2(n_1497),
.B1(n_1504),
.B2(n_1479),
.C(n_1481),
.Y(n_1590)
);

NAND4xp25_ASAP7_75t_L g1591 ( 
.A(n_1561),
.B(n_1513),
.C(n_1487),
.D(n_1529),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1549),
.B(n_1476),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1533),
.B(n_1507),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1543),
.A2(n_1522),
.B(n_1495),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1534),
.B(n_1495),
.Y(n_1595)
);

OAI221xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1546),
.A2(n_1535),
.B1(n_1544),
.B2(n_1543),
.C(n_1537),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1533),
.B(n_1507),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_R g1598 ( 
.A(n_1572),
.B(n_1332),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1572),
.A2(n_1507),
.B1(n_1382),
.B2(n_1500),
.Y(n_1599)
);

OA211x2_ASAP7_75t_L g1600 ( 
.A1(n_1546),
.A2(n_1520),
.B(n_1506),
.C(n_1332),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1534),
.B(n_1477),
.Y(n_1601)
);

OAI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1560),
.A2(n_1515),
.B1(n_1526),
.B2(n_1518),
.C(n_1531),
.Y(n_1602)
);

OAI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1560),
.A2(n_1526),
.B1(n_1518),
.B2(n_1531),
.C(n_1528),
.Y(n_1603)
);

OAI221xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1535),
.A2(n_1467),
.B1(n_1485),
.B2(n_1525),
.C(n_1530),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1555),
.B(n_1523),
.C(n_1513),
.Y(n_1605)
);

OAI21xp33_ASAP7_75t_L g1606 ( 
.A1(n_1535),
.A2(n_1558),
.B(n_1544),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1540),
.A2(n_1524),
.B(n_1461),
.Y(n_1607)
);

OAI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1565),
.A2(n_1528),
.B1(n_1531),
.B2(n_1532),
.C(n_1467),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1538),
.A2(n_1470),
.B1(n_1514),
.B2(n_1519),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1540),
.B(n_1488),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1541),
.B(n_1488),
.Y(n_1611)
);

NAND3xp33_ASAP7_75t_L g1612 ( 
.A(n_1555),
.B(n_1528),
.C(n_1532),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1536),
.A2(n_1453),
.B1(n_1484),
.B2(n_1460),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_SL g1614 ( 
.A1(n_1564),
.A2(n_1496),
.B1(n_1453),
.B2(n_1461),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1551),
.B(n_1343),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1536),
.Y(n_1616)
);

OAI21xp33_ASAP7_75t_L g1617 ( 
.A1(n_1558),
.A2(n_1527),
.B(n_1493),
.Y(n_1617)
);

OA211x2_ASAP7_75t_L g1618 ( 
.A1(n_1552),
.A2(n_1506),
.B(n_1409),
.C(n_1464),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1557),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1552),
.B(n_1562),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1538),
.A2(n_1514),
.B1(n_1519),
.B2(n_1486),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1562),
.B(n_1519),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1538),
.A2(n_1514),
.B1(n_1519),
.B2(n_1486),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1565),
.B(n_1542),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1622),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1591),
.B(n_1573),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1612),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1619),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1601),
.B(n_1595),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1591),
.B(n_1580),
.Y(n_1630)
);

INVx5_ASAP7_75t_L g1631 ( 
.A(n_1624),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1595),
.B(n_1579),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1612),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1587),
.B(n_1565),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1620),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1579),
.B(n_1545),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1573),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1608),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1592),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1588),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1605),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1605),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1616),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1593),
.B(n_1382),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1606),
.B(n_1547),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1606),
.B(n_1548),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1597),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1585),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1610),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1617),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1584),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1617),
.B(n_1548),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1603),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1611),
.B(n_1571),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1604),
.B(n_1557),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1609),
.B(n_1553),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1621),
.B(n_1542),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1632),
.B(n_1551),
.Y(n_1658)
);

NOR4xp25_ASAP7_75t_L g1659 ( 
.A(n_1641),
.B(n_1578),
.C(n_1582),
.D(n_1596),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1637),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1632),
.B(n_1577),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1634),
.B(n_1536),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1635),
.B(n_1553),
.Y(n_1663)
);

NAND2x1p5_ASAP7_75t_L g1664 ( 
.A(n_1631),
.B(n_1564),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1637),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1537),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1637),
.Y(n_1667)
);

BUFx2_ASAP7_75t_L g1668 ( 
.A(n_1636),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1648),
.Y(n_1669)
);

NAND2xp67_ASAP7_75t_L g1670 ( 
.A(n_1653),
.B(n_1586),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1648),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1641),
.B(n_1537),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1642),
.B(n_1590),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1642),
.B(n_1554),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1635),
.B(n_1554),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1632),
.B(n_1551),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1626),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1629),
.B(n_1575),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1629),
.B(n_1575),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1631),
.B(n_1577),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1643),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1643),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1629),
.B(n_1575),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1636),
.B(n_1576),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1650),
.B(n_1556),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1636),
.B(n_1576),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1626),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1650),
.B(n_1556),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1649),
.B(n_1627),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1631),
.B(n_1576),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1652),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1649),
.B(n_1559),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1652),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1627),
.B(n_1559),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1631),
.B(n_1577),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1640),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1628),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1659),
.B(n_1633),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1677),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1673),
.A2(n_1653),
.B1(n_1651),
.B2(n_1638),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1672),
.B(n_1630),
.Y(n_1701)
);

NOR2xp67_ASAP7_75t_SL g1702 ( 
.A(n_1670),
.B(n_1647),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1672),
.B(n_1630),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1662),
.B(n_1666),
.Y(n_1704)
);

AOI21xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1673),
.A2(n_1630),
.B(n_1655),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1662),
.B(n_1633),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1681),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1689),
.B(n_1666),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1669),
.B(n_1638),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1665),
.B(n_1626),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1677),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1668),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1671),
.B(n_1638),
.Y(n_1713)
);

NOR4xp25_ASAP7_75t_L g1714 ( 
.A(n_1687),
.B(n_1653),
.C(n_1651),
.D(n_1583),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1682),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1696),
.B(n_1651),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1663),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_SL g1718 ( 
.A(n_1664),
.B(n_1647),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1658),
.B(n_1631),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1691),
.B(n_1640),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1661),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1661),
.B(n_1631),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1691),
.B(n_1645),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1668),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1658),
.B(n_1631),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1664),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1675),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1694),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1674),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1674),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1685),
.Y(n_1731)
);

NOR2x2_ASAP7_75t_L g1732 ( 
.A(n_1687),
.B(n_1644),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1661),
.Y(n_1733)
);

CKINVDCx16_ASAP7_75t_R g1734 ( 
.A(n_1676),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1693),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1697),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1693),
.A2(n_1655),
.B(n_1656),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1685),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1660),
.A2(n_1657),
.B1(n_1656),
.B2(n_1655),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1688),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1676),
.B(n_1631),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1732),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1732),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1729),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1730),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1704),
.B(n_1665),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1731),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1712),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1740),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1740),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1738),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1724),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1734),
.B(n_1667),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1721),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1707),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1733),
.Y(n_1756)
);

NOR3xp33_ASAP7_75t_L g1757 ( 
.A(n_1698),
.B(n_1697),
.C(n_1667),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1699),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1722),
.B(n_1684),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1705),
.B(n_1688),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1728),
.B(n_1647),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1722),
.B(n_1686),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1706),
.B(n_1692),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1719),
.B(n_1686),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1709),
.B(n_1628),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1708),
.B(n_1645),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1715),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1716),
.Y(n_1769)
);

INVx4_ASAP7_75t_L g1770 ( 
.A(n_1726),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1718),
.B(n_1647),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1719),
.B(n_1664),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1735),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1708),
.B(n_1646),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1735),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_1713),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1701),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1748),
.B(n_1714),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1773),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1773),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1761),
.A2(n_1737),
.B(n_1700),
.Y(n_1781)
);

AOI31xp33_ASAP7_75t_L g1782 ( 
.A1(n_1742),
.A2(n_1718),
.A3(n_1736),
.B(n_1703),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1775),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1743),
.A2(n_1739),
.B1(n_1741),
.B2(n_1726),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1777),
.A2(n_1741),
.B1(n_1726),
.B2(n_1725),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1756),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1752),
.A2(n_1710),
.B1(n_1723),
.B2(n_1657),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1746),
.B(n_1710),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1757),
.A2(n_1657),
.B1(n_1720),
.B2(n_1647),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1753),
.B(n_1754),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1769),
.B(n_1717),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1776),
.A2(n_1699),
.B1(n_1711),
.B2(n_1702),
.Y(n_1792)
);

AO211x2_ASAP7_75t_L g1793 ( 
.A1(n_1744),
.A2(n_1670),
.B(n_1727),
.C(n_1646),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1756),
.A2(n_1741),
.B(n_1725),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1753),
.B(n_1647),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1746),
.B(n_1711),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1775),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1771),
.A2(n_1768),
.B(n_1755),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1765),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1755),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1770),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1768),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1744),
.B(n_1745),
.Y(n_1803)
);

NAND2x1p5_ASAP7_75t_L g1804 ( 
.A(n_1786),
.B(n_1770),
.Y(n_1804)
);

NOR2x1_ASAP7_75t_L g1805 ( 
.A(n_1782),
.B(n_1770),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1778),
.B(n_1647),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1781),
.B(n_1745),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1790),
.B(n_1747),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1782),
.A2(n_1766),
.B1(n_1771),
.B2(n_1767),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1801),
.Y(n_1810)
);

NAND2xp33_ASAP7_75t_L g1811 ( 
.A(n_1788),
.B(n_1570),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1799),
.B(n_1758),
.Y(n_1812)
);

NAND2x1_ASAP7_75t_L g1813 ( 
.A(n_1795),
.B(n_1770),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1796),
.B(n_1747),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1795),
.B(n_1758),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1800),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1802),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1779),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1780),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1783),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_R g1821 ( 
.A(n_1797),
.B(n_1751),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_SL g1822 ( 
.A1(n_1798),
.A2(n_1794),
.B(n_1789),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1803),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1804),
.Y(n_1824)
);

AOI211xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1809),
.A2(n_1822),
.B(n_1807),
.C(n_1810),
.Y(n_1825)
);

NOR3xp33_ASAP7_75t_L g1826 ( 
.A(n_1809),
.B(n_1784),
.C(n_1787),
.Y(n_1826)
);

A2O1A1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1822),
.A2(n_1806),
.B(n_1805),
.C(n_1793),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1814),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1808),
.A2(n_1789),
.B1(n_1787),
.B2(n_1792),
.Y(n_1829)
);

NOR2x1_ASAP7_75t_L g1830 ( 
.A(n_1820),
.B(n_1798),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1811),
.A2(n_1791),
.B(n_1785),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1815),
.A2(n_1749),
.B1(n_1750),
.B2(n_1759),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1816),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_SL g1834 ( 
.A(n_1821),
.B(n_1762),
.C(n_1750),
.Y(n_1834)
);

NAND4xp25_ASAP7_75t_L g1835 ( 
.A(n_1812),
.B(n_1751),
.C(n_1772),
.D(n_1763),
.Y(n_1835)
);

NOR2x1_ASAP7_75t_L g1836 ( 
.A(n_1830),
.B(n_1817),
.Y(n_1836)
);

NAND4xp25_ASAP7_75t_L g1837 ( 
.A(n_1825),
.B(n_1823),
.C(n_1812),
.D(n_1818),
.Y(n_1837)
);

NOR4xp25_ASAP7_75t_L g1838 ( 
.A(n_1827),
.B(n_1819),
.C(n_1749),
.D(n_1750),
.Y(n_1838)
);

NAND4xp75_ASAP7_75t_L g1839 ( 
.A(n_1831),
.B(n_1828),
.C(n_1824),
.D(n_1832),
.Y(n_1839)
);

NOR4xp75_ASAP7_75t_L g1840 ( 
.A(n_1829),
.B(n_1813),
.C(n_1804),
.D(n_1763),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1826),
.A2(n_1749),
.B1(n_1759),
.B2(n_1772),
.Y(n_1841)
);

NAND4xp25_ASAP7_75t_L g1842 ( 
.A(n_1835),
.B(n_1760),
.C(n_1765),
.D(n_1764),
.Y(n_1842)
);

NOR3xp33_ASAP7_75t_L g1843 ( 
.A(n_1834),
.B(n_1759),
.C(n_1767),
.Y(n_1843)
);

NOR3xp33_ASAP7_75t_L g1844 ( 
.A(n_1833),
.B(n_1774),
.C(n_1764),
.Y(n_1844)
);

NAND4xp75_ASAP7_75t_L g1845 ( 
.A(n_1830),
.B(n_1600),
.C(n_1760),
.D(n_1409),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1830),
.Y(n_1846)
);

NOR4xp25_ASAP7_75t_SL g1847 ( 
.A(n_1846),
.B(n_1607),
.C(n_1570),
.D(n_1594),
.Y(n_1847)
);

OAI211xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1836),
.A2(n_1774),
.B(n_1615),
.C(n_1607),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1839),
.B(n_1678),
.Y(n_1849)
);

NOR4xp25_ASAP7_75t_L g1850 ( 
.A(n_1837),
.B(n_1625),
.C(n_1679),
.D(n_1683),
.Y(n_1850)
);

NAND4xp25_ASAP7_75t_L g1851 ( 
.A(n_1841),
.B(n_1618),
.C(n_1600),
.D(n_1695),
.Y(n_1851)
);

NOR3xp33_ASAP7_75t_SL g1852 ( 
.A(n_1842),
.B(n_1599),
.C(n_1644),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1843),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1849),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1853),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1848),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1852),
.Y(n_1857)
);

NOR2x1_ASAP7_75t_L g1858 ( 
.A(n_1851),
.B(n_1845),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1850),
.A2(n_1838),
.B1(n_1844),
.B2(n_1840),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1847),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1849),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1853),
.A2(n_1657),
.B1(n_1599),
.B2(n_1625),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1854),
.Y(n_1863)
);

NAND5xp2_ASAP7_75t_L g1864 ( 
.A(n_1860),
.B(n_1690),
.C(n_1614),
.D(n_1602),
.E(n_1618),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1861),
.Y(n_1865)
);

NAND2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1855),
.B(n_1680),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1856),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1859),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1863),
.Y(n_1869)
);

NOR3xp33_ASAP7_75t_L g1870 ( 
.A(n_1868),
.B(n_1857),
.C(n_1858),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1866),
.B(n_1862),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1871),
.A2(n_1867),
.B1(n_1865),
.B2(n_1864),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1872),
.A2(n_1870),
.B1(n_1869),
.B2(n_1864),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1873),
.A2(n_1695),
.B1(n_1680),
.B2(n_1657),
.Y(n_1874)
);

OA21x2_ASAP7_75t_L g1875 ( 
.A1(n_1873),
.A2(n_1679),
.B(n_1678),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1875),
.A2(n_1639),
.B1(n_1683),
.B2(n_1680),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1874),
.B(n_1563),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1598),
.B1(n_1695),
.B2(n_1563),
.C(n_1623),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1876),
.A2(n_1639),
.B(n_1569),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1878),
.A2(n_1567),
.B(n_1566),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1880),
.A2(n_1879),
.B1(n_1416),
.B2(n_1569),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_1416),
.B1(n_1569),
.B2(n_1654),
.Y(n_1882)
);

AOI211xp5_ASAP7_75t_L g1883 ( 
.A1(n_1882),
.A2(n_1613),
.B(n_1690),
.C(n_1589),
.Y(n_1883)
);


endmodule