module real_aes_14313_n_4 (n_0, n_3, n_2, n_1, n_4);
input n_0;
input n_3;
input n_2;
input n_1;
output n_4;
wire n_16;
wire n_13;
wire n_5;
wire n_15;
wire n_7;
wire n_9;
wire n_12;
wire n_6;
wire n_8;
wire n_14;
wire n_10;
wire n_11;
INVx1_ASAP7_75t_L g8 ( .A(n_0), .Y(n_8) );
INVx1_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
AOI21xp5_ASAP7_75t_L g11 ( .A1(n_1), .A2(n_12), .B(n_13), .Y(n_11) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
NOR3xp33_ASAP7_75t_L g15 ( .A(n_2), .B(n_7), .C(n_16), .Y(n_15) );
INVx1_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_3), .B(n_10), .Y(n_13) );
AOI21xp33_ASAP7_75t_L g4 ( .A1(n_5), .A2(n_14), .B(n_15), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_6), .Y(n_5) );
AOI21xp33_ASAP7_75t_L g6 ( .A1(n_7), .A2(n_9), .B(n_11), .Y(n_6) );
BUFx2_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
HB1xp67_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
INVx1_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
endmodule