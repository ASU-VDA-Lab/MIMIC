module fake_jpeg_19398_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_18),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_71),
.Y(n_79)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_73),
.B(n_50),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_68),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_57),
.B1(n_66),
.B2(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_80),
.B1(n_47),
.B2(n_61),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_48),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_53),
.B1(n_66),
.B2(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_83),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_63),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g85 ( 
.A1(n_79),
.A2(n_73),
.B(n_70),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_87),
.B1(n_97),
.B2(n_0),
.Y(n_104)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_91),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_94),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_64),
.B(n_49),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_50),
.C(n_54),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_60),
.B1(n_65),
.B2(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_103),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_111),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_105),
.B1(n_1),
.B2(n_3),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_20),
.B1(n_41),
.B2(n_40),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_56),
.B1(n_17),
.B2(n_23),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_39),
.B(n_15),
.C(n_27),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_13),
.B1(n_38),
.B2(n_37),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_117),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_116),
.B1(n_119),
.B2(n_104),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_102),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_99),
.C(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_24),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_118),
.B(n_116),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_122),
.C(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_124),
.C(n_110),
.Y(n_127)
);

AOI221xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_113),
.B1(n_119),
.B2(n_106),
.C(n_8),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_107),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_10),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_9),
.A3(n_34),
.B1(n_32),
.B2(n_31),
.C1(n_35),
.C2(n_8),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_4),
.Y(n_133)
);


endmodule