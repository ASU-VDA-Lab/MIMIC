module fake_ariane_3212_n_1967 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1967);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1967;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_59),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_165),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_72),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_81),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_44),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_98),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_83),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_23),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_174),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_25),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_130),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_89),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_187),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_125),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_109),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_175),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_50),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_74),
.Y(n_233)
);

BUFx2_ASAP7_75t_SL g234 ( 
.A(n_39),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_41),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_124),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_155),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_60),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_135),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_17),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_34),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_136),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_53),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_205),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_70),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_1),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_110),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_21),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_8),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_4),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_172),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_46),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_17),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_149),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_182),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_111),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_105),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_169),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_201),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_102),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_20),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_34),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_67),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_71),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_208),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_100),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_53),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_13),
.Y(n_277)
);

HB1xp67_ASAP7_75t_SL g278 ( 
.A(n_21),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_47),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_63),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_82),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_114),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_86),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_115),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_20),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_179),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_84),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_22),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_140),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_3),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_184),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_153),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_141),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_13),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_129),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_103),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_163),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_121),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_2),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_131),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_151),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_200),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_133),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_95),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_69),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_73),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_154),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_116),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_138),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_202),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_66),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_164),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_87),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_29),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_57),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_26),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_158),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_112),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_168),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_40),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_108),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_204),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_10),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_159),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_118),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_123),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_11),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_171),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_167),
.Y(n_330)
);

BUFx2_ASAP7_75t_SL g331 ( 
.A(n_52),
.Y(n_331)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_41),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_26),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_176),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_85),
.Y(n_335)
);

BUFx10_ASAP7_75t_L g336 ( 
.A(n_36),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_113),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_181),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_35),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_57),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_94),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_148),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_139),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_91),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_146),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_54),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_189),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_196),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_16),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_75),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_126),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_142),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_54),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_30),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_170),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_24),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_99),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_147),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_104),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_157),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_28),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_119),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_24),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_60),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_177),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_23),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_106),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_185),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_162),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_90),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_14),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_127),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_51),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_22),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_43),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_27),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_194),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_59),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_14),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_203),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_6),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_166),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_128),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_29),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_186),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_10),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_6),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_132),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_37),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_192),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_19),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_55),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_96),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_161),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_63),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_51),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_78),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_31),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_92),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_8),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_30),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_56),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_45),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g404 ( 
.A(n_27),
.Y(n_404)
);

BUFx10_ASAP7_75t_L g405 ( 
.A(n_47),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_80),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_9),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_33),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_16),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_25),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_101),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_197),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_137),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_268),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_268),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_278),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_266),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_242),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_270),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_386),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_395),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_351),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_404),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_404),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_404),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_404),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_295),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_345),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_213),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_404),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_232),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_245),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_265),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_267),
.Y(n_438)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_272),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_370),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_383),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_332),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_332),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_332),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_211),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_211),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_275),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_336),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_234),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_281),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_336),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_212),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_217),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_315),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_316),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_336),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_250),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_317),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_250),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_339),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_340),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_346),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_248),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_354),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_354),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_356),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_354),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_345),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_405),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_363),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_212),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_284),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_384),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_331),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_391),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_405),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_405),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_218),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_250),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_403),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_218),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_250),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_345),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_409),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_289),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_235),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_289),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_400),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_217),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_220),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_408),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_222),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_408),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_235),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_222),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_250),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_318),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_353),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_252),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_253),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_353),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_253),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_253),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_253),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_255),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_253),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_224),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_210),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_284),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_214),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_338),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_256),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_224),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_215),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_277),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_216),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_459),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_503),
.Y(n_519)
);

INVx5_ASAP7_75t_L g520 ( 
.A(n_429),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_504),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_459),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_490),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_429),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_424),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_425),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_219),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_419),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_426),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_429),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_429),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_512),
.B(n_422),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_468),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_227),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_468),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_419),
.A2(n_243),
.B1(n_387),
.B2(n_240),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_468),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_452),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_509),
.B(n_338),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_468),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_479),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_427),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_430),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_457),
.B(n_236),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_493),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_511),
.B(n_294),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_432),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_418),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_433),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_439),
.B(n_240),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g553 ( 
.A(n_443),
.B(n_221),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_434),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_482),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_421),
.A2(n_387),
.B1(n_389),
.B2(n_243),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_420),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_505),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_493),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_483),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_501),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_421),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_423),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_501),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_452),
.B(n_280),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_498),
.B(n_294),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_498),
.B(n_471),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_483),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_515),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_517),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_445),
.Y(n_571)
);

AND2x6_ASAP7_75t_L g572 ( 
.A(n_483),
.B(n_221),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_471),
.B(n_478),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_483),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_485),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_487),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_488),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_489),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_492),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_496),
.A2(n_514),
.B1(n_508),
.B2(n_444),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_494),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_478),
.B(n_237),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_435),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_436),
.A2(n_241),
.B(n_238),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_437),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_438),
.Y(n_586)
);

AND2x2_ASAP7_75t_SL g587 ( 
.A(n_446),
.B(n_229),
.Y(n_587)
);

INVxp67_ASAP7_75t_SL g588 ( 
.A(n_449),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_447),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_481),
.B(n_273),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_454),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_455),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_458),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_440),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g596 ( 
.A(n_481),
.B(n_246),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_491),
.B(n_276),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_279),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_460),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_441),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_555),
.B(n_558),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_555),
.B(n_431),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_528),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_583),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_528),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_524),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_526),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_526),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_587),
.A2(n_431),
.B1(n_453),
.B2(n_496),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_527),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_463),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_558),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_583),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_583),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_531),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_531),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_544),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_540),
.B(n_417),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_583),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_545),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_545),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_535),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_549),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_583),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_551),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_596),
.B(n_500),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_554),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_566),
.B(n_598),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_534),
.B(n_506),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_587),
.B(n_513),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_553),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_535),
.Y(n_636)
);

AND2x2_ASAP7_75t_SL g637 ( 
.A(n_587),
.B(n_229),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_554),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_561),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_550),
.Y(n_640)
);

INVx6_ASAP7_75t_L g641 ( 
.A(n_583),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_567),
.A2(n_508),
.B1(n_514),
.B2(n_410),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_519),
.Y(n_645)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_584),
.B(n_591),
.C(n_589),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_564),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_564),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_518),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_519),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_521),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_521),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_589),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_548),
.A2(n_428),
.B1(n_499),
.B2(n_495),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_522),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_540),
.B(n_516),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_589),
.Y(n_657)
);

AOI21x1_ASAP7_75t_L g658 ( 
.A1(n_584),
.A2(n_260),
.B(n_251),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_557),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_518),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_522),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_589),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_518),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_518),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_569),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_553),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_595),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_600),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_569),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_546),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_589),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_570),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_R g674 ( 
.A(n_563),
.B(n_428),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_591),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_523),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_553),
.B(n_474),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_552),
.B(n_220),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_552),
.B(n_414),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_535),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_582),
.B(n_223),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_588),
.B(n_548),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_548),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_523),
.Y(n_684)
);

OAI21xp33_ASAP7_75t_SL g685 ( 
.A1(n_570),
.A2(n_486),
.B(n_462),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_591),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_523),
.Y(n_687)
);

BUFx6f_ASAP7_75t_SL g688 ( 
.A(n_548),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_590),
.B(n_597),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_547),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_591),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_541),
.B(n_223),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_541),
.B(n_225),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_591),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_L g695 ( 
.A(n_591),
.B(n_225),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_592),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_523),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_529),
.B(n_541),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_543),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_538),
.B(n_415),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_541),
.B(n_497),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_543),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_543),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_556),
.B(n_416),
.Y(n_704)
);

BUFx4f_ASAP7_75t_L g705 ( 
.A(n_584),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_592),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_565),
.B(n_502),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_535),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_592),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_592),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_592),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_576),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_543),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_585),
.B(n_461),
.Y(n_714)
);

INVxp33_ASAP7_75t_L g715 ( 
.A(n_547),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_SL g716 ( 
.A(n_585),
.B(n_442),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_525),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_576),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_535),
.Y(n_719)
);

AO21x2_ASAP7_75t_L g720 ( 
.A1(n_536),
.A2(n_287),
.B(n_282),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_593),
.A2(n_392),
.B1(n_396),
.B2(n_389),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_576),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_577),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_593),
.A2(n_396),
.B1(n_398),
.B2(n_392),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_577),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_577),
.Y(n_726)
);

AOI21x1_ASAP7_75t_L g727 ( 
.A1(n_584),
.A2(n_260),
.B(n_251),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_525),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_525),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_530),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_586),
.B(n_466),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_532),
.Y(n_732)
);

CKINVDCx6p67_ASAP7_75t_R g733 ( 
.A(n_562),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_532),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_559),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_578),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_578),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_532),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_586),
.B(n_470),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_586),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_578),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_533),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_580),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_572),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_594),
.B(n_290),
.C(n_288),
.Y(n_745)
);

BUFx10_ASAP7_75t_L g746 ( 
.A(n_572),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_533),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_632),
.B(n_599),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_689),
.B(n_599),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_603),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_L g751 ( 
.A(n_607),
.B(n_226),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_671),
.B(n_599),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_637),
.A2(n_401),
.B1(n_402),
.B2(n_398),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_637),
.A2(n_581),
.B1(n_230),
.B2(n_231),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_644),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_637),
.B(n_581),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_611),
.B(n_581),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_633),
.B(n_581),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_730),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_635),
.B(n_579),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_685),
.A2(n_575),
.B(n_480),
.C(n_484),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_744),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_683),
.B(n_228),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_683),
.B(n_228),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_746),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_685),
.A2(n_575),
.B(n_473),
.C(n_475),
.Y(n_766)
);

BUFx8_ASAP7_75t_L g767 ( 
.A(n_659),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_634),
.B(n_579),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_635),
.B(n_579),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_603),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_665),
.A2(n_401),
.B1(n_402),
.B2(n_407),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_666),
.B(n_286),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_666),
.B(n_257),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_677),
.B(n_291),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_705),
.A2(n_572),
.B1(n_465),
.B2(n_442),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_698),
.B(n_301),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_665),
.A2(n_407),
.B1(n_300),
.B2(n_349),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_740),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_683),
.B(n_230),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_613),
.B(n_313),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_607),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_608),
.B(n_231),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_683),
.B(n_233),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_705),
.A2(n_572),
.B1(n_467),
.B2(n_465),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_618),
.A2(n_539),
.B(n_537),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_619),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_619),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_705),
.A2(n_572),
.B1(n_469),
.B2(n_467),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_605),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_623),
.B(n_233),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_605),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_610),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_613),
.B(n_239),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_707),
.A2(n_406),
.B1(n_385),
.B2(n_388),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_669),
.B(n_239),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_669),
.B(n_244),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_740),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_673),
.A2(n_379),
.B1(n_381),
.B2(n_361),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_623),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_625),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_610),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_659),
.Y(n_803)
);

INVx3_ASAP7_75t_R g804 ( 
.A(n_667),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_625),
.A2(n_539),
.B(n_537),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_612),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_673),
.B(n_682),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_629),
.B(n_244),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_629),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_667),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_612),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_631),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_640),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_731),
.B(n_319),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_631),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_731),
.B(n_320),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_731),
.B(n_320),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_638),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_601),
.B(n_388),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_638),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_688),
.A2(n_390),
.B1(n_394),
.B2(n_397),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_679),
.B(n_390),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_SL g823 ( 
.A(n_640),
.B(n_630),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_609),
.B(n_324),
.C(n_321),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_616),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_679),
.B(n_394),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_615),
.B(n_397),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_645),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_615),
.B(n_399),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_602),
.B(n_399),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_615),
.B(n_710),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_701),
.B(n_406),
.Y(n_832)
);

NOR2x1p5_ASAP7_75t_L g833 ( 
.A(n_733),
.B(n_328),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_668),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_668),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_615),
.B(n_412),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_616),
.A2(n_622),
.B1(n_627),
.B2(n_617),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_617),
.A2(n_574),
.B(n_539),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_678),
.B(n_333),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_645),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_739),
.B(n_412),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_656),
.B(n_366),
.C(n_364),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_620),
.A2(n_371),
.B1(n_373),
.B2(n_374),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_622),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_615),
.B(n_296),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_744),
.B(n_297),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_620),
.B(n_559),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_627),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_628),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_628),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_712),
.B(n_375),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_710),
.B(n_298),
.Y(n_852)
);

NOR2x1_ASAP7_75t_L g853 ( 
.A(n_620),
.B(n_444),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_710),
.B(n_303),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_712),
.B(n_376),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_710),
.B(n_650),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_735),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_718),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_722),
.B(n_378),
.Y(n_859)
);

AO221x1_ASAP7_75t_L g860 ( 
.A1(n_721),
.A2(n_456),
.B1(n_469),
.B2(n_476),
.C(n_448),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_620),
.A2(n_306),
.B1(n_350),
.B2(n_362),
.Y(n_861)
);

INVx8_ASAP7_75t_L g862 ( 
.A(n_688),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_722),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_723),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_724),
.B(n_448),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_681),
.B(n_692),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_730),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_700),
.B(n_704),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_723),
.B(n_247),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_725),
.B(n_726),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_725),
.B(n_249),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_650),
.A2(n_572),
.B1(n_477),
.B2(n_451),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_724),
.B(n_451),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_726),
.Y(n_874)
);

BUFx6f_ASAP7_75t_SL g875 ( 
.A(n_700),
.Y(n_875)
);

OAI22xp33_ASAP7_75t_L g876 ( 
.A1(n_642),
.A2(n_456),
.B1(n_464),
.B2(n_477),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_736),
.B(n_254),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_649),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_649),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_710),
.B(n_310),
.Y(n_880)
);

NOR2xp67_ASAP7_75t_L g881 ( 
.A(n_745),
.B(n_568),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_651),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_736),
.B(n_258),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_651),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_652),
.A2(n_337),
.B1(n_358),
.B2(n_343),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_604),
.B(n_334),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_604),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_690),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_674),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_642),
.A2(n_393),
.B(n_341),
.C(n_365),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_693),
.B(n_464),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_641),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_714),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_737),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_737),
.B(n_259),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_604),
.B(n_372),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_741),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_741),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_716),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_655),
.Y(n_900)
);

AND2x6_ASAP7_75t_L g901 ( 
.A(n_662),
.B(n_309),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_655),
.B(n_261),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_606),
.B(n_0),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_715),
.B(n_0),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_688),
.A2(n_380),
.B1(n_413),
.B2(n_327),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_614),
.B(n_309),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_660),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_661),
.B(n_262),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_661),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_781),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_R g911 ( 
.A(n_767),
.B(n_743),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_748),
.B(n_639),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_748),
.B(n_639),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_749),
.B(n_643),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_755),
.B(n_654),
.Y(n_915)
);

NAND2x1p5_ASAP7_75t_L g916 ( 
.A(n_762),
.B(n_744),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_868),
.B(n_803),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_783),
.B(n_643),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_857),
.B(n_759),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_R g920 ( 
.A(n_767),
.B(n_662),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_868),
.A2(n_700),
.B1(n_704),
.B2(n_695),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_888),
.B(n_700),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_787),
.B(n_647),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_788),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_800),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_801),
.B(n_647),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_803),
.B(n_700),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_862),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_862),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_809),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_812),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_815),
.B(n_648),
.Y(n_932)
);

AND2x6_ASAP7_75t_SL g933 ( 
.A(n_865),
.B(n_704),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_835),
.Y(n_934)
);

BUFx8_ASAP7_75t_L g935 ( 
.A(n_875),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_818),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_899),
.B(n_704),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_853),
.B(n_614),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_893),
.B(n_720),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_867),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_756),
.A2(n_646),
.B(n_658),
.Y(n_941)
);

AND2x6_ASAP7_75t_SL g942 ( 
.A(n_873),
.B(n_670),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_889),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_820),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_828),
.Y(n_945)
);

AND3x2_ASAP7_75t_SL g946 ( 
.A(n_876),
.B(n_326),
.C(n_648),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_810),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_834),
.B(n_621),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_772),
.A2(n_641),
.B1(n_694),
.B2(n_691),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_847),
.Y(n_950)
);

INVx5_ASAP7_75t_L g951 ( 
.A(n_862),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_840),
.B(n_720),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_876),
.B(n_621),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_804),
.B(n_621),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_882),
.Y(n_955)
);

NAND3xp33_ASAP7_75t_L g956 ( 
.A(n_795),
.B(n_772),
.C(n_753),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_884),
.B(n_720),
.Y(n_957)
);

BUFx4f_ASAP7_75t_L g958 ( 
.A(n_904),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_903),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_891),
.B(n_626),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_892),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_900),
.B(n_663),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_861),
.A2(n_641),
.B1(n_694),
.B2(n_626),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_SL g964 ( 
.A(n_842),
.B(n_745),
.C(n_264),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_909),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_768),
.B(n_663),
.Y(n_966)
);

BUFx4f_ASAP7_75t_L g967 ( 
.A(n_901),
.Y(n_967)
);

AND2x4_ASAP7_75t_SL g968 ( 
.A(n_872),
.B(n_746),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_807),
.B(n_626),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_858),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_774),
.A2(n_641),
.B1(n_675),
.B2(n_657),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_762),
.B(n_653),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_754),
.A2(n_646),
.B1(n_675),
.B2(n_691),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_776),
.B(n_664),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_773),
.B(n_676),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_892),
.Y(n_976)
);

NOR3xp33_ASAP7_75t_SL g977 ( 
.A(n_771),
.B(n_269),
.C(n_263),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_825),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_891),
.B(n_653),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_825),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_858),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_758),
.B(n_653),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_833),
.B(n_657),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_780),
.B(n_676),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_844),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_824),
.A2(n_702),
.B1(n_703),
.B2(n_697),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_887),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_814),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_846),
.B(n_657),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_822),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_768),
.B(n_684),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_826),
.B(n_872),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_843),
.B(n_777),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_819),
.B(n_684),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_866),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_863),
.B(n_687),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_778),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_863),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_864),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_R g1000 ( 
.A(n_751),
.B(n_670),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_802),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_864),
.B(n_687),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_874),
.B(n_697),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_874),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_894),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_757),
.B(n_794),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_775),
.A2(n_713),
.B1(n_703),
.B2(n_702),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_811),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_778),
.B(n_761),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_887),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_849),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_894),
.Y(n_1012)
);

AOI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_774),
.A2(n_691),
.B1(n_675),
.B2(n_694),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_890),
.B(n_699),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_SL g1015 ( 
.A1(n_875),
.A2(n_326),
.B1(n_746),
.B2(n_355),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_897),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_SL g1017 ( 
.A(n_890),
.B(n_302),
.C(n_271),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_SL g1018 ( 
.A(n_791),
.B(n_304),
.C(n_274),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_799),
.B(n_699),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_866),
.B(n_672),
.Y(n_1020)
);

INVx5_ASAP7_75t_L g1021 ( 
.A(n_765),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_898),
.B(n_713),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_898),
.B(n_672),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_830),
.B(n_686),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_793),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_793),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_806),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_806),
.B(n_686),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_878),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_SL g1030 ( 
.A1(n_775),
.A2(n_293),
.B1(n_283),
.B2(n_285),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_SL g1031 ( 
.A(n_791),
.B(n_305),
.C(n_292),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_848),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_821),
.B(n_696),
.Y(n_1033)
);

AND2x6_ASAP7_75t_L g1034 ( 
.A(n_765),
.B(n_696),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_848),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_850),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_839),
.B(n_706),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_850),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_816),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_846),
.B(n_746),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_879),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_761),
.B(n_706),
.Y(n_1042)
);

NAND2x1p5_ASAP7_75t_L g1043 ( 
.A(n_765),
.B(n_709),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_798),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_765),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_785),
.A2(n_711),
.B1(n_709),
.B2(n_742),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_907),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_796),
.Y(n_1048)
);

AND2x2_ASAP7_75t_SL g1049 ( 
.A(n_785),
.B(n_711),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_782),
.A2(n_299),
.B1(n_307),
.B2(n_308),
.Y(n_1050)
);

OR2x6_ASAP7_75t_L g1051 ( 
.A(n_766),
.B(n_717),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_839),
.B(n_717),
.Y(n_1052)
);

AO22x1_ASAP7_75t_L g1053 ( 
.A1(n_901),
.A2(n_572),
.B1(n_311),
.B2(n_368),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_808),
.A2(n_312),
.B1(n_314),
.B2(n_322),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_752),
.B(n_728),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_837),
.B(n_728),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_763),
.A2(n_323),
.B1(n_325),
.B2(n_329),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_905),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_837),
.B(n_729),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_870),
.B(n_729),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_750),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_770),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_885),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_R g1064 ( 
.A(n_856),
.B(n_624),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_760),
.B(n_732),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_770),
.Y(n_1066)
);

NAND2x2_ASAP7_75t_L g1067 ( 
.A(n_823),
.B(n_1),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_790),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_860),
.B(n_747),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_789),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_763),
.A2(n_680),
.B(n_624),
.C(n_636),
.Y(n_1071)
);

AND2x6_ASAP7_75t_SL g1072 ( 
.A(n_797),
.B(n_3),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_764),
.B(n_624),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_789),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_790),
.Y(n_1075)
);

BUFx4f_ASAP7_75t_L g1076 ( 
.A(n_901),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_792),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_851),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_817),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_769),
.B(n_732),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_792),
.B(n_734),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_855),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_859),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_831),
.A2(n_636),
.B(n_719),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_832),
.B(n_738),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_764),
.A2(n_572),
.B1(n_719),
.B2(n_708),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_841),
.B(n_636),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_950),
.B(n_902),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_917),
.B(n_779),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_929),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_912),
.B(n_908),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_912),
.B(n_779),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_934),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_917),
.B(n_784),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_913),
.A2(n_831),
.B(n_784),
.Y(n_1095)
);

AND3x1_ASAP7_75t_SL g1096 ( 
.A(n_946),
.B(n_4),
.C(n_5),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_913),
.B(n_901),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_929),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_911),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_929),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_956),
.B(n_827),
.C(n_829),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1063),
.B(n_869),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_993),
.A2(n_995),
.B1(n_1074),
.B2(n_1070),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_914),
.A2(n_829),
.B(n_827),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_914),
.B(n_901),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1082),
.B(n_871),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_960),
.B(n_877),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1083),
.B(n_883),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1020),
.B(n_895),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_953),
.A2(n_836),
.B1(n_896),
.B2(n_886),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_SL g1111 ( 
.A1(n_1006),
.A2(n_982),
.B(n_1087),
.C(n_962),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_990),
.B(n_886),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_920),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_966),
.A2(n_836),
.B(n_896),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_928),
.B(n_929),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_941),
.A2(n_727),
.B(n_658),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_966),
.A2(n_786),
.B(n_805),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_991),
.A2(n_906),
.B(n_838),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1078),
.A2(n_906),
.B(n_845),
.C(n_880),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_988),
.B(n_845),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_951),
.B(n_852),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_947),
.A2(n_880),
.B(n_854),
.C(n_852),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1087),
.A2(n_854),
.B(n_680),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_994),
.A2(n_680),
.B(n_719),
.Y(n_1124)
);

O2A1O1Ixp5_ASAP7_75t_L g1125 ( 
.A1(n_979),
.A2(n_708),
.B(n_727),
.C(n_574),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_940),
.B(n_708),
.Y(n_1126)
);

AOI22x1_ASAP7_75t_SL g1127 ( 
.A1(n_1058),
.A2(n_330),
.B1(n_335),
.B2(n_342),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_992),
.B(n_881),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_921),
.A2(n_360),
.B1(n_347),
.B2(n_348),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_970),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_910),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_981),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_919),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_958),
.B(n_344),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_1072),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_935),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_935),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_927),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_958),
.B(n_352),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_998),
.Y(n_1140)
);

AOI33xp33_ASAP7_75t_L g1141 ( 
.A1(n_924),
.A2(n_574),
.A3(n_537),
.B1(n_9),
.B2(n_11),
.B3(n_12),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_967),
.Y(n_1142)
);

AOI222xp33_ASAP7_75t_L g1143 ( 
.A1(n_915),
.A2(n_369),
.B1(n_357),
.B2(n_359),
.C1(n_377),
.C2(n_367),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_922),
.B(n_5),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1009),
.B(n_568),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_925),
.A2(n_411),
.B1(n_382),
.B2(n_345),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_927),
.B(n_937),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1039),
.A2(n_7),
.B(n_12),
.C(n_15),
.Y(n_1148)
);

NOR2xp67_ASAP7_75t_L g1149 ( 
.A(n_951),
.B(n_68),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_950),
.B(n_15),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_SL g1151 ( 
.A(n_977),
.B(n_18),
.C(n_19),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1016),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1048),
.B(n_18),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_937),
.B(n_28),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_943),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_930),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1009),
.B(n_31),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_931),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1030),
.A2(n_968),
.B1(n_959),
.B2(n_1011),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_999),
.B(n_32),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_951),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1004),
.B(n_32),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1005),
.B(n_33),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1060),
.A2(n_923),
.B(n_918),
.Y(n_1164)
);

NOR4xp25_ASAP7_75t_SL g1165 ( 
.A(n_954),
.B(n_946),
.C(n_1033),
.D(n_948),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_933),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_SL g1167 ( 
.A(n_928),
.B(n_951),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1060),
.A2(n_411),
.B(n_382),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_961),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_SL g1170 ( 
.A1(n_1024),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1079),
.A2(n_38),
.B(n_40),
.C(n_42),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1012),
.B(n_38),
.Y(n_1172)
);

INVx5_ASAP7_75t_L g1173 ( 
.A(n_1034),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_918),
.A2(n_411),
.B(n_382),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_923),
.A2(n_411),
.B(n_382),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_980),
.B(n_44),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_926),
.A2(n_411),
.B(n_382),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_936),
.B(n_45),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_983),
.Y(n_1179)
);

OAI22x1_ASAP7_75t_L g1180 ( 
.A1(n_983),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1037),
.A2(n_345),
.B(n_542),
.C(n_535),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1073),
.A2(n_560),
.B(n_542),
.C(n_520),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_944),
.B(n_48),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_945),
.A2(n_49),
.B(n_50),
.C(n_52),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_SL g1185 ( 
.A(n_1067),
.B(n_55),
.C(n_56),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_955),
.B(n_58),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_1001),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_997),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_926),
.A2(n_520),
.B(n_560),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_965),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1061),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1047),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_997),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_932),
.A2(n_61),
.B(n_62),
.C(n_64),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1021),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1044),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_932),
.B(n_64),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1044),
.Y(n_1198)
);

INVxp67_ASAP7_75t_SL g1199 ( 
.A(n_967),
.Y(n_1199)
);

INVxp67_ASAP7_75t_L g1200 ( 
.A(n_1069),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1052),
.B(n_560),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_974),
.B(n_560),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_942),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1015),
.A2(n_560),
.B1(n_542),
.B2(n_520),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1084),
.A2(n_520),
.B(n_542),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1019),
.A2(n_542),
.B1(n_520),
.B2(n_88),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1042),
.B(n_520),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1017),
.A2(n_1042),
.B(n_957),
.C(n_952),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_969),
.A2(n_76),
.B(n_79),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_973),
.A2(n_97),
.B(n_117),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_941),
.A2(n_120),
.B(n_122),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_962),
.A2(n_134),
.B1(n_143),
.B2(n_144),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_987),
.A2(n_145),
.B1(n_150),
.B2(n_156),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1025),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_952),
.B(n_178),
.Y(n_1215)
);

AND3x1_ASAP7_75t_SL g1216 ( 
.A(n_1018),
.B(n_209),
.C(n_190),
.Y(n_1216)
);

XNOR2xp5_ASAP7_75t_L g1217 ( 
.A(n_1031),
.B(n_183),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1021),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_L g1219 ( 
.A(n_1029),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1026),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_938),
.A2(n_198),
.B1(n_207),
.B2(n_1050),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_938),
.B(n_1041),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1062),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1027),
.Y(n_1224)
);

NAND2x1p5_ASAP7_75t_L g1225 ( 
.A(n_1021),
.B(n_1076),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_973),
.A2(n_1085),
.B(n_1055),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1008),
.B(n_985),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1055),
.A2(n_1023),
.B(n_996),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_957),
.A2(n_964),
.B(n_939),
.C(n_1014),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1032),
.B(n_1036),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1023),
.A2(n_996),
.B(n_1002),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1021),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1049),
.B(n_975),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1066),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1035),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1068),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_976),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1038),
.B(n_1002),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1226),
.A2(n_1040),
.B(n_989),
.Y(n_1239)
);

INVx4_ASAP7_75t_SL g1240 ( 
.A(n_1232),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1103),
.B(n_1057),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1117),
.A2(n_1003),
.B(n_1022),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1118),
.A2(n_1003),
.B(n_1022),
.Y(n_1243)
);

CKINVDCx11_ASAP7_75t_R g1244 ( 
.A(n_1137),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1173),
.B(n_1045),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1116),
.A2(n_1071),
.B(n_1028),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1133),
.B(n_978),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1187),
.B(n_1155),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1109),
.A2(n_1040),
.B(n_989),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_L g1250 ( 
.A(n_1100),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1109),
.A2(n_1013),
.B(n_971),
.C(n_984),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1154),
.B(n_1054),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1231),
.A2(n_1028),
.B(n_1081),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1173),
.B(n_1088),
.Y(n_1254)
);

INVx4_ASAP7_75t_L g1255 ( 
.A(n_1173),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1150),
.B(n_1138),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1114),
.A2(n_986),
.B(n_949),
.Y(n_1257)
);

CKINVDCx20_ASAP7_75t_R g1258 ( 
.A(n_1099),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_SL g1259 ( 
.A1(n_1208),
.A2(n_916),
.B(n_1080),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1229),
.A2(n_916),
.B(n_1080),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1131),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1110),
.A2(n_963),
.B(n_1045),
.C(n_987),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1147),
.B(n_1075),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1228),
.A2(n_1081),
.B(n_1043),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1168),
.A2(n_1043),
.B(n_1059),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1164),
.A2(n_1065),
.B(n_1059),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1173),
.B(n_1000),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1101),
.A2(n_1010),
.B(n_1086),
.C(n_1007),
.Y(n_1268)
);

AOI221xp5_ASAP7_75t_SL g1269 ( 
.A1(n_1148),
.A2(n_1171),
.B1(n_1184),
.B2(n_1194),
.C(n_1190),
.Y(n_1269)
);

AOI221x1_ASAP7_75t_L g1270 ( 
.A1(n_1210),
.A2(n_1056),
.B1(n_1065),
.B2(n_1077),
.C(n_1051),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1106),
.B(n_1034),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1174),
.A2(n_1056),
.B(n_972),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1136),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1106),
.B(n_1034),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1156),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1091),
.A2(n_972),
.B(n_1051),
.Y(n_1276)
);

BUFx10_ASAP7_75t_L g1277 ( 
.A(n_1113),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1219),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1211),
.A2(n_1046),
.B(n_1034),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1130),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1091),
.B(n_1064),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1169),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1092),
.A2(n_1053),
.B(n_1095),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1111),
.A2(n_1215),
.B(n_1104),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1215),
.A2(n_1206),
.B(n_1097),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1225),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1203),
.A2(n_1143),
.B1(n_1200),
.B2(n_1144),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1181),
.A2(n_1177),
.A3(n_1175),
.B(n_1128),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1158),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1153),
.B(n_1089),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1097),
.A2(n_1157),
.B(n_1197),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1202),
.A2(n_1123),
.B(n_1205),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1182),
.A2(n_1105),
.A3(n_1238),
.B(n_1233),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1125),
.A2(n_1202),
.B(n_1105),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1124),
.A2(n_1108),
.B(n_1238),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1132),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1189),
.A2(n_1145),
.B(n_1207),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1120),
.B(n_1108),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1232),
.Y(n_1299)
);

AOI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1197),
.A2(n_1201),
.B(n_1145),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1301)
);

NOR3xp33_ASAP7_75t_L g1302 ( 
.A(n_1151),
.B(n_1176),
.C(n_1141),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1201),
.A2(n_1212),
.B(n_1209),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1094),
.A2(n_1096),
.B1(n_1129),
.B2(n_1126),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1230),
.B(n_1214),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1232),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1178),
.A2(n_1186),
.B1(n_1183),
.B2(n_1221),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1230),
.A2(n_1163),
.B(n_1160),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1160),
.A2(n_1172),
.B(n_1162),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1098),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1179),
.B(n_1115),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1220),
.B(n_1235),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1140),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1224),
.B(n_1152),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1115),
.B(n_1198),
.Y(n_1315)
);

NOR2xp67_ASAP7_75t_SL g1316 ( 
.A(n_1100),
.B(n_1218),
.Y(n_1316)
);

AND3x4_ASAP7_75t_L g1317 ( 
.A(n_1185),
.B(n_1135),
.C(n_1127),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1162),
.A2(n_1172),
.B(n_1163),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1191),
.A2(n_1236),
.B1(n_1234),
.B2(n_1223),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1227),
.B(n_1222),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1170),
.A2(n_1186),
.B(n_1134),
.C(n_1139),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1121),
.A2(n_1090),
.B(n_1161),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1146),
.A2(n_1192),
.B(n_1112),
.Y(n_1323)
);

CKINVDCx11_ASAP7_75t_R g1324 ( 
.A(n_1100),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1121),
.A2(n_1090),
.B(n_1161),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_L g1326 ( 
.A(n_1217),
.B(n_1122),
.C(n_1119),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1165),
.B(n_1237),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_SL g1328 ( 
.A1(n_1142),
.A2(n_1199),
.B(n_1213),
.C(n_1218),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_SL g1329 ( 
.A(n_1098),
.B(n_1167),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1180),
.B(n_1159),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1216),
.A2(n_1204),
.A3(n_1149),
.B(n_1196),
.Y(n_1331)
);

BUFx12f_ASAP7_75t_L g1332 ( 
.A(n_1166),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1188),
.B(n_1193),
.Y(n_1333)
);

NOR4xp25_ASAP7_75t_L g1334 ( 
.A(n_1195),
.B(n_1237),
.C(n_1193),
.D(n_1188),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1196),
.A2(n_956),
.B(n_689),
.C(n_1109),
.Y(n_1335)
);

OAI22x1_ASAP7_75t_L g1336 ( 
.A1(n_1102),
.A2(n_642),
.B1(n_921),
.B2(n_868),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1103),
.B(n_803),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1091),
.B(n_1109),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1232),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1226),
.A2(n_1109),
.B(n_1107),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1131),
.Y(n_1341)
);

AND2x6_ASAP7_75t_L g1342 ( 
.A(n_1232),
.B(n_1009),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1133),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1131),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1091),
.B(n_1109),
.Y(n_1345)
);

BUFx12f_ASAP7_75t_L g1346 ( 
.A(n_1113),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1226),
.A2(n_1107),
.B(n_1168),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1091),
.B(n_1109),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_SL g1349 ( 
.A(n_1173),
.B(n_1070),
.Y(n_1349)
);

OAI22x1_ASAP7_75t_L g1350 ( 
.A1(n_1102),
.A2(n_642),
.B1(n_921),
.B2(n_868),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1226),
.A2(n_1109),
.B(n_1107),
.Y(n_1351)
);

BUFx2_ASAP7_75t_R g1352 ( 
.A(n_1099),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1226),
.A2(n_956),
.B(n_1114),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1226),
.A2(n_1107),
.B(n_1168),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1091),
.B(n_1109),
.Y(n_1355)
);

AOI31xp33_ASAP7_75t_L g1356 ( 
.A1(n_1103),
.A2(n_1074),
.A3(n_1070),
.B(n_956),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1226),
.A2(n_956),
.B(n_1114),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1148),
.A2(n_642),
.B(n_956),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1103),
.B(n_1133),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1103),
.B(n_917),
.Y(n_1360)
);

NAND3xp33_ASAP7_75t_L g1361 ( 
.A(n_1143),
.B(n_632),
.C(n_956),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1091),
.B(n_1109),
.Y(n_1362)
);

NOR2xp67_ASAP7_75t_L g1363 ( 
.A(n_1187),
.B(n_857),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1091),
.B(n_1109),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1117),
.A2(n_1118),
.B(n_1116),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1091),
.B(n_1109),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1117),
.A2(n_1118),
.B(n_1116),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1117),
.A2(n_1118),
.B(n_1116),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1226),
.A2(n_1109),
.B(n_1107),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1226),
.A2(n_1109),
.B(n_1107),
.Y(n_1370)
);

AOI21xp33_ASAP7_75t_L g1371 ( 
.A1(n_1103),
.A2(n_1074),
.B(n_1070),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1226),
.A2(n_1109),
.B(n_1107),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1226),
.A2(n_1109),
.B(n_1107),
.Y(n_1373)
);

OAI21xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1211),
.A2(n_1157),
.B(n_1109),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1103),
.B(n_803),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1091),
.B(n_1109),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1103),
.B(n_813),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1093),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1232),
.Y(n_1379)
);

NOR2x1_ASAP7_75t_L g1380 ( 
.A(n_1136),
.B(n_803),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_1133),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1226),
.A2(n_1109),
.B(n_1107),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1117),
.A2(n_1118),
.B(n_1116),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1226),
.A2(n_1109),
.B(n_1107),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1361),
.A2(n_1377),
.B1(n_1241),
.B2(n_1358),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1383),
.A2(n_1292),
.B(n_1347),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1354),
.A2(n_1284),
.B(n_1272),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1353),
.A2(n_1357),
.B(n_1270),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1359),
.B(n_1343),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1293),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_L g1392 ( 
.A(n_1358),
.B(n_1302),
.C(n_1326),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1244),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1256),
.B(n_1320),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1242),
.A2(n_1297),
.B(n_1243),
.Y(n_1395)
);

A2O1A1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1374),
.A2(n_1356),
.B(n_1307),
.C(n_1335),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1353),
.A2(n_1357),
.B(n_1285),
.Y(n_1397)
);

AOI222xp33_ASAP7_75t_L g1398 ( 
.A1(n_1336),
.A2(n_1350),
.B1(n_1330),
.B2(n_1287),
.C1(n_1252),
.C2(n_1307),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1239),
.A2(n_1303),
.B(n_1340),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1265),
.A2(n_1253),
.B(n_1264),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1246),
.A2(n_1266),
.B(n_1300),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1295),
.A2(n_1309),
.B(n_1351),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1369),
.A2(n_1372),
.B(n_1370),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_SL g1404 ( 
.A1(n_1318),
.A2(n_1279),
.B(n_1373),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1382),
.A2(n_1384),
.B(n_1259),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1261),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1283),
.A2(n_1276),
.B(n_1257),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1258),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1290),
.B(n_1360),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1371),
.A2(n_1301),
.B1(n_1345),
.B2(n_1366),
.Y(n_1410)
);

OAI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1356),
.A2(n_1362),
.B1(n_1376),
.B2(n_1338),
.Y(n_1411)
);

NAND2x1p5_ASAP7_75t_L g1412 ( 
.A(n_1255),
.B(n_1316),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1346),
.Y(n_1413)
);

AND2x6_ASAP7_75t_L g1414 ( 
.A(n_1327),
.B(n_1286),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1308),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1318),
.A2(n_1291),
.B(n_1283),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_SL g1417 ( 
.A(n_1352),
.B(n_1349),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1328),
.A2(n_1260),
.B(n_1348),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1308),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1251),
.A2(n_1262),
.B(n_1281),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1337),
.A2(n_1375),
.B1(n_1371),
.B2(n_1304),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1294),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1294),
.A2(n_1325),
.B(n_1322),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1327),
.A2(n_1334),
.B(n_1305),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1281),
.A2(n_1355),
.B(n_1362),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1275),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1305),
.A2(n_1245),
.B(n_1274),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1289),
.Y(n_1428)
);

OAI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1364),
.A2(n_1376),
.B(n_1366),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1245),
.A2(n_1271),
.B(n_1312),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1269),
.A2(n_1268),
.B(n_1312),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1323),
.A2(n_1321),
.B(n_1254),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1364),
.B(n_1298),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1267),
.A2(n_1323),
.B(n_1310),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1293),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1314),
.A2(n_1341),
.B(n_1344),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1282),
.Y(n_1437)
);

INVx5_ASAP7_75t_L g1438 ( 
.A(n_1342),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1280),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1296),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1333),
.A2(n_1319),
.B(n_1313),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1263),
.A2(n_1288),
.B(n_1380),
.Y(n_1442)
);

NAND2x1p5_ASAP7_75t_L g1443 ( 
.A(n_1255),
.B(n_1250),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1288),
.A2(n_1247),
.B(n_1293),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1288),
.A2(n_1248),
.B(n_1329),
.Y(n_1445)
);

AO21x1_ASAP7_75t_L g1446 ( 
.A1(n_1349),
.A2(n_1329),
.B(n_1278),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1342),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1331),
.A2(n_1342),
.B(n_1240),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1273),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1331),
.A2(n_1315),
.B(n_1342),
.Y(n_1450)
);

AOI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1311),
.A2(n_1363),
.B(n_1378),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1331),
.A2(n_1240),
.B(n_1299),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1240),
.A2(n_1299),
.B(n_1339),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1306),
.A2(n_1339),
.B(n_1379),
.Y(n_1454)
);

OR2x6_ASAP7_75t_L g1455 ( 
.A(n_1306),
.B(n_1339),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1317),
.A2(n_1379),
.B1(n_1332),
.B2(n_1277),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1282),
.Y(n_1457)
);

AOI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1358),
.A2(n_566),
.B1(n_876),
.B2(n_498),
.C(n_642),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1293),
.Y(n_1459)
);

OAI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1358),
.A2(n_642),
.B1(n_632),
.B2(n_566),
.C(n_1361),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1294),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1371),
.A2(n_1070),
.B1(n_1074),
.B2(n_876),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1261),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1371),
.A2(n_1070),
.B1(n_1074),
.B2(n_876),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1285),
.A2(n_1284),
.B(n_1318),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1361),
.A2(n_632),
.B(n_956),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1361),
.A2(n_1377),
.B1(n_1241),
.B2(n_956),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1374),
.A2(n_1358),
.B(n_1361),
.C(n_956),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1244),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1327),
.B(n_1254),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1244),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1240),
.B(n_1333),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1261),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1371),
.A2(n_1070),
.B1(n_1074),
.B2(n_876),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1300),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1374),
.B(n_1249),
.Y(n_1477)
);

OAI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1358),
.A2(n_642),
.B1(n_632),
.B2(n_566),
.C(n_1361),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1327),
.B(n_1254),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1381),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1361),
.A2(n_1377),
.B1(n_1241),
.B2(n_956),
.Y(n_1482)
);

OAI21xp33_ASAP7_75t_L g1483 ( 
.A1(n_1361),
.A2(n_632),
.B(n_566),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1285),
.A2(n_1284),
.B(n_1318),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1261),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1359),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1256),
.B(n_1320),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1261),
.Y(n_1488)
);

AO32x2_ASAP7_75t_L g1489 ( 
.A1(n_1307),
.A2(n_1103),
.A3(n_1190),
.B1(n_1030),
.B2(n_885),
.Y(n_1489)
);

INVx5_ASAP7_75t_L g1490 ( 
.A(n_1342),
.Y(n_1490)
);

AO32x2_ASAP7_75t_L g1491 ( 
.A1(n_1307),
.A2(n_1103),
.A3(n_1190),
.B1(n_1030),
.B2(n_885),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1306),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1374),
.A2(n_1239),
.B(n_1284),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1300),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1256),
.B(n_1320),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1374),
.A2(n_1358),
.B(n_1361),
.C(n_956),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1324),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1338),
.B(n_1345),
.Y(n_1501)
);

INVx5_ASAP7_75t_L g1502 ( 
.A(n_1342),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1293),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1361),
.A2(n_632),
.B(n_956),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1359),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1338),
.B(n_1345),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1261),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1371),
.A2(n_1070),
.B1(n_1074),
.B2(n_876),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1261),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1377),
.A2(n_1317),
.B1(n_642),
.B2(n_580),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1255),
.B(n_1173),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1293),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1306),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1358),
.B(n_1361),
.C(n_1241),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1282),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1371),
.A2(n_1070),
.B1(n_1074),
.B2(n_876),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1358),
.A2(n_632),
.B(n_1361),
.C(n_1241),
.Y(n_1520)
);

AO31x2_ASAP7_75t_L g1521 ( 
.A1(n_1270),
.A2(n_1285),
.A3(n_1284),
.B(n_1266),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1300),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1338),
.B(n_1345),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1365),
.A2(n_1368),
.B(n_1367),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1361),
.A2(n_632),
.B(n_956),
.Y(n_1525)
);

BUFx12f_ASAP7_75t_L g1526 ( 
.A(n_1244),
.Y(n_1526)
);

AOI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1284),
.A2(n_1354),
.B(n_1347),
.Y(n_1527)
);

NAND2x1p5_ASAP7_75t_L g1528 ( 
.A(n_1255),
.B(n_1173),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1377),
.A2(n_1063),
.B1(n_876),
.B2(n_865),
.Y(n_1529)
);

INVxp33_ASAP7_75t_L g1530 ( 
.A(n_1394),
.Y(n_1530)
);

NOR2xp67_ASAP7_75t_L g1531 ( 
.A(n_1486),
.B(n_1507),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1471),
.B(n_1479),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1406),
.Y(n_1533)
);

A2O1A1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1460),
.A2(n_1478),
.B(n_1458),
.C(n_1520),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1409),
.B(n_1487),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1467),
.A2(n_1482),
.B(n_1385),
.C(n_1483),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1497),
.B(n_1486),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1494),
.A2(n_1399),
.B(n_1388),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1468),
.A2(n_1498),
.B(n_1520),
.C(n_1396),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1507),
.B(n_1390),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1392),
.A2(n_1396),
.B1(n_1468),
.B2(n_1498),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1516),
.A2(n_1411),
.B(n_1466),
.C(n_1525),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1516),
.A2(n_1506),
.B(n_1411),
.Y(n_1543)
);

O2A1O1Ixp5_ASAP7_75t_L g1544 ( 
.A1(n_1420),
.A2(n_1418),
.B(n_1446),
.C(n_1477),
.Y(n_1544)
);

O2A1O1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1477),
.A2(n_1404),
.B(n_1425),
.C(n_1418),
.Y(n_1545)
);

A2O1A1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1529),
.A2(n_1421),
.B(n_1462),
.C(n_1510),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1481),
.Y(n_1547)
);

AOI221x1_ASAP7_75t_SL g1548 ( 
.A1(n_1456),
.A2(n_1512),
.B1(n_1489),
.B2(n_1491),
.C(n_1523),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1410),
.B(n_1429),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1433),
.B(n_1426),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_SL g1551 ( 
.A1(n_1412),
.A2(n_1431),
.B(n_1513),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1473),
.B(n_1438),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1410),
.B(n_1428),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1462),
.A2(n_1475),
.B1(n_1519),
.B2(n_1510),
.Y(n_1554)
);

NAND4xp25_ASAP7_75t_L g1555 ( 
.A(n_1398),
.B(n_1475),
.C(n_1464),
.D(n_1519),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1463),
.B(n_1474),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1464),
.A2(n_1405),
.B(n_1508),
.C(n_1501),
.Y(n_1557)
);

OA22x2_ASAP7_75t_L g1558 ( 
.A1(n_1471),
.A2(n_1479),
.B1(n_1485),
.B2(n_1511),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1424),
.B(n_1416),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1488),
.B(n_1509),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1438),
.B(n_1490),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1436),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1391),
.A2(n_1435),
.B1(n_1459),
.B2(n_1504),
.C(n_1514),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1424),
.B(n_1416),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1393),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1500),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1397),
.A2(n_1484),
.B(n_1465),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1386),
.A2(n_1469),
.B(n_1499),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1439),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1480),
.A2(n_1505),
.B(n_1503),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1518),
.A2(n_1524),
.B(n_1402),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1491),
.B(n_1417),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1389),
.A2(n_1502),
.B1(n_1500),
.B2(n_1471),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1444),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1440),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1457),
.A2(n_1517),
.B(n_1389),
.C(n_1435),
.Y(n_1576)
);

CKINVDCx11_ASAP7_75t_R g1577 ( 
.A(n_1472),
.Y(n_1577)
);

O2A1O1Ixp5_ASAP7_75t_L g1578 ( 
.A1(n_1451),
.A2(n_1515),
.B(n_1492),
.C(n_1447),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1442),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1461),
.A2(n_1403),
.B(n_1407),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1427),
.B(n_1414),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1454),
.B(n_1455),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1454),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1414),
.B(n_1459),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1443),
.A2(n_1472),
.B1(n_1408),
.B2(n_1470),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1443),
.A2(n_1408),
.B1(n_1470),
.B2(n_1449),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1414),
.B(n_1430),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1448),
.B(n_1445),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1430),
.B(n_1450),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1528),
.A2(n_1450),
.B(n_1476),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1414),
.B(n_1450),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1449),
.A2(n_1422),
.B1(n_1526),
.B2(n_1413),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1476),
.A2(n_1522),
.B(n_1496),
.C(n_1422),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1413),
.A2(n_1522),
.B1(n_1496),
.B2(n_1419),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1415),
.A2(n_1527),
.B1(n_1493),
.B2(n_1495),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1452),
.B(n_1453),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1432),
.B(n_1521),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1452),
.B(n_1441),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1432),
.B(n_1434),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1423),
.B(n_1521),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1493),
.A2(n_1495),
.B1(n_1521),
.B2(n_1401),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1521),
.B(n_1493),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1395),
.Y(n_1603)
);

OA21x2_ASAP7_75t_L g1604 ( 
.A1(n_1400),
.A2(n_1494),
.B(n_1399),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1495),
.B(n_1390),
.Y(n_1605)
);

OA21x2_ASAP7_75t_L g1606 ( 
.A1(n_1494),
.A2(n_1399),
.B(n_1387),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1385),
.A2(n_1478),
.B1(n_1460),
.B2(n_1392),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1512),
.A2(n_1377),
.B1(n_1529),
.B2(n_1317),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1385),
.A2(n_1478),
.B1(n_1460),
.B2(n_1392),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1409),
.B(n_1394),
.Y(n_1610)
);

OA21x2_ASAP7_75t_L g1611 ( 
.A1(n_1494),
.A2(n_1399),
.B(n_1387),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1409),
.B(n_1394),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1437),
.Y(n_1613)
);

O2A1O1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1460),
.A2(n_1478),
.B(n_1482),
.C(n_1467),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1409),
.B(n_1394),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1409),
.B(n_1394),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1494),
.A2(n_1374),
.B(n_1405),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1437),
.Y(n_1618)
);

BUFx4f_ASAP7_75t_SL g1619 ( 
.A(n_1393),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1385),
.A2(n_1478),
.B1(n_1460),
.B2(n_1392),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1494),
.A2(n_1374),
.B(n_1405),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1473),
.B(n_1438),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1486),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1486),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1409),
.B(n_1394),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1385),
.A2(n_1478),
.B1(n_1460),
.B2(n_1392),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1385),
.A2(n_1478),
.B1(n_1460),
.B2(n_1392),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1533),
.Y(n_1628)
);

OR2x6_ASAP7_75t_L g1629 ( 
.A(n_1590),
.B(n_1532),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1617),
.A2(n_1621),
.B(n_1567),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1588),
.B(n_1589),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1541),
.A2(n_1534),
.B1(n_1626),
.B2(n_1620),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1549),
.B(n_1548),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1549),
.B(n_1548),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1562),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1599),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1537),
.B(n_1605),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1580),
.A2(n_1601),
.B(n_1595),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1572),
.B(n_1623),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1600),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1559),
.Y(n_1641)
);

AOI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1595),
.A2(n_1597),
.B(n_1601),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1581),
.B(n_1582),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1624),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1531),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1540),
.B(n_1556),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1553),
.B(n_1547),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1547),
.B(n_1564),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1557),
.B(n_1550),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1569),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1597),
.A2(n_1602),
.B(n_1544),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1575),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1560),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1535),
.B(n_1610),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1612),
.B(n_1615),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1581),
.B(n_1587),
.Y(n_1656)
);

BUFx12f_ASAP7_75t_L g1657 ( 
.A(n_1577),
.Y(n_1657)
);

OA21x2_ASAP7_75t_L g1658 ( 
.A1(n_1603),
.A2(n_1591),
.B(n_1579),
.Y(n_1658)
);

AO21x2_ASAP7_75t_L g1659 ( 
.A1(n_1594),
.A2(n_1593),
.B(n_1576),
.Y(n_1659)
);

INVx5_ASAP7_75t_L g1660 ( 
.A(n_1561),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1584),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1536),
.B(n_1541),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1563),
.A2(n_1584),
.B(n_1574),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1616),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1546),
.A2(n_1543),
.B(n_1598),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1625),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1596),
.B(n_1552),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1583),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1539),
.B(n_1545),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1568),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1614),
.B(n_1542),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1604),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1558),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1558),
.Y(n_1674)
);

AO21x2_ASAP7_75t_L g1675 ( 
.A1(n_1554),
.A2(n_1627),
.B(n_1626),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1607),
.B(n_1627),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1578),
.A2(n_1573),
.B(n_1620),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1530),
.B(n_1592),
.Y(n_1678)
);

AO21x2_ASAP7_75t_L g1679 ( 
.A1(n_1554),
.A2(n_1609),
.B(n_1607),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1660),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1640),
.B(n_1538),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1640),
.B(n_1631),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1635),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1635),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1648),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1631),
.B(n_1622),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1645),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1675),
.A2(n_1555),
.B1(n_1609),
.B2(n_1608),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1670),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1628),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1670),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1658),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1675),
.A2(n_1555),
.B1(n_1592),
.B2(n_1586),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1661),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1658),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1658),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1631),
.B(n_1636),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1631),
.B(n_1636),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1675),
.A2(n_1586),
.B1(n_1585),
.B2(n_1532),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1647),
.B(n_1571),
.Y(n_1702)
);

OR2x6_ASAP7_75t_L g1703 ( 
.A(n_1629),
.B(n_1551),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1675),
.A2(n_1585),
.B1(n_1532),
.B2(n_1619),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1661),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1656),
.B(n_1570),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1656),
.B(n_1570),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1695),
.A2(n_1632),
.B1(n_1676),
.B2(n_1662),
.Y(n_1708)
);

OA21x2_ASAP7_75t_L g1709 ( 
.A1(n_1694),
.A2(n_1638),
.B(n_1672),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1680),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1694),
.A2(n_1633),
.B(n_1634),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1689),
.A2(n_1679),
.B1(n_1634),
.B2(n_1665),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1688),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1683),
.Y(n_1715)
);

NOR3xp33_ASAP7_75t_L g1716 ( 
.A(n_1691),
.B(n_1632),
.C(n_1676),
.Y(n_1716)
);

OAI22xp33_ASAP7_75t_SL g1717 ( 
.A1(n_1701),
.A2(n_1649),
.B1(n_1678),
.B2(n_1673),
.Y(n_1717)
);

OAI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1689),
.A2(n_1671),
.B1(n_1649),
.B2(n_1669),
.C(n_1677),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1695),
.A2(n_1671),
.B1(n_1679),
.B2(n_1669),
.C(n_1641),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1701),
.A2(n_1677),
.B(n_1678),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1691),
.A2(n_1679),
.B1(n_1641),
.B2(n_1665),
.C(n_1639),
.Y(n_1721)
);

NAND4xp25_ASAP7_75t_SL g1722 ( 
.A(n_1701),
.B(n_1679),
.C(n_1654),
.D(n_1655),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1698),
.A2(n_1665),
.B1(n_1639),
.B2(n_1650),
.C(n_1652),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1704),
.A2(n_1665),
.B1(n_1673),
.B2(n_1674),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1692),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1705),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1692),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_SL g1728 ( 
.A1(n_1704),
.A2(n_1657),
.B1(n_1565),
.B2(n_1566),
.Y(n_1728)
);

AO21x2_ASAP7_75t_L g1729 ( 
.A1(n_1697),
.A2(n_1642),
.B(n_1668),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1682),
.B(n_1637),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1682),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1696),
.B(n_1644),
.Y(n_1732)
);

OAI31xp33_ASAP7_75t_SL g1733 ( 
.A1(n_1688),
.A2(n_1700),
.A3(n_1699),
.B(n_1684),
.Y(n_1733)
);

NAND2xp33_ASAP7_75t_R g1734 ( 
.A(n_1687),
.B(n_1677),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_SL g1735 ( 
.A(n_1699),
.B(n_1654),
.C(n_1655),
.D(n_1657),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1699),
.B(n_1646),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1685),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1696),
.B(n_1677),
.C(n_1663),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1705),
.B(n_1646),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1680),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1686),
.B(n_1664),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1686),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1702),
.B(n_1653),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1703),
.A2(n_1643),
.B1(n_1659),
.B2(n_1667),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_L g1745 ( 
.A(n_1719),
.B(n_1698),
.C(n_1630),
.Y(n_1745)
);

OAI21xp33_ASAP7_75t_L g1746 ( 
.A1(n_1716),
.A2(n_1684),
.B(n_1681),
.Y(n_1746)
);

BUFx2_ASAP7_75t_L g1747 ( 
.A(n_1711),
.Y(n_1747)
);

CKINVDCx8_ASAP7_75t_R g1748 ( 
.A(n_1714),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1726),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1725),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1727),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1715),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1708),
.A2(n_1630),
.B(n_1651),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1709),
.Y(n_1754)
);

NOR2x1p5_ASAP7_75t_L g1755 ( 
.A(n_1714),
.B(n_1680),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1733),
.B(n_1700),
.Y(n_1756)
);

AOI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1738),
.A2(n_1693),
.B(n_1690),
.Y(n_1757)
);

INVx4_ASAP7_75t_SL g1758 ( 
.A(n_1728),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1709),
.Y(n_1759)
);

OAI21x1_ASAP7_75t_L g1760 ( 
.A1(n_1720),
.A2(n_1690),
.B(n_1693),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1715),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1732),
.Y(n_1762)
);

AND2x2_ASAP7_75t_SL g1763 ( 
.A(n_1713),
.B(n_1721),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1731),
.B(n_1706),
.Y(n_1764)
);

INVx4_ASAP7_75t_L g1765 ( 
.A(n_1740),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1712),
.Y(n_1766)
);

INVx4_ASAP7_75t_SL g1767 ( 
.A(n_1740),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1709),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1729),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1729),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1712),
.B(n_1706),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1712),
.Y(n_1772)
);

AND2x2_ASAP7_75t_SL g1773 ( 
.A(n_1723),
.B(n_1630),
.Y(n_1773)
);

AOI21xp33_ASAP7_75t_L g1774 ( 
.A1(n_1718),
.A2(n_1659),
.B(n_1630),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1745),
.B(n_1722),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1750),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1748),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1766),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1756),
.B(n_1707),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1745),
.B(n_1742),
.Y(n_1780)
);

NOR2x1_ASAP7_75t_L g1781 ( 
.A(n_1765),
.B(n_1735),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1767),
.B(n_1740),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1754),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1754),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1748),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1750),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1763),
.B(n_1737),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1749),
.B(n_1743),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1767),
.B(n_1771),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1754),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1751),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1754),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1767),
.B(n_1736),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1767),
.B(n_1736),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1767),
.B(n_1710),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1748),
.B(n_1666),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1766),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1763),
.B(n_1737),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1763),
.B(n_1743),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1747),
.Y(n_1800)
);

INVx5_ASAP7_75t_L g1801 ( 
.A(n_1754),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1751),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1759),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1752),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1759),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1772),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1752),
.Y(n_1807)
);

NOR2xp67_ASAP7_75t_L g1808 ( 
.A(n_1765),
.B(n_1744),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1761),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1759),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1771),
.B(n_1764),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1771),
.B(n_1710),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1747),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1764),
.B(n_1730),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1776),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1799),
.B(n_1762),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1785),
.B(n_1746),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1785),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1776),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1799),
.B(n_1762),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1786),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1787),
.B(n_1798),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1775),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1786),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1791),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1791),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1782),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1787),
.B(n_1741),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1777),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1793),
.B(n_1755),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1798),
.B(n_1739),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1802),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1783),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1782),
.B(n_1755),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1813),
.B(n_1763),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1802),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1782),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1813),
.B(n_1746),
.Y(n_1838)
);

OAI33xp33_ASAP7_75t_L g1839 ( 
.A1(n_1775),
.A2(n_1717),
.A3(n_1769),
.B1(n_1770),
.B2(n_1759),
.B3(n_1768),
.Y(n_1839)
);

NAND2x1p5_ASAP7_75t_L g1840 ( 
.A(n_1782),
.B(n_1566),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1788),
.B(n_1753),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1775),
.B(n_1773),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1796),
.B(n_1773),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1796),
.B(n_1773),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1804),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1804),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1780),
.B(n_1773),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1782),
.B(n_1758),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1793),
.B(n_1747),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1807),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1783),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1823),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1849),
.B(n_1777),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1845),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1823),
.B(n_1842),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1827),
.B(n_1777),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1829),
.B(n_1777),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1822),
.B(n_1788),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1839),
.A2(n_1774),
.B1(n_1753),
.B2(n_1724),
.Y(n_1859)
);

INVx1_ASAP7_75t_SL g1860 ( 
.A(n_1818),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1846),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1847),
.A2(n_1774),
.B1(n_1780),
.B2(n_1803),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1850),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1849),
.B(n_1793),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1816),
.B(n_1788),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1817),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1833),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1829),
.B(n_1812),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1815),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1819),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1821),
.Y(n_1871)
);

AOI21xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1848),
.A2(n_1789),
.B(n_1794),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1834),
.B(n_1794),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1848),
.B(n_1827),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1820),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1824),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1825),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1834),
.B(n_1794),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1837),
.Y(n_1879)
);

OAI221xp5_ASAP7_75t_SL g1880 ( 
.A1(n_1852),
.A2(n_1835),
.B1(n_1844),
.B2(n_1843),
.C(n_1841),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1861),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1861),
.Y(n_1882)
);

AOI221xp5_ASAP7_75t_L g1883 ( 
.A1(n_1859),
.A2(n_1817),
.B1(n_1838),
.B2(n_1772),
.C(n_1805),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_SL g1884 ( 
.A1(n_1875),
.A2(n_1789),
.B1(n_1811),
.B2(n_1779),
.Y(n_1884)
);

OAI31xp33_ASAP7_75t_SL g1885 ( 
.A1(n_1874),
.A2(n_1789),
.A3(n_1781),
.B(n_1830),
.Y(n_1885)
);

OAI221xp5_ASAP7_75t_L g1886 ( 
.A1(n_1862),
.A2(n_1808),
.B1(n_1734),
.B2(n_1837),
.C(n_1757),
.Y(n_1886)
);

OAI22xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1855),
.A2(n_1757),
.B1(n_1801),
.B2(n_1840),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1860),
.B(n_1853),
.Y(n_1888)
);

OAI21xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1864),
.A2(n_1811),
.B(n_1779),
.Y(n_1889)
);

OAI321xp33_ASAP7_75t_L g1890 ( 
.A1(n_1855),
.A2(n_1810),
.A3(n_1803),
.B1(n_1805),
.B2(n_1811),
.C(n_1792),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1863),
.Y(n_1891)
);

AOI21xp33_ASAP7_75t_SL g1892 ( 
.A1(n_1866),
.A2(n_1840),
.B(n_1795),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1865),
.B(n_1828),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1864),
.A2(n_1808),
.B1(n_1770),
.B2(n_1769),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1863),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1870),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1870),
.Y(n_1897)
);

OAI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1865),
.A2(n_1801),
.B1(n_1831),
.B2(n_1770),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1853),
.B(n_1814),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1856),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1877),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1883),
.B(n_1877),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1893),
.Y(n_1903)
);

INVx4_ASAP7_75t_L g1904 ( 
.A(n_1881),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1900),
.B(n_1888),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1899),
.B(n_1856),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1883),
.B(n_1879),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1885),
.B(n_1856),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1882),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1880),
.B(n_1857),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1891),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1895),
.B(n_1873),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1884),
.B(n_1868),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1896),
.Y(n_1914)
);

NOR2x1_ASAP7_75t_L g1915 ( 
.A(n_1897),
.B(n_1800),
.Y(n_1915)
);

OAI211xp5_ASAP7_75t_L g1916 ( 
.A1(n_1910),
.A2(n_1880),
.B(n_1872),
.C(n_1892),
.Y(n_1916)
);

NAND3xp33_ASAP7_75t_SL g1917 ( 
.A(n_1905),
.B(n_1886),
.C(n_1894),
.Y(n_1917)
);

AO21x1_ASAP7_75t_L g1918 ( 
.A1(n_1905),
.A2(n_1901),
.B(n_1887),
.Y(n_1918)
);

NOR4xp25_ASAP7_75t_L g1919 ( 
.A(n_1902),
.B(n_1890),
.C(n_1889),
.D(n_1898),
.Y(n_1919)
);

O2A1O1Ixp33_ASAP7_75t_L g1920 ( 
.A1(n_1902),
.A2(n_1867),
.B(n_1869),
.C(n_1854),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1912),
.B(n_1858),
.Y(n_1921)
);

OAI211xp5_ASAP7_75t_L g1922 ( 
.A1(n_1907),
.A2(n_1858),
.B(n_1878),
.C(n_1873),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1908),
.A2(n_1913),
.B(n_1911),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1903),
.A2(n_1867),
.B1(n_1876),
.B2(n_1871),
.C(n_1803),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1906),
.A2(n_1878),
.B(n_1760),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1912),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1909),
.B(n_1800),
.Y(n_1927)
);

AOI322xp5_ASAP7_75t_L g1928 ( 
.A1(n_1914),
.A2(n_1769),
.A3(n_1770),
.B1(n_1803),
.B2(n_1805),
.C1(n_1810),
.C2(n_1768),
.Y(n_1928)
);

OAI322xp33_ASAP7_75t_L g1929 ( 
.A1(n_1923),
.A2(n_1904),
.A3(n_1778),
.B1(n_1806),
.B2(n_1797),
.C1(n_1833),
.C2(n_1851),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1918),
.B(n_1904),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1926),
.B(n_1915),
.Y(n_1931)
);

AOI211xp5_ASAP7_75t_L g1932 ( 
.A1(n_1919),
.A2(n_1778),
.B(n_1797),
.C(n_1806),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1921),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1922),
.B(n_1800),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1927),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1924),
.Y(n_1936)
);

NOR2x1p5_ASAP7_75t_L g1937 ( 
.A(n_1933),
.B(n_1917),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1931),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1930),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1930),
.Y(n_1940)
);

NOR2x1p5_ASAP7_75t_L g1941 ( 
.A(n_1935),
.B(n_1800),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1934),
.B(n_1916),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1936),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1929),
.Y(n_1944)
);

AOI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1943),
.A2(n_1932),
.B1(n_1920),
.B2(n_1925),
.C(n_1805),
.Y(n_1945)
);

OAI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1939),
.A2(n_1928),
.B(n_1801),
.C(n_1851),
.Y(n_1946)
);

NOR2x1_ASAP7_75t_L g1947 ( 
.A(n_1940),
.B(n_1781),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1941),
.Y(n_1948)
);

AOI211xp5_ASAP7_75t_L g1949 ( 
.A1(n_1944),
.A2(n_1836),
.B(n_1832),
.C(n_1826),
.Y(n_1949)
);

BUFx12f_ASAP7_75t_L g1950 ( 
.A(n_1937),
.Y(n_1950)
);

NOR2xp67_ASAP7_75t_L g1951 ( 
.A(n_1950),
.B(n_1938),
.Y(n_1951)
);

A2O1A1Ixp33_ASAP7_75t_L g1952 ( 
.A1(n_1945),
.A2(n_1943),
.B(n_1942),
.C(n_1810),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1947),
.B(n_1801),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1951),
.Y(n_1954)
);

OAI211xp5_ASAP7_75t_L g1955 ( 
.A1(n_1954),
.A2(n_1952),
.B(n_1949),
.C(n_1948),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1955),
.A2(n_1953),
.B1(n_1810),
.B2(n_1784),
.Y(n_1956)
);

OR4x1_ASAP7_75t_L g1957 ( 
.A(n_1955),
.B(n_1946),
.C(n_1807),
.D(n_1809),
.Y(n_1957)
);

AOI221x1_ASAP7_75t_L g1958 ( 
.A1(n_1957),
.A2(n_1784),
.B1(n_1783),
.B2(n_1790),
.C(n_1792),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1956),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_SL g1960 ( 
.A1(n_1958),
.A2(n_1784),
.B(n_1783),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1959),
.A2(n_1792),
.B1(n_1784),
.B2(n_1790),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1961),
.Y(n_1962)
);

AO21x2_ASAP7_75t_L g1963 ( 
.A1(n_1962),
.A2(n_1960),
.B(n_1792),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1963),
.B(n_1801),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1964),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1965),
.A2(n_1790),
.B1(n_1801),
.B2(n_1779),
.Y(n_1966)
);

AOI211xp5_ASAP7_75t_L g1967 ( 
.A1(n_1966),
.A2(n_1790),
.B(n_1618),
.C(n_1613),
.Y(n_1967)
);


endmodule