module fake_netlist_1_6311_n_21 (n_1, n_2, n_4, n_3, n_0, n_21);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_21;
wire n_20;
wire n_5;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_7;
INVx1_ASAP7_75t_L g5 ( .A(n_4), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
CKINVDCx5p33_ASAP7_75t_R g7 ( .A(n_2), .Y(n_7) );
INVx2_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
INVx4_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
NOR3xp33_ASAP7_75t_SL g10 ( .A(n_7), .B(n_0), .C(n_1), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
OR2x2_ASAP7_75t_L g12 ( .A(n_11), .B(n_8), .Y(n_12) );
AND2x4_ASAP7_75t_SL g13 ( .A(n_10), .B(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_13), .B(n_9), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_14), .B(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_15), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
endmodule