module fake_jpeg_22581_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_0),
.B(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_8),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_26),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_11),
.B1(n_20),
.B2(n_16),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_29),
.A2(n_38),
.B1(n_7),
.B2(n_40),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_12),
.B1(n_13),
.B2(n_20),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_5),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_6),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_21),
.B(n_27),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_29),
.C(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_41),
.B(n_39),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_55),
.B(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_62),
.Y(n_64)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_42),
.B(n_44),
.C(n_46),
.D(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_46),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_59),
.C(n_48),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_64),
.C(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_70),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_50),
.Y(n_73)
);


endmodule