module real_aes_1451_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_783, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_783;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_0), .B(n_115), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_1), .A2(n_124), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_2), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_3), .B(n_115), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_4), .B(n_131), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_5), .B(n_131), .Y(n_194) );
INVx1_ASAP7_75t_L g122 ( .A(n_6), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_7), .B(n_131), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g759 ( .A(n_8), .Y(n_759) );
NAND2xp33_ASAP7_75t_L g132 ( .A(n_9), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g456 ( .A(n_10), .B(n_141), .Y(n_456) );
AND2x2_ASAP7_75t_L g516 ( .A(n_11), .B(n_110), .Y(n_516) );
INVx2_ASAP7_75t_L g112 ( .A(n_12), .Y(n_112) );
AOI221x1_ASAP7_75t_L g210 ( .A1(n_13), .A2(n_24), .B1(n_115), .B2(n_124), .C(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_14), .B(n_131), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_15), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_16), .B(n_115), .Y(n_114) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_17), .A2(n_110), .B(n_113), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_18), .B(n_149), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_19), .B(n_131), .Y(n_158) );
AO21x1_ASAP7_75t_L g189 ( .A1(n_20), .A2(n_115), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_21), .B(n_115), .Y(n_521) );
INVx1_ASAP7_75t_L g432 ( .A(n_22), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_23), .A2(n_86), .B1(n_115), .B2(n_461), .Y(n_460) );
NAND2x1_ASAP7_75t_L g180 ( .A(n_25), .B(n_131), .Y(n_180) );
NAND2x1_ASAP7_75t_L g168 ( .A(n_26), .B(n_133), .Y(n_168) );
OA21x2_ASAP7_75t_L g111 ( .A1(n_27), .A2(n_83), .B(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g136 ( .A(n_27), .B(n_83), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_28), .B(n_133), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_29), .B(n_131), .Y(n_130) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_30), .A2(n_141), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_31), .B(n_133), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_32), .A2(n_124), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_33), .B(n_131), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_34), .A2(n_124), .B(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g121 ( .A(n_35), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g125 ( .A(n_35), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g469 ( .A(n_35), .Y(n_469) );
OR2x6_ASAP7_75t_L g430 ( .A(n_36), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_37), .B(n_115), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_38), .B(n_115), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_39), .B(n_131), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_40), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_41), .B(n_133), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_42), .B(n_115), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_43), .A2(n_124), .B(n_452), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_44), .A2(n_124), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_45), .B(n_133), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_46), .B(n_133), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_47), .B(n_115), .Y(n_487) );
INVx1_ASAP7_75t_L g118 ( .A(n_48), .Y(n_118) );
INVx1_ASAP7_75t_L g128 ( .A(n_48), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_49), .B(n_131), .Y(n_454) );
AND2x2_ASAP7_75t_L g476 ( .A(n_50), .B(n_149), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_51), .B(n_133), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_52), .B(n_131), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_53), .B(n_133), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_54), .A2(n_124), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_55), .B(n_115), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_56), .B(n_115), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_57), .A2(n_124), .B(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_58), .Y(n_742) );
AO21x1_ASAP7_75t_L g191 ( .A1(n_59), .A2(n_124), .B(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g527 ( .A(n_60), .B(n_150), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_61), .B(n_115), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_62), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_63), .B(n_133), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_64), .B(n_115), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_65), .B(n_133), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_66), .A2(n_90), .B1(n_124), .B2(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g204 ( .A(n_67), .B(n_150), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_68), .B(n_131), .Y(n_524) );
INVx1_ASAP7_75t_L g120 ( .A(n_69), .Y(n_120) );
INVx1_ASAP7_75t_L g126 ( .A(n_69), .Y(n_126) );
AND2x2_ASAP7_75t_L g172 ( .A(n_70), .B(n_141), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_71), .B(n_133), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_72), .A2(n_124), .B(n_480), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_73), .A2(n_124), .B(n_444), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_74), .A2(n_124), .B(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g499 ( .A(n_75), .B(n_150), .Y(n_499) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_76), .A2(n_99), .B1(n_752), .B2(n_763), .C1(n_771), .C2(n_775), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g765 ( .A1(n_76), .A2(n_434), .B1(n_435), .B2(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_76), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_77), .B(n_149), .Y(n_458) );
INVx1_ASAP7_75t_L g433 ( .A(n_78), .Y(n_433) );
AND2x2_ASAP7_75t_L g140 ( .A(n_79), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_80), .B(n_115), .Y(n_160) );
AND2x2_ASAP7_75t_L g447 ( .A(n_81), .B(n_110), .Y(n_447) );
AND2x2_ASAP7_75t_L g190 ( .A(n_82), .B(n_135), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_84), .B(n_133), .Y(n_159) );
AND2x2_ASAP7_75t_L g184 ( .A(n_85), .B(n_141), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_87), .B(n_131), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_88), .A2(n_124), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_89), .B(n_133), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_91), .A2(n_124), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_92), .B(n_131), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_93), .B(n_131), .Y(n_147) );
BUFx2_ASAP7_75t_L g526 ( .A(n_94), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_95), .Y(n_748) );
BUFx2_ASAP7_75t_L g760 ( .A(n_96), .Y(n_760) );
BUFx2_ASAP7_75t_SL g779 ( .A(n_96), .Y(n_779) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_97), .A2(n_124), .B(n_129), .Y(n_123) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_742), .B(n_743), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_425), .B1(n_434), .B2(n_738), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_103), .A2(n_435), .B1(n_745), .B2(n_746), .Y(n_744) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_346), .Y(n_103) );
NOR3xp33_ASAP7_75t_SL g104 ( .A(n_105), .B(n_258), .C(n_298), .Y(n_104) );
OAI221xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_173), .B1(n_222), .B2(n_237), .C(n_240), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_137), .Y(n_107) );
INVx2_ASAP7_75t_L g255 ( .A(n_108), .Y(n_255) );
AND2x2_ASAP7_75t_L g285 ( .A(n_108), .B(n_286), .Y(n_285) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g223 ( .A(n_109), .B(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g230 ( .A(n_109), .B(n_163), .Y(n_230) );
INVx2_ASAP7_75t_L g236 ( .A(n_109), .Y(n_236) );
AND2x2_ASAP7_75t_L g245 ( .A(n_109), .B(n_139), .Y(n_245) );
INVx1_ASAP7_75t_L g261 ( .A(n_109), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_109), .B(n_307), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_110), .A2(n_521), .B(n_522), .Y(n_520) );
BUFx4f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx3_ASAP7_75t_L g142 ( .A(n_111), .Y(n_142) );
AND2x4_ASAP7_75t_L g135 ( .A(n_112), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_112), .B(n_136), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_123), .B(n_135), .Y(n_113) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_121), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
AND2x6_ASAP7_75t_L g133 ( .A(n_117), .B(n_126), .Y(n_133) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g131 ( .A(n_119), .B(n_128), .Y(n_131) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx5_ASAP7_75t_L g134 ( .A(n_121), .Y(n_134) );
AND2x2_ASAP7_75t_L g127 ( .A(n_122), .B(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_122), .Y(n_464) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
BUFx3_ASAP7_75t_L g465 ( .A(n_125), .Y(n_465) );
INVx2_ASAP7_75t_L g471 ( .A(n_126), .Y(n_471) );
AND2x4_ASAP7_75t_L g467 ( .A(n_127), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g463 ( .A(n_128), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_132), .B(n_134), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_133), .B(n_526), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_134), .A2(n_147), .B(n_148), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_134), .A2(n_158), .B(n_159), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_134), .A2(n_168), .B(n_169), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_134), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_134), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_134), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_134), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_134), .A2(n_445), .B(n_446), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_134), .A2(n_453), .B(n_454), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_134), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_134), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_134), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_134), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_134), .A2(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_SL g154 ( .A(n_135), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_135), .B(n_196), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_135), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_135), .A2(n_487), .B(n_488), .Y(n_486) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_151), .Y(n_137) );
INVx4_ASAP7_75t_L g226 ( .A(n_138), .Y(n_226) );
AND2x2_ASAP7_75t_L g257 ( .A(n_138), .B(n_164), .Y(n_257) );
AND2x2_ASAP7_75t_L g333 ( .A(n_138), .B(n_307), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g375 ( .A(n_138), .B(n_163), .Y(n_375) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_139), .B(n_163), .Y(n_262) );
AND2x2_ASAP7_75t_L g286 ( .A(n_139), .B(n_164), .Y(n_286) );
BUFx2_ASAP7_75t_L g302 ( .A(n_139), .Y(n_302) );
NOR2x1_ASAP7_75t_SL g405 ( .A(n_139), .B(n_307), .Y(n_405) );
OR2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_143), .Y(n_139) );
INVx3_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_142), .A2(n_450), .B(n_456), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_149), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_149), .Y(n_171) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_149), .A2(n_210), .B(n_214), .Y(n_209) );
OA21x2_ASAP7_75t_L g272 ( .A1(n_149), .A2(n_210), .B(n_214), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_149), .A2(n_442), .B(n_443), .Y(n_441) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_149), .A2(n_460), .B(n_466), .Y(n_459) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g282 ( .A(n_151), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_151), .A2(n_349), .B1(n_351), .B2(n_353), .C(n_358), .Y(n_348) );
AND2x2_ASAP7_75t_L g368 ( .A(n_151), .B(n_261), .Y(n_368) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_163), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g224 ( .A(n_153), .Y(n_224) );
INVx1_ASAP7_75t_L g277 ( .A(n_153), .Y(n_277) );
AO21x2_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_161), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_154), .B(n_162), .Y(n_161) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_154), .A2(n_155), .B(n_161), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_160), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_163), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g246 ( .A(n_163), .B(n_234), .Y(n_246) );
INVx2_ASAP7_75t_L g288 ( .A(n_163), .Y(n_288) );
AND2x2_ASAP7_75t_L g421 ( .A(n_163), .B(n_236), .Y(n_421) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_164), .Y(n_278) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_171), .B(n_172), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_166), .B(n_170), .Y(n_165) );
AOI21x1_ASAP7_75t_L g509 ( .A1(n_171), .A2(n_510), .B(n_516), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_205), .C(n_220), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_185), .Y(n_174) );
INVx2_ASAP7_75t_L g335 ( .A(n_175), .Y(n_335) );
AND2x2_ASAP7_75t_L g380 ( .A(n_175), .B(n_257), .Y(n_380) );
BUFx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g325 ( .A(n_176), .Y(n_325) );
AND2x4_ASAP7_75t_SL g340 ( .A(n_176), .B(n_252), .Y(n_340) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_183), .B(n_184), .Y(n_176) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_177), .A2(n_183), .B(n_184), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_182), .Y(n_177) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_183), .A2(n_198), .B(n_204), .Y(n_197) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_183), .A2(n_198), .B(n_204), .Y(n_217) );
AO21x1_ASAP7_75t_SL g492 ( .A1(n_183), .A2(n_493), .B(n_499), .Y(n_492) );
AO21x2_ASAP7_75t_L g550 ( .A1(n_183), .A2(n_493), .B(n_499), .Y(n_550) );
INVx2_ASAP7_75t_L g294 ( .A(n_185), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_185), .B(n_324), .Y(n_350) );
AND2x4_ASAP7_75t_L g383 ( .A(n_185), .B(n_330), .Y(n_383) );
AND2x4_ASAP7_75t_L g185 ( .A(n_186), .B(n_197), .Y(n_185) );
AND2x2_ASAP7_75t_L g221 ( .A(n_186), .B(n_216), .Y(n_221) );
OR2x2_ASAP7_75t_L g251 ( .A(n_186), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_SL g320 ( .A(n_186), .B(n_272), .Y(n_320) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx2_ASAP7_75t_L g265 ( .A(n_187), .Y(n_265) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g239 ( .A(n_188), .Y(n_239) );
OAI21x1_ASAP7_75t_SL g188 ( .A1(n_189), .A2(n_191), .B(n_195), .Y(n_188) );
INVx1_ASAP7_75t_L g196 ( .A(n_190), .Y(n_196) );
INVx2_ASAP7_75t_L g252 ( .A(n_197), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_199), .B(n_203), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_205), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_215), .Y(n_206) );
AND2x2_ASAP7_75t_L g220 ( .A(n_207), .B(n_221), .Y(n_220) );
OR2x2_ASAP7_75t_L g293 ( .A(n_207), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g378 ( .A(n_207), .Y(n_378) );
BUFx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x4_ASAP7_75t_L g238 ( .A(n_208), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g357 ( .A(n_208), .B(n_217), .Y(n_357) );
AND2x2_ASAP7_75t_L g361 ( .A(n_208), .B(n_227), .Y(n_361) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g330 ( .A(n_209), .Y(n_330) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_209), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_215), .B(n_238), .Y(n_314) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_218), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_216), .B(n_239), .Y(n_424) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g228 ( .A(n_217), .B(n_219), .Y(n_228) );
AND2x2_ASAP7_75t_L g310 ( .A(n_217), .B(n_272), .Y(n_310) );
AND2x2_ASAP7_75t_L g329 ( .A(n_217), .B(n_218), .Y(n_329) );
BUFx2_ASAP7_75t_L g250 ( .A(n_218), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_218), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
BUFx3_ASAP7_75t_L g227 ( .A(n_219), .Y(n_227) );
INVxp67_ASAP7_75t_L g270 ( .A(n_219), .Y(n_270) );
INVx1_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
AND2x2_ASAP7_75t_L g279 ( .A(n_221), .B(n_250), .Y(n_279) );
NAND2xp33_ASAP7_75t_L g360 ( .A(n_221), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g397 ( .A(n_221), .B(n_398), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_225), .B1(n_228), .B2(n_229), .C(n_231), .Y(n_222) );
AND2x2_ASAP7_75t_L g326 ( .A(n_223), .B(n_226), .Y(n_326) );
AND2x2_ASAP7_75t_SL g345 ( .A(n_223), .B(n_286), .Y(n_345) );
AND2x2_ASAP7_75t_L g363 ( .A(n_223), .B(n_288), .Y(n_363) );
AND2x2_ASAP7_75t_L g418 ( .A(n_223), .B(n_257), .Y(n_418) );
INVx1_ASAP7_75t_L g234 ( .A(n_224), .Y(n_234) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_224), .Y(n_290) );
CKINVDCx16_ASAP7_75t_R g370 ( .A(n_225), .Y(n_370) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_226), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_226), .B(n_277), .Y(n_352) );
AND2x2_ASAP7_75t_L g319 ( .A(n_227), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g355 ( .A(n_227), .Y(n_355) );
AND2x2_ASAP7_75t_L g264 ( .A(n_228), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_228), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g406 ( .A(n_228), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_228), .B(n_330), .Y(n_416) );
AND2x4_ASAP7_75t_L g332 ( .A(n_229), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g403 ( .A(n_230), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
OR2x2_ASAP7_75t_L g274 ( .A(n_235), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g281 ( .A(n_236), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g312 ( .A(n_236), .B(n_286), .Y(n_312) );
AND2x2_ASAP7_75t_L g386 ( .A(n_236), .B(n_307), .Y(n_386) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g334 ( .A(n_238), .B(n_335), .Y(n_334) );
OAI32xp33_ASAP7_75t_L g399 ( .A1(n_238), .A2(n_400), .A3(n_402), .B1(n_403), .B2(n_406), .Y(n_399) );
AND2x4_ASAP7_75t_L g271 ( .A(n_239), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g369 ( .A(n_239), .B(n_272), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_244), .B1(n_247), .B2(n_253), .Y(n_240) );
INVxp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g358 ( .A1(n_242), .A2(n_256), .B(n_359), .C(n_360), .Y(n_358) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g342 ( .A(n_243), .B(n_270), .Y(n_342) );
INVx1_ASAP7_75t_SL g413 ( .A(n_244), .Y(n_413) );
AND2x4_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
AND2x4_ASAP7_75t_L g316 ( .A(n_246), .B(n_255), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_246), .A2(n_395), .B1(n_396), .B2(n_397), .C(n_399), .Y(n_394) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_251), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI22xp33_ASAP7_75t_L g336 ( .A1(n_254), .A2(n_284), .B1(n_337), .B2(n_338), .Y(n_336) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
OAI211xp5_ASAP7_75t_SL g372 ( .A1(n_255), .A2(n_373), .B(n_381), .C(n_394), .Y(n_372) );
INVx2_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g292 ( .A(n_257), .B(n_261), .Y(n_292) );
OAI211xp5_ASAP7_75t_SL g258 ( .A1(n_259), .A2(n_263), .B(n_266), .C(n_295), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g289 ( .A(n_261), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g409 ( .A(n_261), .B(n_405), .Y(n_409) );
OAI32xp33_ASAP7_75t_L g366 ( .A1(n_262), .A2(n_367), .A3(n_369), .B1(n_370), .B2(n_371), .Y(n_366) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_265), .B(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_273), .B1(n_279), .B2(n_280), .C(n_283), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g423 ( .A(n_270), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_271), .B(n_335), .Y(n_337) );
A2O1A1O1Ixp25_ASAP7_75t_L g408 ( .A1(n_271), .A2(n_340), .B(n_356), .C(n_402), .D(n_409), .Y(n_408) );
AOI31xp33_ASAP7_75t_L g410 ( .A1(n_271), .A2(n_292), .A3(n_402), .B(n_409), .Y(n_410) );
AND2x2_ASAP7_75t_L g324 ( .A(n_272), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_274), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx2_ASAP7_75t_L g401 ( .A(n_276), .Y(n_401) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g396 ( .A(n_277), .B(n_288), .Y(n_396) );
INVx1_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
AND2x2_ASAP7_75t_L g296 ( .A(n_280), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AOI31xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .A3(n_291), .B(n_293), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_286), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g419 ( .A(n_286), .B(n_365), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AND2x2_ASAP7_75t_L g364 ( .A(n_288), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g390 ( .A(n_288), .Y(n_390) );
INVxp67_ASAP7_75t_L g359 ( .A(n_289), .Y(n_359) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g297 ( .A(n_293), .Y(n_297) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND3xp33_ASAP7_75t_SL g298 ( .A(n_299), .B(n_315), .C(n_331), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_308), .B1(n_312), .B2(n_313), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g385 ( .A(n_302), .Y(n_385) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_306), .Y(n_365) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_306), .Y(n_391) );
OR2x2_ASAP7_75t_L g392 ( .A(n_306), .B(n_375), .Y(n_392) );
NAND2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g343 ( .A(n_310), .Y(n_343) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_326), .B2(n_327), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_318), .B(n_321), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_324), .A2(n_329), .B1(n_363), .B2(n_364), .C(n_366), .Y(n_362) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2x1_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g402 ( .A(n_329), .Y(n_402) );
AND2x2_ASAP7_75t_L g339 ( .A(n_330), .B(n_340), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_SL g387 ( .A1(n_330), .A2(n_388), .B(n_392), .C(n_393), .Y(n_387) );
AOI211xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_336), .C(n_341), .Y(n_331) );
AND2x2_ASAP7_75t_L g382 ( .A(n_335), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g393 ( .A(n_340), .Y(n_393) );
AOI21xp33_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_343), .B(n_344), .Y(n_341) );
INVx2_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NOR3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_372), .C(n_407), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_348), .B(n_362), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g371 ( .A(n_356), .Y(n_371) );
INVxp67_ASAP7_75t_L g395 ( .A(n_360), .Y(n_395) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g379 ( .A(n_369), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B1(n_379), .B2(n_380), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_387), .Y(n_381) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g420 ( .A(n_405), .B(n_421), .Y(n_420) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B1(n_411), .B2(n_414), .C(n_417), .Y(n_407) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI31xp33_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_419), .A3(n_420), .B(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx4f_ASAP7_75t_SL g745 ( .A(n_425), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
CKINVDCx11_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
OR2x6_ASAP7_75t_SL g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AND2x6_ASAP7_75t_SL g741 ( .A(n_428), .B(n_430), .Y(n_741) );
OR2x2_ASAP7_75t_L g751 ( .A(n_428), .B(n_430), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_428), .B(n_429), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx3_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_SL g435 ( .A(n_436), .B(n_634), .Y(n_435) );
NOR3xp33_ASAP7_75t_SL g436 ( .A(n_437), .B(n_543), .C(n_575), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_472), .B1(n_500), .B2(n_517), .C(n_528), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_448), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g506 ( .A(n_440), .B(n_449), .Y(n_506) );
INVx4_ASAP7_75t_L g534 ( .A(n_440), .Y(n_534) );
AND2x4_ASAP7_75t_SL g574 ( .A(n_440), .B(n_508), .Y(n_574) );
BUFx2_ASAP7_75t_L g584 ( .A(n_440), .Y(n_584) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_440), .B(n_589), .Y(n_650) );
AND2x2_ASAP7_75t_L g659 ( .A(n_440), .B(n_587), .Y(n_659) );
OR2x2_ASAP7_75t_L g667 ( .A(n_440), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g693 ( .A(n_440), .B(n_532), .Y(n_693) );
AND2x4_ASAP7_75t_L g712 ( .A(n_440), .B(n_713), .Y(n_712) );
OR2x6_ASAP7_75t_L g440 ( .A(n_441), .B(n_447), .Y(n_440) );
INVx2_ASAP7_75t_SL g625 ( .A(n_448), .Y(n_625) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_457), .Y(n_448) );
AND2x2_ASAP7_75t_L g532 ( .A(n_449), .B(n_509), .Y(n_532) );
INVx2_ASAP7_75t_L g559 ( .A(n_449), .Y(n_559) );
INVx2_ASAP7_75t_L g589 ( .A(n_449), .Y(n_589) );
AND2x2_ASAP7_75t_L g603 ( .A(n_449), .B(n_508), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_455), .Y(n_450) );
AND2x2_ASAP7_75t_L g533 ( .A(n_457), .B(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g556 ( .A(n_457), .Y(n_556) );
BUFx3_ASAP7_75t_L g570 ( .A(n_457), .Y(n_570) );
AND2x2_ASAP7_75t_L g599 ( .A(n_457), .B(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
AND2x4_ASAP7_75t_L g504 ( .A(n_458), .B(n_459), .Y(n_504) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_465), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
NOR2x1p5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g605 ( .A(n_472), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_483), .Y(n_472) );
OR2x2_ASAP7_75t_L g716 ( .A(n_473), .B(n_517), .Y(n_716) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g572 ( .A(n_474), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_474), .B(n_483), .Y(n_633) );
OR2x2_ASAP7_75t_L g731 ( .A(n_474), .B(n_653), .Y(n_731) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g542 ( .A(n_475), .B(n_518), .Y(n_542) );
OR2x2_ASAP7_75t_SL g552 ( .A(n_475), .B(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g563 ( .A(n_475), .Y(n_563) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_475), .Y(n_614) );
NAND2x1_ASAP7_75t_L g620 ( .A(n_475), .B(n_519), .Y(n_620) );
AND2x2_ASAP7_75t_L g645 ( .A(n_475), .B(n_485), .Y(n_645) );
OR2x2_ASAP7_75t_L g666 ( .A(n_475), .B(n_549), .Y(n_666) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g561 ( .A(n_483), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_483), .A2(n_655), .B(n_658), .C(n_660), .Y(n_654) );
AND2x2_ASAP7_75t_L g727 ( .A(n_483), .B(n_503), .Y(n_727) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_492), .Y(n_483) );
INVx1_ASAP7_75t_L g594 ( .A(n_484), .Y(n_594) );
AND2x2_ASAP7_75t_L g664 ( .A(n_484), .B(n_519), .Y(n_664) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g538 ( .A(n_485), .Y(n_538) );
OR2x2_ASAP7_75t_L g553 ( .A(n_485), .B(n_519), .Y(n_553) );
INVx1_ASAP7_75t_L g569 ( .A(n_485), .Y(n_569) );
AND2x2_ASAP7_75t_L g581 ( .A(n_485), .B(n_492), .Y(n_581) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_485), .Y(n_687) );
NOR2x1_ASAP7_75t_SL g518 ( .A(n_492), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
INVxp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .Y(n_501) );
OR2x2_ASAP7_75t_L g651 ( .A(n_502), .B(n_586), .Y(n_651) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_503), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g733 ( .A(n_503), .B(n_630), .Y(n_733) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g578 ( .A(n_504), .B(n_559), .Y(n_578) );
AND2x2_ASAP7_75t_L g674 ( .A(n_504), .B(n_587), .Y(n_674) );
INVx1_ASAP7_75t_L g591 ( .A(n_505), .Y(n_591) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g641 ( .A(n_506), .Y(n_641) );
INVx2_ASAP7_75t_L g608 ( .A(n_507), .Y(n_608) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g558 ( .A(n_508), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g588 ( .A(n_508), .Y(n_588) );
INVx1_ASAP7_75t_L g713 ( .A(n_508), .Y(n_713) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_509), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
OR2x2_ASAP7_75t_L g684 ( .A(n_517), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_SL g539 ( .A(n_519), .Y(n_539) );
OR2x2_ASAP7_75t_L g562 ( .A(n_519), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g573 ( .A(n_519), .B(n_549), .Y(n_573) );
AND2x2_ASAP7_75t_L g647 ( .A(n_519), .B(n_563), .Y(n_647) );
BUFx2_ASAP7_75t_L g730 ( .A(n_519), .Y(n_730) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_527), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_535), .B(n_540), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g682 ( .A(n_531), .B(n_604), .Y(n_682) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g541 ( .A(n_532), .B(n_534), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_533), .B(n_603), .Y(n_704) );
INVx1_ASAP7_75t_L g734 ( .A(n_533), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_534), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_534), .B(n_670), .Y(n_707) );
INVxp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
AND2x4_ASAP7_75t_SL g571 ( .A(n_537), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_537), .B(n_565), .Y(n_718) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_538), .B(n_620), .Y(n_676) );
AND2x2_ASAP7_75t_L g694 ( .A(n_538), .B(n_647), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_539), .B(n_581), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_539), .A2(n_585), .B(n_627), .C(n_632), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_539), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_541), .A2(n_614), .B1(n_722), .B2(n_728), .C(n_732), .Y(n_721) );
INVx1_ASAP7_75t_SL g709 ( .A(n_542), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_554), .B1(n_560), .B2(n_564), .C(n_783), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_551), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g619 ( .A(n_548), .Y(n_619) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g593 ( .A(n_549), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g624 ( .A(n_549), .B(n_569), .Y(n_624) );
INVx2_ASAP7_75t_L g657 ( .A(n_549), .Y(n_657) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OAI32xp33_ASAP7_75t_L g708 ( .A1(n_552), .A2(n_599), .A3(n_630), .B1(n_709), .B2(n_710), .Y(n_708) );
OR2x2_ASAP7_75t_L g679 ( .A(n_553), .B(n_666), .Y(n_679) );
INVx1_ASAP7_75t_L g689 ( .A(n_554), .Y(n_689) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
INVx2_ASAP7_75t_L g604 ( .A(n_555), .Y(n_604) );
AND2x2_ASAP7_75t_L g675 ( .A(n_555), .B(n_650), .Y(n_675) );
OR2x2_ASAP7_75t_L g706 ( .A(n_555), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_556), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g600 ( .A(n_559), .Y(n_600) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx2_ASAP7_75t_SL g565 ( .A(n_562), .Y(n_565) );
OR2x2_ASAP7_75t_L g652 ( .A(n_562), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_563), .B(n_581), .Y(n_580) );
NOR2xp67_ASAP7_75t_L g686 ( .A(n_563), .B(n_687), .Y(n_686) );
BUFx2_ASAP7_75t_L g699 ( .A(n_563), .Y(n_699) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B(n_571), .C(n_574), .Y(n_564) );
AND2x2_ASAP7_75t_L g714 ( .A(n_566), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
BUFx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g640 ( .A(n_570), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_570), .B(n_574), .Y(n_661) );
AND2x2_ASAP7_75t_L g692 ( .A(n_570), .B(n_693), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_572), .A2(n_703), .B(n_705), .C(n_708), .Y(n_702) );
AOI222xp33_ASAP7_75t_L g576 ( .A1(n_573), .A2(n_577), .B1(n_579), .B2(n_582), .C1(n_590), .C2(n_592), .Y(n_576) );
AND2x2_ASAP7_75t_L g644 ( .A(n_573), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g577 ( .A(n_574), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g598 ( .A(n_574), .Y(n_598) );
NAND4xp25_ASAP7_75t_L g575 ( .A(n_576), .B(n_595), .C(n_616), .D(n_626), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_578), .B(n_584), .Y(n_638) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g646 ( .A(n_581), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_SL g653 ( .A(n_581), .Y(n_653) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_583), .A2(n_617), .B(n_621), .C(n_625), .Y(n_616) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_584), .B(n_599), .Y(n_720) );
OR2x2_ASAP7_75t_L g724 ( .A(n_584), .B(n_610), .Y(n_724) );
INVx1_ASAP7_75t_L g697 ( .A(n_585), .Y(n_697) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_SL g631 ( .A(n_588), .Y(n_631) );
INVx1_ASAP7_75t_L g611 ( .A(n_589), .Y(n_611) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_591), .B(n_628), .Y(n_627) );
BUFx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g615 ( .A(n_593), .Y(n_615) );
AOI322xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .A3(n_599), .B1(n_601), .B2(n_605), .C1(n_606), .C2(n_612), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_SL g677 ( .A1(n_598), .A2(n_678), .B(n_679), .C(n_680), .Y(n_677) );
INVx1_ASAP7_75t_L g700 ( .A(n_599), .Y(n_700) );
NOR2xp67_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g658 ( .A(n_604), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_610), .Y(n_680) );
INVx2_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx3_ASAP7_75t_L g623 ( .A(n_620), .Y(n_623) );
OR2x2_ASAP7_75t_L g691 ( .A(n_620), .B(n_653), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_620), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_SL g723 ( .A(n_624), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_625), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND3xp33_ASAP7_75t_SL g728 ( .A(n_633), .B(n_729), .C(n_731), .Y(n_728) );
NOR3xp33_ASAP7_75t_SL g634 ( .A(n_635), .B(n_672), .C(n_701), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_636), .B(n_654), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_639), .B(n_642), .C(n_648), .Y(n_636) );
OAI31xp33_ASAP7_75t_L g681 ( .A1(n_637), .A2(n_659), .A3(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx2_ASAP7_75t_L g696 ( .A(n_644), .Y(n_696) );
INVx1_ASAP7_75t_L g671 ( .A(n_646), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B(n_652), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g698 ( .A(n_656), .B(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g737 ( .A(n_657), .Y(n_737) );
OAI22xp33_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_662), .B1(n_667), .B2(n_671), .Y(n_660) );
INVx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_666), .Y(n_678) );
OR2x2_ASAP7_75t_L g729 ( .A(n_666), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g672 ( .A(n_673), .B(n_681), .C(n_688), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B(n_676), .C(n_677), .Y(n_673) );
INVx2_ASAP7_75t_L g710 ( .A(n_674), .Y(n_710) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_692), .B2(n_694), .C(n_695), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_698), .B2(n_700), .Y(n_695) );
NAND3xp33_ASAP7_75t_SL g701 ( .A(n_702), .B(n_711), .C(n_721), .Y(n_701) );
INVxp33_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B1(n_717), .B2(n_719), .Y(n_711) );
INVx2_ASAP7_75t_L g725 ( .A(n_712), .Y(n_725) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp33_ASAP7_75t_SL g732 ( .A1(n_731), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx6p67_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx4_ASAP7_75t_SL g746 ( .A(n_739), .Y(n_746) );
INVx3_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g743 ( .A1(n_742), .A2(n_744), .B(n_747), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_761), .Y(n_754) );
INVxp67_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_757), .B(n_760), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OR2x2_ASAP7_75t_SL g774 ( .A(n_758), .B(n_760), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g776 ( .A1(n_758), .A2(n_777), .B(n_780), .Y(n_776) );
INVx1_ASAP7_75t_SL g768 ( .A(n_761), .Y(n_768) );
NOR2xp33_ASAP7_75t_SL g769 ( .A(n_761), .B(n_770), .Y(n_769) );
BUFx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
BUFx2_ASAP7_75t_L g781 ( .A(n_762), .Y(n_781) );
INVxp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_767), .B(n_769), .Y(n_764) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
CKINVDCx9p33_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
CKINVDCx11_ASAP7_75t_R g777 ( .A(n_778), .Y(n_777) );
CKINVDCx8_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
endmodule