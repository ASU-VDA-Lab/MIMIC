module fake_jpeg_5639_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_0),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_23),
.B1(n_17),
.B2(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_25),
.Y(n_64)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_15),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_40),
.B1(n_36),
.B2(n_35),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_61),
.B1(n_65),
.B2(n_68),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_36),
.B1(n_35),
.B2(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_36),
.B1(n_26),
.B2(n_23),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_18),
.B1(n_17),
.B2(n_28),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_11),
.B1(n_14),
.B2(n_4),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_20),
.B1(n_19),
.B2(n_18),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_75),
.Y(n_96)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_37),
.B1(n_32),
.B2(n_8),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_22),
.C(n_21),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_82),
.C(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_83),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_42),
.A2(n_22),
.B(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_91),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_76),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_1),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_83),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_76),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_109),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_120),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_61),
.C(n_80),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_118),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_99),
.B1(n_90),
.B2(n_84),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_81),
.B(n_32),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_122),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_72),
.C(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_2),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_37),
.B(n_3),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_135),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_115),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_137),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_101),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_136),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_140),
.Y(n_152)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_121),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_113),
.B(n_118),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_114),
.B1(n_131),
.B2(n_111),
.Y(n_156)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_117),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g153 ( 
.A(n_142),
.B(n_124),
.C(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_156),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_146),
.C(n_139),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_129),
.B1(n_95),
.B2(n_132),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_138),
.B1(n_145),
.B2(n_84),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_111),
.B1(n_131),
.B2(n_95),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_104),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_160),
.B(n_163),
.Y(n_170)
);

FAx1_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_147),
.CI(n_140),
.CON(n_160),
.SN(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_148),
.C(n_143),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_164),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_152),
.B(n_89),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_122),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_160),
.B(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_98),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_92),
.C(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_158),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_170),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_153),
.B1(n_158),
.B2(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_176),
.A2(n_171),
.B(n_173),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_175),
.C(n_103),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_12),
.Y(n_179)
);


endmodule