module fake_ibex_1010_n_649 (n_85, n_84, n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_649);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_649;

wire n_151;
wire n_599;
wire n_507;
wire n_540;
wire n_395;
wire n_171;
wire n_103;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_108;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_255;
wire n_175;
wire n_586;
wire n_638;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_94;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_645;
wire n_500;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_556;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_106;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_550;
wire n_169;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_109;
wire n_127;
wire n_121;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_122;
wire n_523;
wire n_116;
wire n_614;
wire n_370;
wire n_431;
wire n_574;
wire n_289;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_136;
wire n_261;
wire n_521;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_437;
wire n_602;
wire n_355;
wire n_474;
wire n_594;
wire n_636;
wire n_407;
wire n_102;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_623;
wire n_585;
wire n_530;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_576;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_488;
wire n_139;
wire n_514;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_98;
wire n_129;
wire n_613;
wire n_267;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_643;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_554;
wire n_553;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_365;
wire n_605;
wire n_539;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_624;
wire n_411;
wire n_135;
wire n_520;
wire n_512;
wire n_615;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_627;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_582;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_218;
wire n_314;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_633;
wire n_532;
wire n_95;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_118;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_639;
wire n_303;
wire n_362;
wire n_93;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_501;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_311;
wire n_406;
wire n_606;
wire n_97;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_631;
wire n_260;
wire n_620;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_159;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_14),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_22),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_61),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g108 ( 
.A(n_74),
.Y(n_108)
);

INVxp33_ASAP7_75t_SL g109 ( 
.A(n_36),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_16),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_38),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_39),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_2),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_11),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_15),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_25),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_17),
.B(n_3),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_0),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_2),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_65),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_19),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_20),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_54),
.Y(n_148)
);

NOR2xp67_ASAP7_75t_L g149 ( 
.A(n_41),
.B(n_29),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_75),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_82),
.Y(n_151)
);

INVxp33_ASAP7_75t_SL g152 ( 
.A(n_45),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_12),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_42),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_33),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_53),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_32),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_43),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_52),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_55),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_48),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_59),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_1),
.Y(n_168)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_111),
.B(n_1),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

BUFx8_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

NAND2x1p5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_46),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_3),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_97),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_4),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_100),
.B(n_5),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g184 ( 
.A(n_121),
.B(n_63),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_100),
.B(n_7),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_9),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_97),
.B(n_9),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_96),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_133),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_106),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_106),
.B(n_148),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_129),
.B(n_24),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_137),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_95),
.B(n_30),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_139),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_140),
.B(n_31),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_127),
.B(n_34),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_35),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_192),
.Y(n_234)
);

NAND2xp33_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_143),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_200),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_201),
.B(n_109),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_198),
.B(n_162),
.Y(n_241)
);

AO221x1_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_150),
.B1(n_126),
.B2(n_158),
.C(n_157),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_160),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_152),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_152),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_151),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_L g248 ( 
.A(n_184),
.B(n_173),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

AOI221xp5_ASAP7_75t_L g250 ( 
.A1(n_169),
.A2(n_126),
.B1(n_136),
.B2(n_150),
.C(n_122),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_159),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_203),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_172),
.B(n_124),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_187),
.A2(n_93),
.B1(n_107),
.B2(n_108),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_180),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_156),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_168),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_200),
.B(n_155),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_168),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_173),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_180),
.Y(n_262)
);

BUFx8_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_200),
.B(n_149),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_37),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_40),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_177),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_223),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_188),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_185),
.A2(n_79),
.B1(n_80),
.B2(n_84),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_214),
.B(n_233),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_191),
.B(n_91),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_181),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_214),
.B(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_193),
.Y(n_276)
);

NOR2x1p5_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_174),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_193),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_179),
.B(n_189),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_185),
.A2(n_183),
.B1(n_169),
.B2(n_210),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_230),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_181),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_194),
.B(n_208),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_194),
.B(n_208),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_195),
.B(n_209),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_218),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_195),
.B(n_209),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_197),
.B(n_231),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g291 ( 
.A(n_210),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_176),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_L g293 ( 
.A(n_184),
.B(n_229),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_197),
.B(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_178),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_199),
.B(n_220),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_190),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_190),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_199),
.B(n_212),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_207),
.B(n_224),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_213),
.B(n_219),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_213),
.B(n_219),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_223),
.B(n_227),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_184),
.Y(n_304)
);

OR2x2_ASAP7_75t_SL g305 ( 
.A(n_251),
.B(n_205),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_258),
.A2(n_227),
.B1(n_218),
.B2(n_184),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_246),
.B(n_225),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_260),
.A2(n_186),
.B1(n_170),
.B2(n_175),
.Y(n_308)
);

OR2x6_ASAP7_75t_SL g309 ( 
.A(n_251),
.B(n_167),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_279),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_238),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_167),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_182),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_244),
.B(n_217),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_267),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_281),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_245),
.B(n_182),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_272),
.B(n_275),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_261),
.B(n_186),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_240),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_253),
.B(n_234),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_239),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_283),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_236),
.B(n_269),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_263),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_255),
.Y(n_333)
);

BUFx8_ASAP7_75t_L g334 ( 
.A(n_291),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_280),
.B(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_254),
.B(n_257),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_241),
.B(n_243),
.Y(n_338)
);

OR2x6_ASAP7_75t_L g339 ( 
.A(n_264),
.B(n_259),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_241),
.B(n_243),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_259),
.B(n_300),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

AND2x6_ASAP7_75t_L g346 ( 
.A(n_270),
.B(n_276),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_252),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_292),
.Y(n_349)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_302),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_293),
.A2(n_278),
.B1(n_289),
.B2(n_290),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_294),
.A2(n_296),
.B1(n_298),
.B2(n_297),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_271),
.A2(n_235),
.B1(n_266),
.B2(n_265),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_249),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_256),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_262),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_274),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_304),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_282),
.A2(n_247),
.B1(n_242),
.B2(n_226),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_303),
.B(n_216),
.Y(n_363)
);

AND3x1_ASAP7_75t_SL g364 ( 
.A(n_250),
.B(n_277),
.C(n_171),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_238),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_248),
.B(n_293),
.C(n_303),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_238),
.Y(n_367)
);

AND3x1_ASAP7_75t_SL g368 ( 
.A(n_250),
.B(n_277),
.C(n_171),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_291),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_303),
.B(n_216),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_303),
.B(n_216),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_303),
.B(n_216),
.Y(n_372)
);

NAND3xp33_ASAP7_75t_SL g373 ( 
.A(n_247),
.B(n_250),
.C(n_232),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_237),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_238),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_238),
.Y(n_376)
);

CKINVDCx6p67_ASAP7_75t_R g377 ( 
.A(n_309),
.Y(n_377)
);

INVx3_ASAP7_75t_SL g378 ( 
.A(n_369),
.Y(n_378)
);

BUFx12f_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

AOI222xp33_ASAP7_75t_L g380 ( 
.A1(n_311),
.A2(n_373),
.B1(n_318),
.B2(n_328),
.C1(n_372),
.C2(n_371),
.Y(n_380)
);

BUFx12f_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_341),
.B(n_345),
.Y(n_382)
);

O2A1O1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_363),
.A2(n_370),
.B(n_333),
.C(n_322),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_341),
.A2(n_364),
.B1(n_368),
.B2(n_337),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_330),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_332),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_317),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_312),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_344),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_337),
.A2(n_339),
.B1(n_335),
.B2(n_307),
.Y(n_393)
);

O2A1O1Ixp33_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_325),
.B(n_314),
.C(n_315),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_326),
.B(n_339),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_313),
.B(n_376),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_339),
.B(n_375),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_319),
.B(n_365),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_321),
.B(n_367),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_331),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

INVx8_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_355),
.A2(n_352),
.B1(n_354),
.B2(n_327),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_374),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_310),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_324),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_316),
.Y(n_411)
);

OR2x6_ASAP7_75t_L g412 ( 
.A(n_305),
.B(n_323),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_308),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_346),
.B(n_306),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_346),
.B(n_348),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_356),
.Y(n_416)
);

OAI21xp33_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_357),
.B(n_358),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_360),
.A2(n_356),
.B(n_359),
.C(n_350),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_350),
.A2(n_341),
.B1(n_311),
.B2(n_345),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_311),
.B(n_345),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_341),
.B(n_311),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_341),
.B(n_311),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_309),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

NAND2x2_ASAP7_75t_L g428 ( 
.A(n_334),
.B(n_277),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_338),
.A2(n_293),
.B(n_340),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

NAND3xp33_ASAP7_75t_L g432 ( 
.A(n_362),
.B(n_250),
.C(n_280),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_351),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_318),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_341),
.A2(n_311),
.B1(n_345),
.B2(n_340),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_338),
.A2(n_293),
.B(n_340),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_311),
.B(n_345),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_366),
.A2(n_307),
.B(n_320),
.C(n_322),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_345),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_345),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_341),
.A2(n_311),
.B1(n_345),
.B2(n_340),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_317),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_311),
.A2(n_351),
.B1(n_345),
.B2(n_312),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_362),
.B(n_250),
.C(n_280),
.Y(n_444)
);

BUFx2_ASAP7_75t_SL g445 ( 
.A(n_330),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_317),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_351),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_421),
.Y(n_448)
);

NOR2x1_ASAP7_75t_R g449 ( 
.A(n_379),
.B(n_381),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_426),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_424),
.Y(n_451)
);

BUFx4f_ASAP7_75t_SL g452 ( 
.A(n_377),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_391),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_435),
.A2(n_441),
.B1(n_382),
.B2(n_398),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_431),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_387),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_397),
.B(n_392),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_395),
.B(n_393),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

BUFx8_ASAP7_75t_SL g465 ( 
.A(n_434),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_420),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_403),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_438),
.A2(n_430),
.B(n_436),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_378),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_383),
.B(n_384),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_407),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_409),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_380),
.B(n_443),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_406),
.A2(n_394),
.B(n_414),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_404),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_427),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_402),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_429),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_411),
.B(n_432),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_442),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_446),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_447),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_444),
.B(n_412),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_433),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

AO32x1_ASAP7_75t_L g498 ( 
.A1(n_413),
.A2(n_416),
.A3(n_418),
.B1(n_417),
.B2(n_412),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_415),
.A2(n_428),
.B(n_425),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_437),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_379),
.B(n_381),
.Y(n_501)
);

AO21x1_ASAP7_75t_SL g502 ( 
.A1(n_389),
.A2(n_401),
.B(n_400),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_437),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_437),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_379),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_437),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_437),
.B(n_421),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_408),
.A2(n_394),
.B(n_415),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_421),
.B(n_437),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_426),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_437),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_511),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_453),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_455),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_453),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_456),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_459),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_460),
.B(n_462),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_476),
.B(n_448),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_472),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_511),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_458),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_465),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_465),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_468),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_463),
.B(n_454),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_469),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_504),
.B(n_488),
.Y(n_530)
);

NOR4xp25_ASAP7_75t_SL g531 ( 
.A(n_505),
.B(n_470),
.C(n_489),
.D(n_480),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_488),
.A2(n_494),
.B1(n_463),
.B2(n_503),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_474),
.B(n_500),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_494),
.A2(n_463),
.B1(n_471),
.B2(n_496),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_477),
.B(n_512),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_475),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_473),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_475),
.B(n_506),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_467),
.B(n_487),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_464),
.B(n_490),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_497),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_497),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_482),
.B(n_478),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_524),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_517),
.Y(n_545)
);

NAND4xp25_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_501),
.C(n_492),
.D(n_491),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_524),
.Y(n_547)
);

NAND4xp25_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_485),
.C(n_483),
.D(n_479),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_540),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_517),
.A2(n_452),
.B1(n_478),
.B2(n_470),
.Y(n_550)
);

AOI221xp5_ASAP7_75t_L g551 ( 
.A1(n_515),
.A2(n_466),
.B1(n_461),
.B2(n_505),
.C(n_508),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_517),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_516),
.B(n_484),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_514),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_522),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_517),
.Y(n_556)
);

AOI33xp33_ASAP7_75t_L g557 ( 
.A1(n_519),
.A2(n_449),
.A3(n_452),
.B1(n_499),
.B2(n_493),
.B3(n_484),
.Y(n_557)
);

NAND3xp33_ASAP7_75t_SL g558 ( 
.A(n_531),
.B(n_478),
.C(n_486),
.Y(n_558)
);

NOR2x1_ASAP7_75t_L g559 ( 
.A(n_517),
.B(n_481),
.Y(n_559)
);

INVx3_ASAP7_75t_SL g560 ( 
.A(n_517),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_521),
.A2(n_482),
.B1(n_499),
.B2(n_486),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_528),
.B(n_482),
.Y(n_562)
);

AOI211x1_ASAP7_75t_L g563 ( 
.A1(n_530),
.A2(n_498),
.B(n_481),
.C(n_482),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_516),
.B(n_493),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_450),
.Y(n_565)
);

NAND4xp25_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_495),
.C(n_457),
.D(n_510),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_514),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_519),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_518),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_513),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_527),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_562),
.B(n_535),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_535),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_544),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_547),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_571),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_560),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_569),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_572),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_549),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_560),
.Y(n_582)
);

OAI32xp33_ASAP7_75t_L g583 ( 
.A1(n_546),
.A2(n_538),
.A3(n_542),
.B1(n_541),
.B2(n_537),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_568),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_567),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_555),
.B(n_520),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_553),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_539),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_548),
.B(n_525),
.Y(n_589)
);

AOI21xp33_ASAP7_75t_SL g590 ( 
.A1(n_589),
.A2(n_550),
.B(n_526),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_574),
.B(n_529),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_582),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_585),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_581),
.B(n_557),
.Y(n_594)
);

OR2x6_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_552),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_584),
.B(n_557),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_576),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_565),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_576),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_578),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_598),
.B(n_573),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_600),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_592),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_592),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_597),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_599),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_594),
.B(n_575),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_596),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_593),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_593),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_595),
.A2(n_583),
.B(n_579),
.Y(n_611)
);

NOR3x1_ASAP7_75t_L g612 ( 
.A(n_607),
.B(n_558),
.C(n_566),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_608),
.B(n_591),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_607),
.B(n_577),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_605),
.Y(n_615)
);

AOI211xp5_ASAP7_75t_L g616 ( 
.A1(n_604),
.A2(n_590),
.B(n_583),
.C(n_603),
.Y(n_616)
);

NAND4xp75_ASAP7_75t_L g617 ( 
.A(n_611),
.B(n_563),
.C(n_559),
.D(n_586),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_602),
.B(n_545),
.Y(n_618)
);

AOI211xp5_ASAP7_75t_L g619 ( 
.A1(n_601),
.A2(n_551),
.B(n_552),
.C(n_570),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_609),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_615),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_613),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_616),
.B(n_561),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_613),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_614),
.B(n_606),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_620),
.B(n_591),
.Y(n_626)
);

AOI311xp33_ASAP7_75t_L g627 ( 
.A1(n_619),
.A2(n_580),
.A3(n_588),
.B(n_610),
.C(n_587),
.Y(n_627)
);

NAND2x1_ASAP7_75t_SL g628 ( 
.A(n_612),
.B(n_556),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_618),
.Y(n_629)
);

XOR2x1_ASAP7_75t_L g630 ( 
.A(n_627),
.B(n_531),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_624),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_623),
.B(n_545),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_628),
.B(n_617),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_625),
.Y(n_634)
);

NAND2x1p5_ASAP7_75t_L g635 ( 
.A(n_629),
.B(n_570),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_631),
.Y(n_636)
);

AND2x2_ASAP7_75t_SL g637 ( 
.A(n_633),
.B(n_630),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_634),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_633),
.A2(n_623),
.B(n_621),
.Y(n_639)
);

NOR2x1p5_ASAP7_75t_L g640 ( 
.A(n_636),
.B(n_622),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_638),
.B(n_639),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_638),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_637),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_641),
.Y(n_644)
);

OR3x1_ASAP7_75t_L g645 ( 
.A(n_640),
.B(n_632),
.C(n_635),
.Y(n_645)
);

AOI221xp5_ASAP7_75t_SL g646 ( 
.A1(n_641),
.A2(n_626),
.B1(n_543),
.B2(n_536),
.C(n_539),
.Y(n_646)
);

OAI32xp33_ASAP7_75t_L g647 ( 
.A1(n_643),
.A2(n_644),
.A3(n_645),
.B1(n_646),
.B2(n_523),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_647),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_648),
.A2(n_533),
.B(n_543),
.Y(n_649)
);


endmodule