module real_jpeg_18674_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_0),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_0),
.Y(n_138)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_0),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_1),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_2),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_2),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_2),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_2),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_2),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_2),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_2),
.B(n_330),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_3),
.Y(n_126)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_3),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_4),
.Y(n_200)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_5),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_5),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_5),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_6),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_6),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_7),
.B(n_27),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_7),
.B(n_65),
.Y(n_64)
);

AND2x4_ASAP7_75t_SL g83 ( 
.A(n_7),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_7),
.B(n_113),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g158 ( 
.A(n_7),
.B(n_159),
.Y(n_158)
);

AND2x4_ASAP7_75t_SL g256 ( 
.A(n_7),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_7),
.B(n_316),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_8),
.A2(n_13),
.B1(n_39),
.B2(n_42),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_8),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_8),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_8),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_8),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_8),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_8),
.B(n_69),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_8),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_8),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_9),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_9),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_9),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_9),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_9),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_9),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_9),
.B(n_365),
.Y(n_364)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_11),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_11),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_11),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_11),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_11),
.B(n_126),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_13),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_13),
.B(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_13),
.Y(n_248)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_14),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_14),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_58),
.Y(n_57)
);

AND2x4_ASAP7_75t_SL g88 ( 
.A(n_15),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_15),
.B(n_110),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_15),
.B(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_15),
.B(n_213),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_16),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_223),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_221),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_172),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_20),
.B(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_100),
.C(n_139),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_22),
.A2(n_23),
.B1(n_100),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_60),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_24),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.C(n_47),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_25),
.B(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_29),
.C(n_33),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_32),
.Y(n_314)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_34),
.Y(n_351)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_37),
.A2(n_38),
.B1(n_47),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_38),
.A2(n_240),
.B(n_247),
.Y(n_239)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_41),
.Y(n_310)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_45),
.Y(n_282)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_47),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.C(n_57),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_48),
.A2(n_49),
.B1(n_57),
.B2(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_48),
.A2(n_49),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_54),
.B(n_144),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_73),
.B1(n_98),
.B2(n_99),
.Y(n_60)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_62),
.B(n_182),
.C(n_183),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_64),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_64),
.B(n_255),
.C(n_260),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_64),
.A2(n_183),
.B1(n_260),
.B2(n_261),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_67),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_68),
.Y(n_182)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_87),
.C(n_92),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_74),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_83),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_75),
.A2(n_83),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_75),
.Y(n_238)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_79),
.B(n_236),
.Y(n_235)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_83),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_83),
.B(n_297),
.Y(n_296)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_100),
.Y(n_229)
);

XNOR2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_128),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_102),
.B(n_116),
.C(n_128),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_111),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_103),
.A2(n_111),
.B1(n_112),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_111),
.B(n_280),
.C(n_283),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_111),
.A2(n_112),
.B1(n_280),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_114),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_117),
.B(n_125),
.C(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_125),
.A2(n_127),
.B1(n_199),
.B2(n_204),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_131),
.C(n_135),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_134),
.Y(n_263)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_140),
.B(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_165),
.C(n_169),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_141),
.B(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.C(n_151),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_143),
.B(n_289),
.Y(n_288)
);

XNOR2x1_ASAP7_75t_L g289 ( 
.A(n_146),
.B(n_151),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_147),
.B(n_150),
.Y(n_287)
);

NOR2x1_ASAP7_75t_R g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_158),
.C(n_162),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_152),
.B(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_157),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_158),
.A2(n_162),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_158),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_158),
.B(n_339),
.C(n_341),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_158),
.A2(n_277),
.B1(n_341),
.B2(n_342),
.Y(n_354)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_160),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_161),
.Y(n_360)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_162),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_169),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.C(n_176),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_194),
.B1(n_219),
.B2(n_220),
.Y(n_177)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_194),
.Y(n_220)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_290),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.C(n_267),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_227),
.B(n_231),
.Y(n_393)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.C(n_264),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_264),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.C(n_254),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_239),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_237),
.B(n_298),
.C(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_255),
.B(n_381),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g328 ( 
.A(n_256),
.B(n_259),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_256),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_256),
.A2(n_348),
.B1(n_349),
.B2(n_362),
.Y(n_361)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_268),
.B(n_270),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.C(n_288),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_271),
.B(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_273),
.B(n_288),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.C(n_286),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_274),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_279),
.B(n_287),
.Y(n_376)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_323),
.Y(n_322)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_392),
.C(n_393),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_387),
.B(n_391),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_372),
.B(n_386),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_333),
.B(n_371),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_319),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_295),
.B(n_319),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_303),
.C(n_311),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_303),
.A2(n_304),
.B1(n_311),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_305),
.B(n_309),
.Y(n_340)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_311),
.Y(n_337)
);

AO22x1_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_315),
.B1(n_317),
.B2(n_318),
.Y(n_311)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_315),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_317),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_318),
.B(n_364),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_325),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_321),
.B(n_325),
.C(n_385),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_322),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_326),
.B(n_328),
.C(n_329),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_345),
.B(n_370),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_SL g370 ( 
.A(n_335),
.B(n_338),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_339),
.A2(n_340),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_355),
.B(n_369),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_352),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_352),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_349),
.Y(n_362)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_363),
.B(n_368),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_361),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_361),
.Y(n_368)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_384),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_SL g386 ( 
.A(n_373),
.B(n_384),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_377),
.B2(n_378),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_379),
.C(n_383),
.Y(n_388)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_388),
.B(n_389),
.Y(n_391)
);


endmodule