module real_jpeg_3868_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_0),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_0),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_0),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_0),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_0),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_0),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_0),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_1),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_1),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_1),
.B(n_190),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_1),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_1),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_1),
.B(n_393),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_1),
.B(n_108),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_2),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_2),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_2),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_3),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_3),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_3),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_3),
.B(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_4),
.Y(n_174)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_4),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_5),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_5),
.B(n_64),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_5),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_5),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_5),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_5),
.B(n_116),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_5),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_5),
.B(n_416),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_6),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_7),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_7),
.B(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_7),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_7),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_7),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_7),
.B(n_190),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_7),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_7),
.B(n_192),
.Y(n_417)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_9),
.Y(n_540)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_10),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_10),
.Y(n_300)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_12),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_12),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_12),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_12),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_12),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_12),
.B(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_13),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_13),
.Y(n_332)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_15),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_15),
.B(n_146),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_15),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_15),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_15),
.B(n_71),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_15),
.B(n_396),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_15),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_16),
.B(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_16),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_16),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_16),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_16),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_16),
.B(n_187),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_16),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_16),
.B(n_377),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_17),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_17),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_17),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_17),
.B(n_176),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_17),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_17),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_17),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_18),
.B(n_44),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_18),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_18),
.B(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_18),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_18),
.B(n_28),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_18),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_18),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_18),
.B(n_424),
.Y(n_423)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_538),
.B(n_541),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_40),
.B(n_78),
.C(n_537),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_24),
.B(n_48),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.C(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_26),
.A2(n_31),
.B1(n_39),
.B2(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_31),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_52),
.C(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_33),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_34),
.B(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_74),
.C(n_76),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_63),
.C(n_67),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_50),
.B(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_52),
.A2(n_57),
.B1(n_70),
.B2(n_118),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_54),
.Y(n_160)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_55),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_68),
.C(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_63),
.B(n_67),
.Y(n_125)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_66),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_68),
.A2(n_69),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_70),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_70),
.A2(n_111),
.B1(n_112),
.B2(n_118),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_73),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_73),
.Y(n_344)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_73),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_129),
.B(n_536),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_126),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_80),
.B(n_126),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_123),
.C(n_124),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_81),
.A2(n_82),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_106),
.C(n_119),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_83),
.A2(n_84),
.B1(n_512),
.B2(n_514),
.Y(n_511)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_94),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_90),
.C(n_94),
.Y(n_123)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_93),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.C(n_101),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_95),
.B(n_502),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_502)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_105),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_106),
.A2(n_119),
.B1(n_120),
.B2(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_106),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_118),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_107),
.B(n_508),
.Y(n_507)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_111),
.A2(n_112),
.B1(n_206),
.B2(n_211),
.Y(n_205)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_112),
.B(n_201),
.C(n_206),
.Y(n_509)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_117),
.Y(n_294)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_117),
.Y(n_340)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_123),
.B(n_124),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_530),
.B(n_535),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_495),
.B(n_527),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_302),
.B(n_494),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_257),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_133),
.B(n_257),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_198),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_134),
.B(n_199),
.C(n_236),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_171),
.C(n_180),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_135),
.B(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_147),
.C(n_161),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_136),
.B(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_140),
.C(n_143),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_142),
.B(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_146),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_147),
.A2(n_148),
.B1(n_161),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_157),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_149),
.B(n_157),
.Y(n_470)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_152),
.B(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_156),
.Y(n_223)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_156),
.Y(n_419)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_160),
.Y(n_362)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_161),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_162),
.B(n_164),
.C(n_168),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_167),
.B1(n_168),
.B2(n_170),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_166),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_166),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_167),
.B(n_206),
.C(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_167),
.A2(n_168),
.B1(n_206),
.B2(n_211),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_171),
.B(n_180),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_175),
.B(n_177),
.C(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_178),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_178),
.B(n_241),
.C(n_250),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.C(n_195),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_181),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_189),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_182),
.B(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_186),
.B(n_189),
.Y(n_269)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_191),
.B(n_195),
.Y(n_286)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_193),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_194),
.Y(n_219)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_236),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_212),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_200),
.B(n_213),
.C(n_224),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_210),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_224),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.C(n_220),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_220),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_224),
.Y(n_544)
);

FAx1_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.CI(n_235),
.CON(n_224),
.SN(n_224)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_225),
.B(n_231),
.C(n_235),
.Y(n_510)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_229),
.Y(n_416)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_230),
.Y(n_397)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_234),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_251),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_238),
.B(n_240),
.C(n_251),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.C(n_255),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_255),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.C(n_264),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_259),
.B(n_262),
.Y(n_490)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_264),
.B(n_490),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_284),
.C(n_287),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_266),
.B(n_483),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.C(n_277),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_267),
.A2(n_268),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_270),
.A2(n_271),
.B(n_273),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_270),
.B(n_277),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.C(n_282),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_438)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_282),
.B(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_283),
.B(n_374),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_287),
.Y(n_484)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_298),
.C(n_301),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_289),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.C(n_295),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_290),
.B(n_450),
.Y(n_449)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_293),
.A2(n_295),
.B1(n_296),
.B2(n_451),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_293),
.Y(n_451)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_298),
.B(n_301),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_488),
.B(n_493),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_475),
.B(n_487),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_457),
.B(n_474),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_431),
.B(n_456),
.Y(n_305)
);

AOI21x1_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_401),
.B(n_430),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_366),
.B(n_400),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_346),
.B(n_365),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_323),
.B(n_345),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_320),
.B(n_322),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_318),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_315),
.Y(n_324)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_325),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_336),
.B2(n_337),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_339),
.C(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_333),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_333),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_364),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_364),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_356),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_355),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_355),
.C(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_354),
.Y(n_371)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_356),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_384),
.C(n_385),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_363),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_363),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_369),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_382),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_383),
.C(n_386),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_373),
.C(n_375),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_378),
.B1(n_379),
.B2(n_381),
.Y(n_375)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_376),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_381),
.Y(n_411)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_SL g425 ( 
.A(n_380),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_395),
.C(n_398),
.Y(n_428)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_392),
.A2(n_395),
.B1(n_398),
.B2(n_399),
.Y(n_391)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_392),
.Y(n_398)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_394),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_395),
.Y(n_399)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_429),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_429),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_413),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_412),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_404),
.B(n_412),
.C(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_411),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_410),
.Y(n_405)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_410),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_411),
.B(n_445),
.C(n_446),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_413),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_420),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_422),
.C(n_427),
.Y(n_434)
);

BUFx24_ASAP7_75t_SL g546 ( 
.A(n_414),
.Y(n_546)
);

FAx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_417),
.CI(n_418),
.CON(n_414),
.SN(n_414)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_415),
.B(n_417),
.C(n_418),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_422),
.B1(n_427),
.B2(n_428),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_426),
.Y(n_441)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_454),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_454),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_443),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_435),
.C(n_443),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_439),
.B2(n_440),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_466),
.C(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_448),
.C(n_453),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_449),
.B1(n_452),
.B2(n_453),
.Y(n_447)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_448),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_449),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_473),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_473),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_459),
.B(n_464),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_463),
.C(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_461),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_468),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_469),
.C(n_471),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_485),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_485),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_477),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_482),
.C(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_491),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_491),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_523),
.Y(n_495)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_496),
.A2(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_516),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_516),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_499),
.B1(n_505),
.B2(n_515),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_498),
.B(n_506),
.C(n_511),
.Y(n_534)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.C(n_503),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_518),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_501),
.A2(n_503),
.B1(n_504),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_501),
.Y(n_519)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_505),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_511),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_509),
.C(n_510),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_521),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_510),
.Y(n_521)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_512),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.C(n_522),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_520),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_525),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_524),
.B(n_526),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_524),
.B(n_526),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_534),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_534),
.Y(n_535)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_532),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx13_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_540),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_543),
.Y(n_541)
);


endmodule