module fake_ibex_524_n_842 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_158, n_132, n_157, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_842);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_158;
input n_132;
input n_157;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_842;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_747;
wire n_500;
wire n_645;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_798;
wire n_732;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_281;
wire n_758;
wire n_636;
wire n_594;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_385;
wire n_342;
wire n_233;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g159 ( 
.A(n_42),
.Y(n_159)
);

NOR2xp67_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_6),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_71),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_75),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_156),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_2),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_68),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_66),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_108),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_27),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_57),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_35),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_31),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_139),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_26),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_114),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_55),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_13),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_15),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_3),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_4),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_125),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_32),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_6),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_51),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_89),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_97),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_80),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_5),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_54),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_95),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_103),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_45),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_33),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_24),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_63),
.Y(n_212)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_33),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_39),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_119),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_23),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_76),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_133),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_84),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_32),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_79),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_19),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_106),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_81),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_72),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_48),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_35),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_43),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_91),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_41),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_142),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_121),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_17),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_112),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_46),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_117),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_9),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_11),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_102),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_144),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_38),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_14),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_69),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_85),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_132),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_29),
.B(n_110),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_70),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_21),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_49),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_23),
.Y(n_255)
);

OAI22x1_ASAP7_75t_R g256 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

AND2x6_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_36),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_170),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_179),
.B(n_0),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_163),
.B(n_1),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_169),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g268 ( 
.A1(n_200),
.A2(n_77),
.B(n_154),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g269 ( 
.A(n_194),
.B(n_37),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_170),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_7),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_175),
.B(n_8),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_198),
.A2(n_231),
.B1(n_209),
.B2(n_212),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_167),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_175),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_183),
.B(n_9),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_170),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_222),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_177),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_177),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_172),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_173),
.Y(n_286)
);

BUFx8_ASAP7_75t_L g287 ( 
.A(n_170),
.Y(n_287)
);

OA21x2_ASAP7_75t_L g288 ( 
.A1(n_200),
.A2(n_82),
.B(n_153),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_190),
.B(n_10),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_220),
.B(n_12),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_187),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_170),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_170),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_210),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_207),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_164),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_219),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_225),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_238),
.B(n_16),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_206),
.A2(n_228),
.B1(n_241),
.B2(n_212),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_243),
.B(n_16),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_224),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_190),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_207),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_217),
.Y(n_307)
);

AND2x6_ASAP7_75t_L g308 ( 
.A(n_216),
.B(n_40),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_217),
.A2(n_87),
.B(n_150),
.Y(n_309)
);

BUFx8_ASAP7_75t_L g310 ( 
.A(n_159),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_216),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_218),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_255),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_206),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_232),
.B(n_25),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_218),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_245),
.B(n_25),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_232),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_166),
.B(n_27),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_189),
.B(n_28),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_195),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_209),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_180),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_304),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_289),
.B(n_182),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_304),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_273),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_263),
.B(n_188),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_289),
.B(n_184),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_263),
.B(n_192),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_265),
.B(n_201),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_258),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_259),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_287),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_262),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_258),
.A2(n_234),
.B1(n_214),
.B2(n_215),
.Y(n_346)
);

BUFx4f_ASAP7_75t_L g347 ( 
.A(n_275),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_271),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_271),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_323),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_L g354 ( 
.A(n_258),
.B(n_161),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_257),
.B(n_193),
.Y(n_355)
);

AOI22x1_ASAP7_75t_L g356 ( 
.A1(n_279),
.A2(n_230),
.B1(n_202),
.B2(n_197),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_279),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_323),
.B(n_203),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_258),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_275),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_287),
.B(n_264),
.C(n_278),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_296),
.Y(n_363)
);

BUFx6f_ASAP7_75t_SL g364 ( 
.A(n_299),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_306),
.Y(n_365)
);

OR2x6_ASAP7_75t_L g366 ( 
.A(n_314),
.B(n_160),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_286),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_286),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_258),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_262),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_L g373 ( 
.A1(n_315),
.A2(n_324),
.B1(n_267),
.B2(n_274),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_306),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_294),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_297),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_307),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_285),
.B(n_196),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_305),
.Y(n_379)
);

INVx8_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_269),
.B(n_199),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_259),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_266),
.B(n_204),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_292),
.B(n_205),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_301),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_L g387 ( 
.A(n_308),
.B(n_162),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_310),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_291),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_308),
.B(n_208),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_272),
.B(n_221),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_312),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_298),
.B(n_185),
.Y(n_398)
);

AOI21x1_ASAP7_75t_L g399 ( 
.A1(n_309),
.A2(n_229),
.B(n_233),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_310),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_320),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_270),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_268),
.A2(n_240),
.B(n_248),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_270),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_270),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_311),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_283),
.B(n_252),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_284),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_318),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_270),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_283),
.B(n_213),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_L g414 ( 
.A1(n_295),
.A2(n_255),
.B1(n_223),
.B2(n_253),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_L g415 ( 
.A(n_321),
.B(n_254),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_276),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_318),
.B(n_237),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_319),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_336),
.A2(n_303),
.B1(n_300),
.B2(n_282),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_351),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_340),
.B(n_165),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

O2A1O1Ixp5_ASAP7_75t_L g425 ( 
.A1(n_405),
.A2(n_337),
.B(n_327),
.C(n_399),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_340),
.B(n_174),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_347),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_332),
.A2(n_228),
.B1(n_241),
.B2(n_242),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_374),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_383),
.B(n_393),
.Y(n_433)
);

AND3x1_ASAP7_75t_L g434 ( 
.A(n_335),
.B(n_256),
.C(n_251),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_377),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_370),
.B(n_178),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_333),
.A2(n_403),
.B1(n_336),
.B2(n_346),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_378),
.A2(n_239),
.B(n_249),
.C(n_250),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_346),
.A2(n_236),
.B1(n_186),
.B2(n_191),
.Y(n_441)
);

AND3x1_ASAP7_75t_L g442 ( 
.A(n_335),
.B(n_30),
.C(n_34),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_338),
.B(n_227),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_380),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_348),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_352),
.B(n_171),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_354),
.A2(n_288),
.B(n_268),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_339),
.B(n_235),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_327),
.B(n_181),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_347),
.Y(n_452)
);

AOI21x1_ASAP7_75t_L g453 ( 
.A1(n_337),
.A2(n_268),
.B(n_288),
.Y(n_453)
);

BUFx5_ASAP7_75t_L g454 ( 
.A(n_392),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_362),
.B(n_244),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_359),
.B(n_288),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_355),
.B(n_284),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_394),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_390),
.B(n_413),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_413),
.B(n_276),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_364),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_397),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_364),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_373),
.A2(n_302),
.B1(n_290),
.B2(n_281),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_367),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_369),
.B(n_378),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_384),
.B(n_280),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_343),
.B(n_280),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_415),
.B(n_280),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_381),
.B(n_280),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_387),
.B(n_290),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_392),
.B(n_302),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_356),
.Y(n_476)
);

OR2x2_ASAP7_75t_SL g477 ( 
.A(n_376),
.B(n_44),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_330),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_361),
.B(n_47),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_366),
.B(n_50),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_330),
.B(n_52),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_388),
.B(n_53),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_373),
.B(n_331),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_331),
.A2(n_56),
.B(n_58),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_334),
.B(n_60),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_366),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_334),
.B(n_65),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_326),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_410),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_421),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_447),
.B(n_414),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_447),
.B(n_414),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_439),
.A2(n_366),
.B1(n_386),
.B2(n_328),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_424),
.B(n_401),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_449),
.A2(n_341),
.B(n_375),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_425),
.A2(n_341),
.B(n_375),
.Y(n_499)
);

NOR3xp33_ASAP7_75t_L g500 ( 
.A(n_429),
.B(n_371),
.C(n_344),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_430),
.B(n_349),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_439),
.A2(n_372),
.B1(n_358),
.B2(n_357),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_420),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_425),
.A2(n_368),
.B(n_350),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_456),
.A2(n_372),
.B(n_350),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_430),
.B(n_358),
.Y(n_509)
);

O2A1O1Ixp33_ASAP7_75t_L g510 ( 
.A1(n_483),
.A2(n_368),
.B(n_329),
.C(n_379),
.Y(n_510)
);

NAND2x1_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_385),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_436),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_453),
.A2(n_402),
.B(n_391),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_418),
.A2(n_400),
.B(n_402),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_462),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_428),
.B(n_452),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_478),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_419),
.B(n_410),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_419),
.B(n_433),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_459),
.B(n_410),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_433),
.B(n_410),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_438),
.B(n_448),
.Y(n_522)
);

CKINVDCx8_ASAP7_75t_R g523 ( 
.A(n_480),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_432),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_436),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_468),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_465),
.A2(n_404),
.B1(n_412),
.B2(n_407),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_476),
.A2(n_406),
.B(n_416),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_451),
.B(n_440),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_L g531 ( 
.A(n_455),
.B(n_73),
.C(n_74),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_446),
.Y(n_532)
);

AO32x1_ASAP7_75t_L g533 ( 
.A1(n_486),
.A2(n_382),
.A3(n_342),
.B1(n_86),
.B2(n_90),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_477),
.A2(n_444),
.B1(n_458),
.B2(n_466),
.Y(n_534)
);

O2A1O1Ixp33_ASAP7_75t_L g535 ( 
.A1(n_460),
.A2(n_78),
.B(n_83),
.C(n_92),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_462),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_464),
.B(n_93),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_463),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_480),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_422),
.A2(n_94),
.B(n_96),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_443),
.B(n_155),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_436),
.B(n_98),
.Y(n_544)
);

OA22x2_ASAP7_75t_L g545 ( 
.A1(n_480),
.A2(n_149),
.B1(n_104),
.B2(n_109),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_464),
.B(n_113),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_473),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_427),
.A2(n_124),
.B(n_126),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_436),
.B(n_127),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_450),
.B(n_128),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_467),
.B(n_129),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_434),
.B(n_148),
.Y(n_552)
);

AOI221xp5_ASAP7_75t_L g553 ( 
.A1(n_442),
.A2(n_130),
.B1(n_137),
.B2(n_138),
.C(n_140),
.Y(n_553)
);

CKINVDCx10_ASAP7_75t_R g554 ( 
.A(n_482),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_441),
.B(n_479),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_490),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_457),
.B(n_491),
.Y(n_557)
);

BUFx4f_ASAP7_75t_L g558 ( 
.A(n_491),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_469),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_470),
.B(n_145),
.Y(n_560)
);

INVx3_ASAP7_75t_SL g561 ( 
.A(n_437),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_474),
.A2(n_475),
.B(n_472),
.Y(n_563)
);

NOR3xp33_ASAP7_75t_L g564 ( 
.A(n_481),
.B(n_487),
.C(n_485),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_L g565 ( 
.A(n_481),
.B(n_485),
.C(n_484),
.Y(n_565)
);

BUFx8_ASAP7_75t_L g566 ( 
.A(n_454),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_445),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_496),
.B(n_454),
.Y(n_568)
);

O2A1O1Ixp5_ASAP7_75t_SL g569 ( 
.A1(n_534),
.A2(n_549),
.B(n_544),
.C(n_547),
.Y(n_569)
);

OA21x2_ASAP7_75t_L g570 ( 
.A1(n_529),
.A2(n_454),
.B(n_498),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_499),
.A2(n_506),
.B(n_527),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_508),
.A2(n_563),
.B(n_530),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_545),
.A2(n_546),
.B(n_543),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_522),
.A2(n_519),
.B1(n_523),
.B2(n_555),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_494),
.B(n_503),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_509),
.B(n_504),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_505),
.B(n_507),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_492),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_524),
.B(n_539),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_526),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_501),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_495),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_517),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_552),
.A2(n_559),
.B1(n_546),
.B2(n_553),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_515),
.B(n_500),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_497),
.B(n_516),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_516),
.B(n_561),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_566),
.Y(n_589)
);

AOI221xp5_ASAP7_75t_SL g590 ( 
.A1(n_518),
.A2(n_510),
.B1(n_535),
.B2(n_542),
.C(n_548),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_520),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_521),
.A2(n_557),
.B(n_514),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_567),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_538),
.B(n_558),
.Y(n_594)
);

O2A1O1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_531),
.A2(n_550),
.B(n_551),
.C(n_562),
.Y(n_595)
);

AO31x2_ASAP7_75t_L g596 ( 
.A1(n_533),
.A2(n_512),
.A3(n_525),
.B(n_560),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_SL g597 ( 
.A1(n_536),
.A2(n_540),
.B(n_554),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_511),
.A2(n_512),
.B(n_525),
.Y(n_598)
);

AO31x2_ASAP7_75t_L g599 ( 
.A1(n_533),
.A2(n_525),
.A3(n_566),
.B(n_537),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_492),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_R g601 ( 
.A(n_523),
.B(n_421),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_503),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_503),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_492),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_492),
.Y(n_605)
);

AO21x2_ASAP7_75t_L g606 ( 
.A1(n_565),
.A2(n_564),
.B(n_449),
.Y(n_606)
);

AO31x2_ASAP7_75t_L g607 ( 
.A1(n_498),
.A2(n_449),
.A3(n_506),
.B(n_499),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_503),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_493),
.B(n_439),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_556),
.B(n_380),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_522),
.A2(n_527),
.B(n_530),
.C(n_519),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_503),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_508),
.A2(n_425),
.B(n_499),
.Y(n_614)
);

AO32x2_ASAP7_75t_L g615 ( 
.A1(n_534),
.A2(n_502),
.A3(n_486),
.B1(n_528),
.B2(n_541),
.Y(n_615)
);

AOI221xp5_ASAP7_75t_SL g616 ( 
.A1(n_522),
.A2(n_519),
.B1(n_483),
.B2(n_530),
.C(n_440),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_496),
.B(n_386),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_493),
.B(n_439),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_493),
.B(n_439),
.Y(n_619)
);

OA21x2_ASAP7_75t_L g620 ( 
.A1(n_513),
.A2(n_449),
.B(n_405),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_493),
.B(n_439),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_493),
.B(n_439),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_493),
.B(n_439),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_566),
.Y(n_624)
);

BUFx12f_ASAP7_75t_L g625 ( 
.A(n_497),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_541),
.B(n_421),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_508),
.A2(n_425),
.B(n_499),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_496),
.B(n_386),
.Y(n_628)
);

OAI22x1_ASAP7_75t_L g629 ( 
.A1(n_541),
.A2(n_301),
.B1(n_274),
.B2(n_371),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_496),
.B(n_386),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_522),
.A2(n_519),
.B1(n_523),
.B2(n_530),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_522),
.A2(n_527),
.B(n_530),
.C(n_519),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_493),
.B(n_439),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_503),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_523),
.B(n_340),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_493),
.B(n_439),
.Y(n_636)
);

A2O1A1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_522),
.A2(n_527),
.B(n_530),
.C(n_519),
.Y(n_637)
);

BUFx12f_ASAP7_75t_L g638 ( 
.A(n_497),
.Y(n_638)
);

NAND3xp33_ASAP7_75t_L g639 ( 
.A(n_565),
.B(n_465),
.C(n_553),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_602),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_582),
.B(n_618),
.Y(n_641)
);

AOI21xp33_ASAP7_75t_SL g642 ( 
.A1(n_597),
.A2(n_574),
.B(n_631),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_574),
.A2(n_631),
.B1(n_585),
.B2(n_576),
.Y(n_643)
);

CKINVDCx11_ASAP7_75t_R g644 ( 
.A(n_625),
.Y(n_644)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_601),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_603),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_609),
.B(n_619),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_608),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_578),
.Y(n_649)
);

NAND2x1_ASAP7_75t_L g650 ( 
.A(n_573),
.B(n_584),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_633),
.B(n_621),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_622),
.A2(n_623),
.B1(n_636),
.B2(n_586),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_575),
.B(n_577),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_638),
.Y(n_655)
);

NAND3xp33_ASAP7_75t_L g656 ( 
.A(n_585),
.B(n_616),
.C(n_569),
.Y(n_656)
);

AO21x2_ASAP7_75t_L g657 ( 
.A1(n_614),
.A2(n_627),
.B(n_606),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_607),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_611),
.A2(n_595),
.B(n_592),
.Y(n_659)
);

OA21x2_ASAP7_75t_L g660 ( 
.A1(n_590),
.A2(n_639),
.B(n_616),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_613),
.Y(n_661)
);

INVx8_ASAP7_75t_L g662 ( 
.A(n_626),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_607),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_607),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_620),
.A2(n_598),
.B(n_570),
.Y(n_665)
);

AO222x2_ASAP7_75t_L g666 ( 
.A1(n_587),
.A2(n_629),
.B1(n_626),
.B2(n_597),
.C1(n_628),
.C2(n_617),
.Y(n_666)
);

INVx6_ASAP7_75t_L g667 ( 
.A(n_604),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_612),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_577),
.B(n_583),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_605),
.Y(n_670)
);

AO21x1_ASAP7_75t_L g671 ( 
.A1(n_591),
.A2(n_568),
.B(n_579),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_604),
.Y(n_672)
);

BUFx2_ASAP7_75t_SL g673 ( 
.A(n_589),
.Y(n_673)
);

OA21x2_ASAP7_75t_L g674 ( 
.A1(n_596),
.A2(n_599),
.B(n_634),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_588),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_600),
.Y(n_676)
);

AOI22x1_ASAP7_75t_L g677 ( 
.A1(n_580),
.A2(n_581),
.B1(n_593),
.B2(n_624),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_594),
.A2(n_610),
.B(n_635),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_635),
.A2(n_615),
.B(n_630),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_615),
.A2(n_639),
.B(n_527),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_599),
.B(n_615),
.Y(n_681)
);

BUFx2_ASAP7_75t_R g682 ( 
.A(n_588),
.Y(n_682)
);

AO31x2_ASAP7_75t_L g683 ( 
.A1(n_571),
.A2(n_572),
.A3(n_632),
.B(n_611),
.Y(n_683)
);

OR3x4_ASAP7_75t_SL g684 ( 
.A(n_589),
.B(n_624),
.C(n_523),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_582),
.B(n_618),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_589),
.B(n_624),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_618),
.B(n_633),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_578),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_611),
.A2(n_637),
.B(n_632),
.C(n_585),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_578),
.Y(n_690)
);

NAND2x1p5_ASAP7_75t_L g691 ( 
.A(n_604),
.B(n_492),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_607),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_602),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_618),
.B(n_633),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_604),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_582),
.B(n_618),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_602),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_695),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_658),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_672),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_SL g701 ( 
.A1(n_643),
.A2(n_695),
.B1(n_677),
.B2(n_667),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_650),
.B(n_662),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_663),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_662),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_664),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_653),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_667),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_688),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_662),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_690),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_667),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_692),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_654),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_641),
.B(n_685),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_686),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_670),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_R g718 ( 
.A1(n_666),
.A2(n_647),
.B1(n_684),
.B2(n_697),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_687),
.B(n_694),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_662),
.B(n_679),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_691),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_691),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_683),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_640),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_641),
.B(n_685),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_696),
.B(n_669),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_683),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_652),
.B(n_651),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_683),
.Y(n_729)
);

AO21x2_ASAP7_75t_L g730 ( 
.A1(n_656),
.A2(n_659),
.B(n_680),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_646),
.Y(n_731)
);

OR2x6_ASAP7_75t_L g732 ( 
.A(n_673),
.B(n_678),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_676),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_652),
.B(n_642),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_668),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_648),
.B(n_693),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_661),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_674),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_689),
.B(n_657),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_699),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_739),
.B(n_699),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_705),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_718),
.A2(n_671),
.B1(n_666),
.B2(n_675),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_739),
.B(n_657),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_703),
.B(n_674),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_713),
.B(n_681),
.Y(n_746)
);

INVx5_ASAP7_75t_L g747 ( 
.A(n_702),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_720),
.B(n_665),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_706),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_728),
.B(n_660),
.Y(n_750)
);

INVxp67_ASAP7_75t_SL g751 ( 
.A(n_714),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_723),
.B(n_727),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_718),
.A2(n_675),
.B1(n_660),
.B2(n_686),
.Y(n_753)
);

CKINVDCx14_ASAP7_75t_R g754 ( 
.A(n_716),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_740),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_741),
.B(n_738),
.Y(n_756)
);

AND2x4_ASAP7_75t_SL g757 ( 
.A(n_754),
.B(n_716),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_746),
.B(n_729),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_743),
.A2(n_734),
.B1(n_726),
.B2(n_715),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_742),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_740),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_750),
.B(n_709),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_751),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_750),
.B(n_715),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_747),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_746),
.B(n_730),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_743),
.B(n_655),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_752),
.B(n_730),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_752),
.B(n_730),
.Y(n_769)
);

NAND2x1p5_ASAP7_75t_L g770 ( 
.A(n_747),
.B(n_698),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_764),
.B(n_751),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_755),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_761),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_767),
.B(n_733),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_764),
.B(n_744),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_766),
.B(n_745),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_760),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_758),
.B(n_734),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_758),
.B(n_749),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_766),
.B(n_745),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_765),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_765),
.B(n_748),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_776),
.B(n_768),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_776),
.B(n_768),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_772),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_774),
.B(n_753),
.C(n_763),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_777),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_772),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_775),
.B(n_762),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_773),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_780),
.B(n_769),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_780),
.B(n_769),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_782),
.B(n_756),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_773),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_783),
.B(n_779),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_783),
.B(n_778),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_786),
.B(n_775),
.Y(n_797)
);

NOR4xp25_ASAP7_75t_L g798 ( 
.A(n_789),
.B(n_753),
.C(n_759),
.D(n_737),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_787),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_793),
.A2(n_754),
.B(n_781),
.Y(n_800)
);

AO22x1_ASAP7_75t_L g801 ( 
.A1(n_793),
.A2(n_781),
.B1(n_782),
.B2(n_765),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_789),
.A2(n_771),
.B1(n_782),
.B2(n_770),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_785),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_788),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_797),
.B(n_791),
.Y(n_805)
);

OAI221xp5_ASAP7_75t_L g806 ( 
.A1(n_798),
.A2(n_701),
.B1(n_784),
.B2(n_794),
.C(n_790),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_797),
.B(n_791),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_796),
.B(n_792),
.Y(n_808)
);

NAND4xp75_ASAP7_75t_L g809 ( 
.A(n_805),
.B(n_800),
.C(n_795),
.D(n_644),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_808),
.Y(n_810)
);

AOI322xp5_ASAP7_75t_L g811 ( 
.A1(n_807),
.A2(n_792),
.A3(n_717),
.B1(n_735),
.B2(n_804),
.C1(n_803),
.C2(n_799),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_811),
.B(n_802),
.Y(n_812)
);

NOR3xp33_ASAP7_75t_SL g813 ( 
.A(n_809),
.B(n_645),
.C(n_806),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_812),
.B(n_813),
.C(n_644),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_813),
.A2(n_810),
.B1(n_801),
.B2(n_799),
.Y(n_815)
);

CKINVDCx6p67_ASAP7_75t_R g816 ( 
.A(n_814),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_815),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_817),
.B(n_686),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_816),
.B(n_682),
.Y(n_819)
);

XOR2x1_ASAP7_75t_L g820 ( 
.A(n_819),
.B(n_816),
.Y(n_820)
);

OA21x2_ASAP7_75t_L g821 ( 
.A1(n_818),
.A2(n_684),
.B(n_722),
.Y(n_821)
);

XOR2x2_ASAP7_75t_L g822 ( 
.A(n_819),
.B(n_719),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_822),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_820),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_821),
.A2(n_700),
.B1(n_721),
.B2(n_707),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_821),
.A2(n_747),
.B1(n_757),
.B2(n_770),
.Y(n_826)
);

NAND4xp75_ASAP7_75t_L g827 ( 
.A(n_821),
.B(n_721),
.C(n_708),
.D(n_736),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_SL g828 ( 
.A(n_824),
.B(n_708),
.Y(n_828)
);

OAI21xp33_ASAP7_75t_L g829 ( 
.A1(n_823),
.A2(n_711),
.B(n_704),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_827),
.Y(n_830)
);

OAI21x1_ASAP7_75t_SL g831 ( 
.A1(n_825),
.A2(n_710),
.B(n_725),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_826),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_824),
.A2(n_700),
.B(n_732),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_824),
.A2(n_732),
.B(n_724),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_830),
.B(n_710),
.C(n_712),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_832),
.A2(n_747),
.B1(n_757),
.B2(n_732),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_833),
.B(n_731),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_834),
.A2(n_710),
.B1(n_732),
.B2(n_747),
.Y(n_838)
);

AOI31xp67_ASAP7_75t_SL g839 ( 
.A1(n_837),
.A2(n_828),
.A3(n_829),
.B(n_831),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_835),
.B(n_836),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_840),
.B(n_704),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_838),
.B1(n_839),
.B2(n_712),
.Y(n_842)
);


endmodule