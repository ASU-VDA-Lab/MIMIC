module fake_jpeg_7970_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx2_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx3_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_28),
.Y(n_67)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_19),
.B1(n_26),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_51),
.B1(n_57),
.B2(n_61),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_52),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

AO22x2_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_23),
.B1(n_18),
.B2(n_17),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_41),
.B1(n_34),
.B2(n_23),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_59),
.B1(n_63),
.B2(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_61),
.B1(n_41),
.B2(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_86),
.B1(n_85),
.B2(n_89),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_44),
.B(n_34),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_79),
.C(n_68),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_38),
.C(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_38),
.Y(n_82)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_41),
.B1(n_34),
.B2(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_94),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_28),
.B1(n_25),
.B2(n_32),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_89),
.B1(n_29),
.B2(n_16),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_16),
.B1(n_27),
.B2(n_25),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_32),
.B1(n_27),
.B2(n_29),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_49),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_35),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_96),
.A2(n_106),
.B1(n_112),
.B2(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_120),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_24),
.Y(n_150)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_111),
.B1(n_95),
.B2(n_87),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_115),
.B1(n_121),
.B2(n_91),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_76),
.B1(n_79),
.B2(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_48),
.B1(n_65),
.B2(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_117),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_50),
.B1(n_46),
.B2(n_33),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_35),
.C(n_43),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_22),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_90),
.B1(n_83),
.B2(n_87),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_22),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_143),
.C(n_150),
.Y(n_165)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_83),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_138),
.B(n_151),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_90),
.B1(n_81),
.B2(n_80),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_148),
.B1(n_120),
.B2(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_103),
.B(n_43),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_145),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_92),
.B(n_88),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_70),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_95),
.B1(n_88),
.B2(n_12),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_100),
.A2(n_66),
.B1(n_62),
.B2(n_21),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_62),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_96),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_0),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_97),
.Y(n_161)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_116),
.C(n_105),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_165),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_117),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_109),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_122),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_108),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_111),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_129),
.B(n_123),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_136),
.B1(n_128),
.B2(n_132),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_24),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_179),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_183),
.B1(n_184),
.B2(n_202),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_189),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_143),
.B1(n_132),
.B2(n_146),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_146),
.B1(n_128),
.B2(n_133),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_161),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_135),
.B1(n_125),
.B2(n_137),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_194),
.B1(n_205),
.B2(n_177),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_188),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_138),
.A3(n_150),
.B1(n_151),
.B2(n_130),
.C1(n_148),
.C2(n_124),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_199),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_197),
.C(n_199),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_152),
.A2(n_138),
.B1(n_150),
.B2(n_144),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_151),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_144),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_175),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_155),
.A2(n_157),
.B(n_162),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_170),
.B(n_174),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_178),
.A2(n_144),
.B1(n_24),
.B2(n_31),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_24),
.B1(n_20),
.B2(n_3),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_214),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_166),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_210),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

AO21x2_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_189),
.B(n_201),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_213),
.B1(n_219),
.B2(n_183),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_164),
.B1(n_160),
.B2(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_215),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

AO22x1_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_171),
.B1(n_157),
.B2(n_159),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_166),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_227),
.C(n_230),
.Y(n_231)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_168),
.C(n_158),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_158),
.C(n_163),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_241),
.B1(n_245),
.B2(n_209),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_204),
.C(n_184),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_237),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_248),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_179),
.C(n_156),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_220),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_251),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_173),
.B1(n_205),
.B2(n_202),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_177),
.B1(n_179),
.B2(n_182),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_222),
.B1(n_228),
.B2(n_227),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_209),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_210),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_24),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_258),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_259),
.B(n_266),
.Y(n_270)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_219),
.B(n_224),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_268),
.B(n_269),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_215),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_231),
.C(n_243),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_265),
.Y(n_281)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_267),
.B(n_251),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_223),
.B(n_9),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_238),
.A2(n_223),
.B(n_2),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_233),
.B(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_11),
.C(n_14),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_234),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_260),
.B(n_20),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_268),
.B(n_269),
.C(n_265),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_240),
.C(n_243),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_283),
.Y(n_291)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_8),
.C(n_15),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_8),
.C(n_14),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_7),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_260),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_286),
.C(n_287),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_279),
.A2(n_272),
.B1(n_276),
.B2(n_254),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_280),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_7),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_7),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_292),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_276),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_297),
.Y(n_306)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_295),
.A2(n_275),
.A3(n_273),
.B1(n_280),
.B2(n_270),
.C1(n_11),
.C2(n_12),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_12),
.C(n_13),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_303),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_291),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_20),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_10),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_293),
.B(n_287),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_310),
.B(n_311),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_20),
.B(n_13),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_13),
.C(n_5),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_315),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_4),
.B(n_5),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_318),
.C(n_320),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_313),
.A2(n_300),
.B1(n_302),
.B2(n_6),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_6),
.B1(n_319),
.B2(n_321),
.Y(n_323)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_323),
.Y(n_324)
);

XNOR2x2_ASAP7_75t_SL g325 ( 
.A(n_324),
.B(n_6),
.Y(n_325)
);


endmodule