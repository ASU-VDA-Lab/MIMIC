module fake_ariane_3272_n_1710 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1710);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1710;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_114),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_100),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_65),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_3),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_137),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_82),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_107),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_47),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_116),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_86),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_117),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_85),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_120),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_68),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_1),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_6),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_49),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_94),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_56),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_21),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_88),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_118),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_81),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_40),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_43),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_61),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_29),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_10),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_15),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_52),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_57),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_20),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_35),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_78),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_26),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_22),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_51),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_90),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_20),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_48),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_98),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_127),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_99),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_62),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_34),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_92),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_136),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_122),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_54),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_45),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_7),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_74),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_32),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_12),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_22),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_66),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_17),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_47),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_110),
.Y(n_231)
);

BUFx8_ASAP7_75t_SL g232 ( 
.A(n_121),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_139),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_111),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_73),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_84),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_5),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_53),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_145),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_143),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_103),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_67),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_72),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_21),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_80),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_44),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_16),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_44),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_41),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_13),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_64),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_25),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_95),
.Y(n_257)
);

BUFx8_ASAP7_75t_SL g258 ( 
.A(n_146),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_87),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_25),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_93),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_9),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_13),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_23),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_115),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_36),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_23),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_104),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_96),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_147),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_125),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_48),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_34),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_150),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_30),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_141),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_15),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_39),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_42),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_16),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_19),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_58),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_91),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_26),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_3),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_134),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_133),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_39),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_59),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_4),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_10),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_38),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_45),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_9),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_29),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_75),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_70),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_37),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_0),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_71),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_226),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_253),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_253),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_253),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_232),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_253),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_258),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_158),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_177),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_188),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_250),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_260),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_278),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_160),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_278),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_160),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_189),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_212),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_191),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_192),
.Y(n_336)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_252),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_212),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_229),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_175),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_274),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_267),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_175),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_211),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_196),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_229),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_201),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_229),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_229),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_230),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_230),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_164),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_266),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_230),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_274),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_276),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_230),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_249),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_270),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_249),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_202),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_249),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_249),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_167),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_167),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_261),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_281),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_281),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_204),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_155),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_182),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_155),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_194),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_194),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_200),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_200),
.Y(n_377)
);

CKINVDCx6p67_ASAP7_75t_R g378 ( 
.A(n_338),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_315),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_315),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_309),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_340),
.B(n_208),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_304),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_326),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_304),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g386 ( 
.A(n_305),
.B(n_228),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_151),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_305),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_372),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_306),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_307),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_307),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_221),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_311),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_329),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_308),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_310),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_310),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

NOR2x1_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_261),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_221),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_313),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_314),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_331),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_314),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_354),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_318),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_319),
.B(n_228),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_319),
.Y(n_416)
);

AND3x2_ASAP7_75t_L g417 ( 
.A(n_321),
.B(n_353),
.C(n_344),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_322),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_322),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_317),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_341),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_324),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_356),
.B(n_182),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_324),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_320),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_325),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_L g429 ( 
.A(n_330),
.B(n_205),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_333),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_327),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_327),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_336),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_360),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_345),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_328),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_328),
.B(n_152),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_332),
.A2(n_162),
.B(n_156),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_332),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_334),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_334),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_335),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_335),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_339),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_371),
.B(n_373),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_430),
.A2(n_337),
.B1(n_293),
.B2(n_295),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_343),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_430),
.B(n_347),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_379),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_425),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_436),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g455 ( 
.A(n_411),
.B(n_271),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_411),
.B(n_303),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_R g462 ( 
.A(n_434),
.B(n_316),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_362),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_385),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_427),
.B(n_370),
.Y(n_468)
);

AND3x2_ASAP7_75t_L g469 ( 
.A(n_421),
.B(n_286),
.C(n_282),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_395),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_408),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_394),
.B(n_271),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_385),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_421),
.B(n_342),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_387),
.B(n_373),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_386),
.A2(n_292),
.B1(n_287),
.B2(n_294),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_386),
.B(n_374),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_394),
.B(n_352),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_398),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_386),
.B(n_374),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_398),
.Y(n_487)
);

INVx8_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

AO22x2_ASAP7_75t_L g489 ( 
.A1(n_394),
.A2(n_210),
.B1(n_377),
.B2(n_375),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_386),
.B(n_415),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_391),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_417),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_387),
.B(n_375),
.Y(n_495)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_389),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_417),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_389),
.B(n_161),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_382),
.B(n_415),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_425),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_389),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_389),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_406),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_415),
.B(n_376),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_423),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_415),
.B(n_376),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_L g512 ( 
.A(n_406),
.B(n_161),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_424),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_424),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_406),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_382),
.B(n_163),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_441),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_394),
.B(n_163),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_442),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_391),
.B(n_392),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_406),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_446),
.B(n_165),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_404),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_392),
.B(n_377),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_446),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_446),
.B(n_165),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_443),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_443),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_393),
.B(n_348),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_435),
.B(n_233),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_393),
.B(n_301),
.C(n_296),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_406),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_409),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_446),
.B(n_166),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_406),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_396),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_429),
.B(n_357),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_404),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_416),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_446),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_416),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_384),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_439),
.A2(n_288),
.B1(n_270),
.B2(n_236),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_438),
.B(n_166),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_416),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_438),
.B(n_172),
.Y(n_554)
);

INVx6_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

INVx8_ASAP7_75t_L g556 ( 
.A(n_400),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_416),
.B(n_172),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_396),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_416),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_426),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_426),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_390),
.A2(n_235),
.B1(n_263),
.B2(n_290),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_426),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_399),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_399),
.B(n_168),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_426),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_400),
.B(n_173),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_397),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_426),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_422),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_403),
.B(n_366),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_390),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_401),
.B(n_348),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_401),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_426),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_426),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_407),
.B(n_349),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_407),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_431),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_431),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_431),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_403),
.B(n_366),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_413),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_431),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_413),
.B(n_349),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_414),
.Y(n_586)
);

INVxp33_ASAP7_75t_SL g587 ( 
.A(n_378),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_431),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_431),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_431),
.Y(n_590)
);

AO21x2_ASAP7_75t_L g591 ( 
.A1(n_414),
.A2(n_178),
.B(n_170),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_400),
.B(n_173),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_439),
.A2(n_235),
.B1(n_290),
.B2(n_263),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_418),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_400),
.B(n_174),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_418),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_450),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_493),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_544),
.B(n_400),
.Y(n_599)
);

NAND2x1p5_ASAP7_75t_L g600 ( 
.A(n_531),
.B(n_439),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_478),
.B(n_470),
.Y(n_601)
);

INVx8_ASAP7_75t_L g602 ( 
.A(n_488),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_583),
.B(n_405),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_459),
.B(n_478),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_549),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_447),
.B(n_169),
.C(n_164),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_479),
.B(n_405),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_459),
.B(n_378),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_495),
.B(n_405),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_501),
.B(n_405),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_531),
.A2(n_428),
.B1(n_444),
.B2(n_440),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_463),
.B(n_405),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_450),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_547),
.B(n_455),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_524),
.A2(n_420),
.B(n_419),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_547),
.B(n_410),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_493),
.B(n_439),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_455),
.B(n_410),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_455),
.B(n_410),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_454),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_455),
.B(n_410),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_583),
.B(n_174),
.Y(n_623)
);

INVx8_ASAP7_75t_L g624 ( 
.A(n_488),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_455),
.B(n_571),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_564),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_519),
.B(n_410),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_564),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_540),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_454),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_540),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_543),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_448),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_448),
.B(n_378),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_583),
.B(n_298),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_543),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_528),
.B(n_420),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_455),
.B(n_428),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_571),
.B(n_432),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_470),
.B(n_435),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_457),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_491),
.A2(n_432),
.B1(n_444),
.B2(n_440),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_528),
.B(n_433),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_528),
.B(n_433),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_457),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_481),
.A2(n_439),
.B1(n_233),
.B2(n_288),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_558),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_460),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_460),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_558),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_574),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_471),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_545),
.B(n_298),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_593),
.A2(n_270),
.B1(n_288),
.B2(n_445),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_582),
.B(n_437),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_545),
.B(n_437),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_545),
.B(n_291),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_593),
.A2(n_445),
.B1(n_412),
.B2(n_291),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_574),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_473),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_527),
.B(n_412),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_578),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_578),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_461),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_461),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_473),
.B(n_169),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_483),
.B(n_412),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_483),
.B(n_412),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_586),
.A2(n_293),
.B1(n_295),
.B2(n_297),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_556),
.B(n_209),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_565),
.A2(n_207),
.B(n_193),
.C(n_195),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_448),
.B(n_368),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_466),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_SL g674 ( 
.A1(n_562),
.A2(n_297),
.B1(n_300),
.B2(n_227),
.Y(n_674)
);

NOR3xp33_ASAP7_75t_L g675 ( 
.A(n_468),
.B(n_227),
.C(n_300),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_466),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_483),
.B(n_171),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_456),
.B(n_181),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_586),
.A2(n_240),
.B1(n_239),
.B2(n_254),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_448),
.B(n_368),
.Y(n_680)
);

INVxp33_ASAP7_75t_L g681 ( 
.A(n_562),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_568),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_483),
.B(n_184),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_472),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_488),
.B(n_217),
.Y(n_685)
);

CKINVDCx14_ASAP7_75t_R g686 ( 
.A(n_471),
.Y(n_686)
);

NOR2xp67_ASAP7_75t_L g687 ( 
.A(n_570),
.B(n_369),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_532),
.B(n_222),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_594),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_456),
.B(n_197),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_594),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_488),
.B(n_223),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_541),
.B(n_225),
.Y(n_693)
);

NOR3xp33_ASAP7_75t_L g694 ( 
.A(n_449),
.B(n_247),
.C(n_251),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_488),
.B(n_262),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_482),
.B(n_486),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_494),
.B(n_369),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_507),
.B(n_264),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_510),
.B(n_272),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_472),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_572),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_476),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_476),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_552),
.B(n_273),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_596),
.B(n_279),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_484),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_596),
.B(n_280),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_474),
.B(n_283),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_484),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_474),
.B(n_153),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_474),
.B(n_154),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_474),
.A2(n_198),
.B1(n_218),
.B2(n_219),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_489),
.A2(n_591),
.B1(n_474),
.B2(n_550),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_474),
.B(n_451),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_492),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_474),
.B(n_157),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_451),
.B(n_159),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_458),
.B(n_176),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_458),
.B(n_179),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_464),
.B(n_180),
.Y(n_720)
);

NAND2x1p5_ASAP7_75t_L g721 ( 
.A(n_494),
.B(n_224),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_465),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_464),
.B(n_185),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_492),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_467),
.B(n_186),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_467),
.B(n_187),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_456),
.B(n_237),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_529),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_465),
.B(n_346),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_475),
.B(n_190),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_506),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_477),
.B(n_199),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_489),
.A2(n_445),
.B1(n_299),
.B2(n_284),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_506),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_456),
.B(n_238),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_535),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_554),
.B(n_241),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_508),
.Y(n_738)
);

BUFx5_ASAP7_75t_L g739 ( 
.A(n_477),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_480),
.B(n_487),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_499),
.B(n_244),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_573),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_465),
.B(n_203),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_577),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_585),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_556),
.A2(n_248),
.B1(n_255),
.B2(n_259),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_508),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_480),
.B(n_206),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_487),
.B(n_213),
.Y(n_749)
);

INVxp33_ASAP7_75t_L g750 ( 
.A(n_453),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_509),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_485),
.B(n_277),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_490),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_499),
.B(n_346),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_490),
.B(n_214),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_485),
.B(n_183),
.Y(n_756)
);

BUFx12f_ASAP7_75t_L g757 ( 
.A(n_453),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_497),
.B(n_511),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_509),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_513),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_L g761 ( 
.A1(n_536),
.A2(n_364),
.B1(n_363),
.B2(n_361),
.C(n_358),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_522),
.B(n_0),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_497),
.B(n_215),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_511),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_518),
.B(n_216),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_SL g766 ( 
.A(n_652),
.B(n_462),
.C(n_592),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_599),
.A2(n_556),
.B1(n_595),
.B2(n_567),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_632),
.Y(n_768)
);

BUFx4f_ASAP7_75t_L g769 ( 
.A(n_757),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_SL g770 ( 
.A(n_607),
.B(n_538),
.C(n_518),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_SL g771 ( 
.A1(n_637),
.A2(n_517),
.B(n_590),
.C(n_553),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_637),
.B(n_489),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_643),
.B(n_587),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_636),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_643),
.B(n_489),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_633),
.A2(n_587),
.B1(n_500),
.B2(n_512),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_728),
.B(n_521),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_597),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_647),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_650),
.Y(n_780)
);

NOR3xp33_ASAP7_75t_SL g781 ( 
.A(n_653),
.B(n_538),
.C(n_285),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_697),
.B(n_521),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_634),
.B(n_556),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_614),
.Y(n_784)
);

NAND2x1p5_ASAP7_75t_L g785 ( 
.A(n_598),
.B(n_533),
.Y(n_785)
);

NOR2x1p5_ASAP7_75t_L g786 ( 
.A(n_722),
.B(n_452),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_697),
.B(n_533),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_651),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_659),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_614),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_662),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_663),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_660),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_696),
.B(n_513),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_621),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_646),
.A2(n_658),
.B1(n_733),
.B2(n_674),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_602),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_736),
.B(n_515),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_605),
.A2(n_500),
.B1(n_512),
.B2(n_557),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_742),
.B(n_515),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_602),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_621),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_615),
.B(n_619),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_611),
.A2(n_610),
.B(n_608),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_701),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_600),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_630),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_624),
.B(n_629),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_744),
.B(n_516),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_757),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_646),
.A2(n_591),
.B1(n_534),
.B2(n_530),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_745),
.B(n_516),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_689),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_639),
.B(n_520),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_631),
.B(n_485),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_691),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_762),
.A2(n_557),
.B1(n_555),
.B2(n_496),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_630),
.Y(n_818)
);

AND2x6_ASAP7_75t_SL g819 ( 
.A(n_640),
.B(n_634),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_762),
.A2(n_555),
.B1(n_496),
.B2(n_503),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_658),
.A2(n_591),
.B1(n_537),
.B2(n_534),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_609),
.B(n_498),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_688),
.A2(n_693),
.B1(n_704),
.B2(n_672),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_733),
.A2(n_537),
.B1(n_526),
.B2(n_523),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_655),
.B(n_520),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_722),
.B(n_498),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_613),
.A2(n_542),
.B(n_589),
.Y(n_827)
);

NOR2x2_ASAP7_75t_L g828 ( 
.A(n_634),
.B(n_502),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_604),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_753),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_698),
.B(n_523),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_764),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_601),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_699),
.B(n_526),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_680),
.B(n_469),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_688),
.A2(n_555),
.B1(n_496),
.B2(n_503),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_672),
.B(n_498),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_606),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_721),
.B(n_530),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_721),
.B(n_590),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_729),
.B(n_503),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_682),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_741),
.B(n_514),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_754),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_641),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_754),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_686),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_685),
.B(n_498),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_741),
.B(n_514),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_713),
.A2(n_548),
.B1(n_589),
.B2(n_588),
.Y(n_850)
);

INVx5_ASAP7_75t_L g851 ( 
.A(n_604),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_645),
.Y(n_852)
);

CKINVDCx6p67_ASAP7_75t_R g853 ( 
.A(n_666),
.Y(n_853)
);

INVx5_ASAP7_75t_L g854 ( 
.A(n_604),
.Y(n_854)
);

AND2x6_ASAP7_75t_L g855 ( 
.A(n_620),
.B(n_622),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_645),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_693),
.A2(n_555),
.B1(n_496),
.B2(n_553),
.Y(n_857)
);

NAND2xp33_ASAP7_75t_L g858 ( 
.A(n_739),
.B(n_498),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_648),
.Y(n_859)
);

AO22x1_ASAP7_75t_L g860 ( 
.A1(n_681),
.A2(n_242),
.B1(n_231),
.B2(n_234),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_743),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_739),
.B(n_504),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_667),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_740),
.A2(n_560),
.B(n_588),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_677),
.B(n_514),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_750),
.B(n_517),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_683),
.B(n_590),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_669),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_626),
.B(n_517),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_687),
.B(n_525),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_692),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_628),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_648),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_668),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_625),
.B(n_542),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_604),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_708),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_737),
.B(n_525),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_649),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_737),
.B(n_525),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_684),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_SL g882 ( 
.A(n_746),
.B(n_220),
.Y(n_882)
);

BUFx3_ASAP7_75t_L g883 ( 
.A(n_704),
.Y(n_883)
);

AOI211xp5_ASAP7_75t_L g884 ( 
.A1(n_675),
.A2(n_584),
.B(n_581),
.C(n_580),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_649),
.Y(n_885)
);

BUFx2_ASAP7_75t_SL g886 ( 
.A(n_695),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_627),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_705),
.B(n_539),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_644),
.B(n_539),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_644),
.A2(n_539),
.B1(n_553),
.B2(n_580),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_664),
.Y(n_891)
);

NOR2x1p5_ASAP7_75t_L g892 ( 
.A(n_707),
.B(n_546),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_656),
.B(n_657),
.Y(n_893)
);

AND3x1_ASAP7_75t_L g894 ( 
.A(n_694),
.B(n_584),
.C(n_581),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_654),
.B(n_548),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_684),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_713),
.A2(n_579),
.B1(n_576),
.B2(n_575),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_700),
.Y(n_898)
);

NOR2x1_ASAP7_75t_L g899 ( 
.A(n_623),
.B(n_551),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_600),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_635),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_654),
.B(n_551),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_679),
.B(n_355),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_627),
.B(n_560),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_661),
.A2(n_575),
.B1(n_569),
.B2(n_563),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_603),
.B(n_714),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_603),
.B(n_561),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_700),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_702),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_765),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_618),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_758),
.A2(n_569),
.B(n_563),
.Y(n_912)
);

INVxp67_ASAP7_75t_L g913 ( 
.A(n_661),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_717),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_638),
.B(n_559),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_739),
.B(n_617),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_718),
.B(n_559),
.Y(n_917)
);

OR2x2_ASAP7_75t_SL g918 ( 
.A(n_710),
.B(n_183),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_612),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_703),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_618),
.Y(n_921)
);

OR2x2_ASAP7_75t_SL g922 ( 
.A(n_711),
.B(n_716),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_739),
.B(n_559),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_703),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_706),
.B(n_559),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_706),
.A2(n_709),
.B1(n_724),
.B2(n_760),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_709),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_715),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_719),
.B(n_504),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_720),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_761),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_715),
.B(n_504),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_724),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_731),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_731),
.B(n_504),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_665),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_712),
.B(n_566),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_SL g938 ( 
.A(n_723),
.B(n_725),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_665),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_726),
.B(n_566),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_734),
.B(n_566),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_734),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_738),
.Y(n_943)
);

O2A1O1Ixp5_ASAP7_75t_L g944 ( 
.A1(n_938),
.A2(n_642),
.B(n_690),
.C(n_678),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_823),
.B(n_738),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_910),
.B(n_730),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_883),
.B(n_931),
.Y(n_947)
);

OAI21xp33_ASAP7_75t_L g948 ( 
.A1(n_868),
.A2(n_671),
.B(n_670),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_SL g949 ( 
.A1(n_893),
.A2(n_616),
.B(n_749),
.C(n_748),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_797),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_919),
.A2(n_763),
.B1(n_732),
.B2(n_755),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_SL g952 ( 
.A(n_847),
.B(n_735),
.C(n_678),
.Y(n_952)
);

AO32x2_ASAP7_75t_L g953 ( 
.A1(n_871),
.A2(n_901),
.A3(n_767),
.B1(n_771),
.B2(n_796),
.Y(n_953)
);

O2A1O1Ixp5_ASAP7_75t_L g954 ( 
.A1(n_848),
.A2(n_690),
.B(n_727),
.C(n_752),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_838),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_R g956 ( 
.A(n_769),
.B(n_747),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_773),
.B(n_727),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_797),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_778),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_SL g960 ( 
.A1(n_796),
.A2(n_302),
.B1(n_243),
.B2(n_245),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_914),
.B(n_751),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_769),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_784),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_R g964 ( 
.A(n_766),
.B(n_759),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_882),
.A2(n_833),
.B1(n_853),
.B2(n_893),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_833),
.B(n_751),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_827),
.A2(n_676),
.B(n_673),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_790),
.Y(n_968)
);

OAI21xp33_ASAP7_75t_L g969 ( 
.A1(n_887),
.A2(n_289),
.B(n_246),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_804),
.A2(n_566),
.B(n_505),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_887),
.B(n_566),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_913),
.A2(n_505),
.B(n_756),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_863),
.B(n_874),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_793),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_768),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_913),
.A2(n_505),
.B(n_756),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_923),
.A2(n_505),
.B(n_257),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_774),
.Y(n_978)
);

NAND3xp33_ASAP7_75t_SL g979 ( 
.A(n_861),
.B(n_265),
.C(n_268),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_793),
.A2(n_269),
.B1(n_275),
.B2(n_361),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_842),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_786),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_779),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_862),
.A2(n_916),
.B(n_794),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_795),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_884),
.B(n_351),
.C(n_350),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_SL g987 ( 
.A(n_801),
.B(n_183),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_930),
.B(n_2),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_SL g989 ( 
.A1(n_810),
.A2(n_783),
.B1(n_776),
.B2(n_894),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_801),
.B(n_8),
.Y(n_990)
);

O2A1O1Ixp5_ASAP7_75t_L g991 ( 
.A1(n_940),
.A2(n_8),
.B(n_11),
.C(n_12),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_783),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_930),
.A2(n_14),
.B(n_18),
.C(n_24),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_777),
.A2(n_789),
.B1(n_780),
.B2(n_813),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_822),
.A2(n_14),
.B(n_18),
.C(n_24),
.Y(n_995)
);

INVxp67_ASAP7_75t_L g996 ( 
.A(n_805),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_872),
.Y(n_997)
);

AO32x2_ASAP7_75t_L g998 ( 
.A1(n_771),
.A2(n_775),
.A3(n_772),
.B1(n_811),
.B2(n_922),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_783),
.B(n_27),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_835),
.B(n_27),
.Y(n_1000)
);

INVx1_ASAP7_75t_SL g1001 ( 
.A(n_866),
.Y(n_1001)
);

OR2x4_ASAP7_75t_L g1002 ( 
.A(n_788),
.B(n_28),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_844),
.B(n_28),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_SL g1004 ( 
.A1(n_889),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_R g1005 ( 
.A(n_819),
.B(n_76),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_841),
.B(n_31),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_791),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_R g1008 ( 
.A(n_886),
.B(n_33),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_808),
.B(n_36),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_792),
.B(n_37),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_903),
.B(n_38),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_802),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_846),
.B(n_40),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_862),
.A2(n_89),
.B(n_140),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_841),
.B(n_41),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_916),
.A2(n_97),
.B(n_132),
.Y(n_1016)
);

OA22x2_ASAP7_75t_L g1017 ( 
.A1(n_816),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_837),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_770),
.A2(n_46),
.B(n_50),
.C(n_55),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_830),
.B(n_63),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_832),
.B(n_69),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_799),
.A2(n_102),
.B1(n_109),
.B2(n_112),
.Y(n_1022)
);

NOR2x1_ASAP7_75t_L g1023 ( 
.A(n_770),
.B(n_826),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_940),
.A2(n_126),
.B(n_128),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_828),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_906),
.B(n_131),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_888),
.A2(n_815),
.B(n_880),
.C(n_878),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_782),
.A2(n_787),
.B1(n_811),
.B2(n_825),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_781),
.A2(n_929),
.B(n_917),
.C(n_906),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_911),
.B(n_921),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_864),
.A2(n_912),
.B(n_904),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_R g1032 ( 
.A(n_851),
.B(n_854),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_864),
.A2(n_912),
.B(n_917),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_781),
.B(n_860),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_851),
.B(n_854),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_870),
.A2(n_892),
.B1(n_803),
.B2(n_855),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_870),
.A2(n_803),
.B1(n_855),
.B2(n_915),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_854),
.B(n_876),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_920),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_929),
.A2(n_831),
.B(n_834),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_814),
.B(n_798),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_865),
.A2(n_867),
.B(n_869),
.C(n_809),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_898),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_895),
.A2(n_902),
.B(n_935),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_925),
.A2(n_932),
.B(n_941),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_800),
.B(n_812),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_909),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_877),
.B(n_881),
.Y(n_1048)
);

AO32x1_ASAP7_75t_L g1049 ( 
.A1(n_924),
.A2(n_928),
.A3(n_942),
.B1(n_933),
.B2(n_934),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_806),
.A2(n_900),
.B(n_915),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_806),
.A2(n_900),
.B(n_907),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_807),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_839),
.B(n_879),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_817),
.A2(n_824),
.B1(n_857),
.B2(n_820),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_818),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_876),
.B(n_849),
.Y(n_1056)
);

INVx4_ASAP7_75t_L g1057 ( 
.A(n_876),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_845),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_824),
.A2(n_836),
.B1(n_821),
.B2(n_785),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_785),
.A2(n_843),
.B(n_840),
.C(n_907),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_899),
.A2(n_829),
.B(n_937),
.C(n_896),
.Y(n_1061)
);

NAND3xp33_ASAP7_75t_SL g1062 ( 
.A(n_890),
.B(n_905),
.C(n_821),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_850),
.A2(n_897),
.B(n_855),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_908),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_927),
.A2(n_897),
.B(n_850),
.C(n_852),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_856),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_911),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_943),
.B(n_911),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_859),
.B(n_939),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_873),
.B(n_936),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_885),
.B(n_891),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_1035),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_1031),
.A2(n_926),
.B(n_918),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_947),
.B(n_943),
.Y(n_1074)
);

INVx5_ASAP7_75t_L g1075 ( 
.A(n_1035),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1070),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_974),
.B(n_926),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_965),
.B(n_921),
.Y(n_1078)
);

OR2x6_ASAP7_75t_L g1079 ( 
.A(n_999),
.B(n_803),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_1059),
.A2(n_803),
.A3(n_875),
.B(n_1054),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_994),
.A2(n_973),
.B1(n_988),
.B2(n_1010),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_951),
.A2(n_949),
.B(n_1041),
.Y(n_1082)
);

NOR4xp25_ASAP7_75t_L g1083 ( 
.A(n_993),
.B(n_875),
.C(n_948),
.D(n_1019),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_967),
.A2(n_875),
.B(n_1045),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_981),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_973),
.B(n_875),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_992),
.B(n_962),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_SL g1088 ( 
.A1(n_945),
.A2(n_1028),
.B(n_1046),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_984),
.A2(n_970),
.B(n_1044),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_SL g1090 ( 
.A1(n_971),
.A2(n_951),
.B(n_1029),
.C(n_1004),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1054),
.A2(n_1042),
.B(n_1027),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_944),
.A2(n_1023),
.B(n_1022),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1020),
.A2(n_1021),
.B(n_957),
.C(n_1011),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_975),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1022),
.A2(n_1062),
.B(n_991),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1060),
.A2(n_976),
.B(n_972),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_961),
.B(n_1001),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_960),
.A2(n_1000),
.B1(n_1017),
.B2(n_989),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1051),
.A2(n_1024),
.B(n_1016),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1001),
.B(n_966),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_946),
.A2(n_1015),
.B(n_1006),
.C(n_1009),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_955),
.Y(n_1102)
);

CKINVDCx11_ASAP7_75t_R g1103 ( 
.A(n_997),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_992),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_978),
.B(n_983),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1007),
.B(n_1039),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1050),
.A2(n_954),
.B(n_977),
.Y(n_1107)
);

INVx3_ASAP7_75t_SL g1108 ( 
.A(n_982),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1065),
.A2(n_1063),
.B(n_1028),
.Y(n_1109)
);

AND3x4_ASAP7_75t_L g1110 ( 
.A(n_999),
.B(n_952),
.C(n_1003),
.Y(n_1110)
);

NOR2x1_ASAP7_75t_SL g1111 ( 
.A(n_1030),
.B(n_1038),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1043),
.Y(n_1112)
);

AOI31xp67_ASAP7_75t_L g1113 ( 
.A1(n_1036),
.A2(n_1037),
.A3(n_1056),
.B(n_1026),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_959),
.Y(n_1114)
);

OAI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1002),
.A2(n_1017),
.B1(n_980),
.B2(n_1063),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1061),
.A2(n_1014),
.B(n_1068),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_1069),
.A2(n_1049),
.A3(n_1047),
.B(n_1071),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1034),
.A2(n_969),
.B(n_995),
.C(n_1013),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1048),
.B(n_1003),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1032),
.B(n_950),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_956),
.Y(n_1121)
);

INVx6_ASAP7_75t_SL g1122 ( 
.A(n_1030),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_996),
.B(n_979),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_1049),
.A2(n_1071),
.A3(n_1055),
.B(n_1052),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1058),
.Y(n_1125)
);

AOI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_964),
.A2(n_986),
.B(n_1053),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_950),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_963),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_1025),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_958),
.A2(n_1012),
.B(n_1066),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_968),
.A2(n_985),
.B(n_1064),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1018),
.B(n_1008),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1067),
.B(n_1057),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_990),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1002),
.B(n_950),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1067),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1067),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_953),
.A2(n_998),
.B(n_987),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1005),
.A2(n_1057),
.B1(n_953),
.B2(n_998),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_998),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_948),
.A2(n_823),
.B(n_883),
.C(n_762),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1054),
.A2(n_913),
.B(n_887),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_975),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1031),
.A2(n_967),
.B(n_1033),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_973),
.B(n_1041),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_965),
.B(n_823),
.Y(n_1146)
);

NOR4xp25_ASAP7_75t_L g1147 ( 
.A(n_993),
.B(n_796),
.C(n_948),
.D(n_1019),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_975),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_975),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_955),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1152)
);

INVxp67_ASAP7_75t_SL g1153 ( 
.A(n_974),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1033),
.A2(n_1059),
.A3(n_1040),
.B(n_1054),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_955),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1031),
.A2(n_967),
.B(n_1033),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_1063),
.B(n_587),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_SL g1158 ( 
.A1(n_994),
.A2(n_1041),
.B(n_945),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_975),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1160)
);

NOR2xp67_ASAP7_75t_SL g1161 ( 
.A(n_962),
.B(n_652),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1033),
.A2(n_1031),
.B(n_1063),
.Y(n_1162)
);

OR2x6_ASAP7_75t_L g1163 ( 
.A(n_999),
.B(n_783),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1035),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_975),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_975),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_947),
.B(n_605),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_955),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1031),
.A2(n_967),
.B(n_1033),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_994),
.A2(n_823),
.B1(n_919),
.B2(n_796),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_965),
.B(n_823),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1033),
.A2(n_1031),
.B(n_1063),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_947),
.B(n_338),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_960),
.A2(n_823),
.B1(n_868),
.B2(n_796),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_947),
.B(n_833),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_1033),
.A2(n_1059),
.A3(n_1040),
.B(n_1054),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_947),
.B(n_605),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1054),
.A2(n_913),
.B(n_887),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1070),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1070),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_994),
.A2(n_823),
.B1(n_919),
.B2(n_796),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_947),
.B(n_338),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1054),
.A2(n_913),
.B(n_887),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_965),
.B(n_823),
.Y(n_1188)
);

INVx5_ASAP7_75t_L g1189 ( 
.A(n_1035),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_SL g1190 ( 
.A1(n_994),
.A2(n_973),
.B(n_1060),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1031),
.A2(n_967),
.B(n_1033),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1033),
.A2(n_1059),
.A3(n_1040),
.B(n_1054),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_975),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_948),
.A2(n_823),
.B(n_883),
.C(n_762),
.Y(n_1194)
);

NOR4xp25_ASAP7_75t_L g1195 ( 
.A(n_993),
.B(n_796),
.C(n_948),
.D(n_1019),
.Y(n_1195)
);

OAI22x1_ASAP7_75t_L g1196 ( 
.A1(n_965),
.A2(n_823),
.B1(n_593),
.B2(n_425),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_975),
.Y(n_1197)
);

BUFx12f_ASAP7_75t_L g1198 ( 
.A(n_962),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_948),
.A2(n_823),
.B(n_883),
.C(n_762),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_947),
.B(n_605),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_975),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1033),
.A2(n_858),
.B(n_804),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_SL g1204 ( 
.A1(n_1081),
.A2(n_1190),
.B(n_1180),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1153),
.B(n_1106),
.Y(n_1205)
);

NOR3xp33_ASAP7_75t_L g1206 ( 
.A(n_1081),
.B(n_1093),
.C(n_1170),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1174),
.A2(n_1098),
.B1(n_1170),
.B2(n_1184),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_1077),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1184),
.A2(n_1141),
.B(n_1194),
.C(n_1200),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1144),
.A2(n_1169),
.B(n_1156),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1105),
.Y(n_1211)
);

OAI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1174),
.A2(n_1098),
.B1(n_1157),
.B2(n_1115),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1175),
.B(n_1167),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1196),
.A2(n_1188),
.B1(n_1146),
.B2(n_1171),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1100),
.B(n_1094),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1157),
.A2(n_1109),
.B1(n_1180),
.B2(n_1186),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1142),
.A2(n_1186),
.B1(n_1110),
.B2(n_1095),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1072),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1150),
.A2(n_1203),
.B(n_1199),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1143),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1124),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1148),
.Y(n_1222)
);

BUFx4_ASAP7_75t_SL g1223 ( 
.A(n_1129),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1152),
.A2(n_1160),
.B(n_1179),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1149),
.Y(n_1225)
);

CKINVDCx14_ASAP7_75t_R g1226 ( 
.A(n_1103),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1159),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1191),
.A2(n_1089),
.B(n_1187),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1178),
.A2(n_1181),
.B(n_1099),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1155),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1198),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1165),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1161),
.B(n_1102),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1084),
.A2(n_1096),
.B(n_1107),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1173),
.B(n_1185),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1166),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1193),
.Y(n_1237)
);

INVx6_ASAP7_75t_L g1238 ( 
.A(n_1075),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1123),
.A2(n_1177),
.B1(n_1201),
.B2(n_1135),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1102),
.B(n_1119),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1142),
.A2(n_1092),
.B1(n_1118),
.B2(n_1091),
.Y(n_1241)
);

INVx8_ASAP7_75t_L g1242 ( 
.A(n_1163),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1138),
.A2(n_1109),
.B(n_1082),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1197),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1151),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1079),
.A2(n_1101),
.B1(n_1145),
.B2(n_1134),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1116),
.A2(n_1130),
.B(n_1172),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1087),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1145),
.B(n_1097),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1202),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1140),
.A2(n_1139),
.B1(n_1126),
.B2(n_1182),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1117),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1131),
.A2(n_1086),
.B(n_1126),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_1147),
.B(n_1195),
.C(n_1158),
.Y(n_1254)
);

CKINVDCx11_ASAP7_75t_R g1255 ( 
.A(n_1108),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_SL g1256 ( 
.A(n_1121),
.B(n_1189),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1088),
.A2(n_1162),
.B(n_1090),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1076),
.A2(n_1183),
.B1(n_1079),
.B2(n_1112),
.Y(n_1258)
);

INVx8_ASAP7_75t_L g1259 ( 
.A(n_1163),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1125),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1085),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1122),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1154),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1132),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1086),
.B(n_1128),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1072),
.Y(n_1266)
);

BUFx2_ASAP7_75t_SL g1267 ( 
.A(n_1075),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1114),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1117),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1117),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1147),
.A2(n_1195),
.B(n_1083),
.C(n_1078),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1164),
.B(n_1072),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1189),
.B(n_1164),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_L g1274 ( 
.A(n_1083),
.B(n_1137),
.C(n_1074),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1111),
.A2(n_1080),
.A3(n_1073),
.B(n_1136),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1133),
.A2(n_1192),
.B(n_1176),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1104),
.B(n_1120),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1133),
.A2(n_1113),
.B(n_1154),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1080),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1122),
.A2(n_1080),
.B1(n_1127),
.B2(n_1154),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1176),
.A2(n_1152),
.B(n_1150),
.Y(n_1281)
);

BUFx2_ASAP7_75t_R g1282 ( 
.A(n_1176),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1192),
.B(n_1174),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1192),
.A2(n_1196),
.B1(n_562),
.B2(n_796),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1144),
.A2(n_1169),
.B(n_1156),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_SL g1286 ( 
.A1(n_1081),
.A2(n_1190),
.B(n_1180),
.Y(n_1286)
);

OAI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1098),
.A2(n_1174),
.B1(n_1110),
.B2(n_1171),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1081),
.A2(n_1093),
.B(n_1194),
.C(n_1141),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1175),
.B(n_974),
.Y(n_1289)
);

CKINVDCx6p67_ASAP7_75t_R g1290 ( 
.A(n_1103),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1168),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1145),
.B(n_1167),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1198),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1144),
.A2(n_1169),
.B(n_1156),
.Y(n_1294)
);

AND2x2_ASAP7_75t_SL g1295 ( 
.A(n_1157),
.B(n_1147),
.Y(n_1295)
);

BUFx8_ASAP7_75t_L g1296 ( 
.A(n_1198),
.Y(n_1296)
);

AO221x2_ASAP7_75t_L g1297 ( 
.A1(n_1081),
.A2(n_1170),
.B1(n_1184),
.B2(n_1115),
.C(n_1095),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1093),
.A2(n_1081),
.B(n_823),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1196),
.A2(n_562),
.B1(n_796),
.B2(n_1170),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1072),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1144),
.A2(n_1169),
.B(n_1156),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1093),
.A2(n_1081),
.B(n_823),
.Y(n_1302)
);

NAND3xp33_ASAP7_75t_L g1303 ( 
.A(n_1093),
.B(n_1081),
.C(n_1141),
.Y(n_1303)
);

AOI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1091),
.A2(n_1082),
.B(n_1081),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1144),
.A2(n_1169),
.B(n_1156),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1153),
.B(n_1106),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1198),
.Y(n_1307)
);

CKINVDCx16_ASAP7_75t_R g1308 ( 
.A(n_1198),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1168),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1174),
.A2(n_1184),
.B1(n_1170),
.B2(n_1098),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1144),
.A2(n_1169),
.B(n_1156),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1144),
.A2(n_1169),
.B(n_1156),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1174),
.A2(n_1098),
.B1(n_1184),
.B2(n_1170),
.Y(n_1313)
);

BUFx2_ASAP7_75t_SL g1314 ( 
.A(n_1168),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1093),
.A2(n_1174),
.B1(n_1081),
.B2(n_823),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1105),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_SL g1317 ( 
.A(n_1161),
.B(n_652),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1144),
.A2(n_1169),
.B(n_1156),
.Y(n_1318)
);

CKINVDCx14_ASAP7_75t_R g1319 ( 
.A(n_1103),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1093),
.A2(n_1081),
.B(n_823),
.Y(n_1320)
);

AND2x2_ASAP7_75t_SL g1321 ( 
.A(n_1157),
.B(n_1147),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1093),
.A2(n_1174),
.B1(n_1081),
.B2(n_823),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1240),
.B(n_1213),
.Y(n_1323)
);

OA21x2_ASAP7_75t_L g1324 ( 
.A1(n_1219),
.A2(n_1224),
.B(n_1281),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1205),
.B(n_1306),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1298),
.A2(n_1320),
.B(n_1302),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1313),
.A2(n_1216),
.B1(n_1207),
.B2(n_1310),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1216),
.A2(n_1310),
.B1(n_1217),
.B2(n_1322),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1315),
.A2(n_1206),
.B(n_1288),
.C(n_1241),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1206),
.A2(n_1288),
.B(n_1283),
.C(n_1254),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1220),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1289),
.B(n_1245),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1219),
.A2(n_1224),
.B(n_1281),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1314),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1283),
.A2(n_1303),
.B(n_1209),
.C(n_1271),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1208),
.B(n_1274),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1292),
.B(n_1249),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1230),
.B(n_1248),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1287),
.B(n_1239),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1297),
.B(n_1211),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1299),
.A2(n_1212),
.B1(n_1214),
.B2(n_1209),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1222),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1299),
.A2(n_1212),
.B1(n_1214),
.B2(n_1284),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1257),
.A2(n_1297),
.B(n_1204),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1257),
.A2(n_1297),
.B(n_1286),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1284),
.A2(n_1235),
.B1(n_1321),
.B2(n_1295),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1316),
.B(n_1215),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1229),
.A2(n_1228),
.B(n_1234),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1232),
.B(n_1236),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1263),
.Y(n_1351)
);

AOI221x1_ASAP7_75t_SL g1352 ( 
.A1(n_1235),
.A2(n_1246),
.B1(n_1237),
.B2(n_1244),
.C(n_1250),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1296),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1295),
.B(n_1321),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1223),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1261),
.A2(n_1304),
.B1(n_1251),
.B2(n_1258),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1260),
.B(n_1277),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1265),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1291),
.B(n_1309),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1208),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1273),
.A2(n_1276),
.B(n_1231),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1251),
.A2(n_1258),
.B1(n_1264),
.B2(n_1282),
.Y(n_1362)
);

OAI22x1_ASAP7_75t_L g1363 ( 
.A1(n_1262),
.A2(n_1293),
.B1(n_1307),
.B2(n_1276),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1272),
.B(n_1233),
.Y(n_1364)
);

O2A1O1Ixp5_ASAP7_75t_L g1365 ( 
.A1(n_1269),
.A2(n_1270),
.B(n_1279),
.C(n_1252),
.Y(n_1365)
);

O2A1O1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1317),
.A2(n_1243),
.B(n_1231),
.C(n_1256),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1280),
.B(n_1268),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1243),
.A2(n_1218),
.B(n_1266),
.C(n_1300),
.Y(n_1368)
);

OR2x6_ASAP7_75t_L g1369 ( 
.A(n_1242),
.B(n_1259),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1242),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1218),
.B(n_1266),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1300),
.B(n_1319),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1242),
.B(n_1259),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1247),
.A2(n_1278),
.B(n_1210),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1226),
.A2(n_1319),
.B(n_1252),
.C(n_1221),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1253),
.A2(n_1267),
.B(n_1238),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1226),
.B(n_1290),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1308),
.B(n_1238),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1285),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1275),
.B(n_1255),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1285),
.A2(n_1301),
.B(n_1294),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1294),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1301),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1301),
.B(n_1223),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1296),
.A2(n_1305),
.B1(n_1311),
.B2(n_1312),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1318),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1240),
.B(n_1213),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1240),
.B(n_1213),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1313),
.A2(n_1216),
.B1(n_1174),
.B2(n_1207),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1220),
.Y(n_1390)
);

NOR2xp67_ASAP7_75t_L g1391 ( 
.A(n_1208),
.B(n_1274),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1240),
.B(n_1213),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1219),
.A2(n_1224),
.B(n_1281),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1223),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1205),
.B(n_1306),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1219),
.A2(n_1224),
.B(n_1281),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1240),
.B(n_1213),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1315),
.A2(n_1322),
.B(n_1093),
.C(n_1081),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1276),
.Y(n_1399)
);

O2A1O1Ixp5_ASAP7_75t_L g1400 ( 
.A1(n_1298),
.A2(n_1320),
.B(n_1302),
.C(n_1315),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1220),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1220),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1220),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1324),
.B(n_1333),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1382),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1324),
.B(n_1333),
.Y(n_1406)
);

OAI21xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1354),
.A2(n_1328),
.B(n_1344),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1326),
.B(n_1398),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1325),
.B(n_1395),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1335),
.A2(n_1381),
.B(n_1330),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1360),
.B(n_1340),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1374),
.Y(n_1412)
);

AO21x2_ASAP7_75t_L g1413 ( 
.A1(n_1335),
.A2(n_1330),
.B(n_1346),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1343),
.A2(n_1341),
.B1(n_1389),
.B2(n_1327),
.Y(n_1414)
);

NOR2x1_ASAP7_75t_SL g1415 ( 
.A(n_1369),
.B(n_1385),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1324),
.B(n_1333),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1379),
.A2(n_1345),
.B(n_1365),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1386),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1374),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1393),
.B(n_1396),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1399),
.A2(n_1383),
.B(n_1391),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1348),
.B(n_1350),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1331),
.Y(n_1423)
);

AOI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1329),
.A2(n_1400),
.B1(n_1352),
.B2(n_1356),
.C(n_1339),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1342),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1374),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1351),
.B(n_1358),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1351),
.B(n_1390),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1376),
.B(n_1361),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1401),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1400),
.A2(n_1336),
.B(n_1366),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1402),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1403),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1386),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1384),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1368),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1349),
.Y(n_1437)
);

AOI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1363),
.A2(n_1380),
.B(n_1371),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1367),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1332),
.B(n_1323),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1357),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1347),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1362),
.A2(n_1337),
.B(n_1364),
.Y(n_1443)
);

BUFx2_ASAP7_75t_SL g1444 ( 
.A(n_1418),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1404),
.B(n_1397),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1404),
.B(n_1387),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1404),
.B(n_1406),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1427),
.B(n_1388),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1406),
.B(n_1392),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1432),
.B(n_1442),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1421),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1406),
.B(n_1338),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1416),
.B(n_1420),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1416),
.B(n_1420),
.Y(n_1454)
);

CKINVDCx14_ASAP7_75t_R g1455 ( 
.A(n_1434),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1421),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1410),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1414),
.A2(n_1375),
.B1(n_1334),
.B2(n_1378),
.C(n_1355),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1408),
.B(n_1359),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1408),
.A2(n_1369),
.B1(n_1370),
.B2(n_1373),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1405),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1412),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1409),
.B(n_1372),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1437),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1409),
.B(n_1422),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1441),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1457),
.B(n_1415),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1463),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1452),
.Y(n_1469)
);

CKINVDCx16_ASAP7_75t_R g1470 ( 
.A(n_1466),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1457),
.B(n_1415),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1457),
.B(n_1415),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1461),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1459),
.B(n_1394),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1464),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1445),
.B(n_1440),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1457),
.A2(n_1424),
.B1(n_1407),
.B2(n_1431),
.C(n_1414),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1445),
.B(n_1440),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1464),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1448),
.B(n_1422),
.Y(n_1480)
);

OAI211xp5_ASAP7_75t_L g1481 ( 
.A1(n_1459),
.A2(n_1407),
.B(n_1424),
.C(n_1431),
.Y(n_1481)
);

AOI33xp33_ASAP7_75t_L g1482 ( 
.A1(n_1447),
.A2(n_1453),
.A3(n_1454),
.B1(n_1449),
.B2(n_1446),
.B3(n_1445),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1451),
.A2(n_1413),
.B1(n_1436),
.B2(n_1411),
.C(n_1410),
.Y(n_1483)
);

INVx4_ASAP7_75t_L g1484 ( 
.A(n_1462),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1448),
.B(n_1409),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1446),
.B(n_1440),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1446),
.B(n_1435),
.Y(n_1487)
);

AOI211xp5_ASAP7_75t_L g1488 ( 
.A1(n_1458),
.A2(n_1460),
.B(n_1436),
.C(n_1434),
.Y(n_1488)
);

AOI33xp33_ASAP7_75t_L g1489 ( 
.A1(n_1447),
.A2(n_1436),
.A3(n_1430),
.B1(n_1423),
.B2(n_1425),
.B3(n_1433),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1461),
.Y(n_1490)
);

OR2x6_ASAP7_75t_L g1491 ( 
.A(n_1444),
.B(n_1429),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1449),
.B(n_1435),
.Y(n_1492)
);

OAI31xp33_ASAP7_75t_L g1493 ( 
.A1(n_1458),
.A2(n_1413),
.A3(n_1434),
.B(n_1410),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1451),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1466),
.A2(n_1413),
.B1(n_1410),
.B2(n_1443),
.Y(n_1495)
);

OAI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1451),
.A2(n_1411),
.B1(n_1418),
.B2(n_1443),
.C(n_1442),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1452),
.B(n_1441),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1455),
.A2(n_1465),
.B1(n_1463),
.B2(n_1448),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1465),
.B(n_1428),
.Y(n_1499)
);

NAND4xp25_ASAP7_75t_L g1500 ( 
.A(n_1447),
.B(n_1419),
.C(n_1412),
.D(n_1426),
.Y(n_1500)
);

OAI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1456),
.A2(n_1418),
.B1(n_1443),
.B2(n_1442),
.C(n_1438),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1461),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1473),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1494),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1473),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1482),
.B(n_1453),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1490),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1491),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1469),
.B(n_1478),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1475),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1481),
.A2(n_1456),
.B(n_1443),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1493),
.A2(n_1413),
.B(n_1429),
.Y(n_1512)
);

OR2x6_ASAP7_75t_L g1513 ( 
.A(n_1467),
.B(n_1429),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1489),
.B(n_1450),
.Y(n_1514)
);

NOR2x1_ASAP7_75t_L g1515 ( 
.A(n_1500),
.B(n_1377),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1490),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1470),
.B(n_1460),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1502),
.Y(n_1518)
);

INVx4_ASAP7_75t_SL g1519 ( 
.A(n_1491),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1485),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1485),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1499),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1491),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1475),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1479),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1499),
.Y(n_1526)
);

NOR2x1p5_ASAP7_75t_L g1527 ( 
.A(n_1500),
.B(n_1463),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1480),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1480),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1494),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1493),
.A2(n_1429),
.B(n_1417),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1494),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1503),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1532),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1527),
.B(n_1478),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1514),
.B(n_1468),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1519),
.B(n_1494),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1514),
.B(n_1450),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1528),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1511),
.B(n_1483),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1510),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1503),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1510),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1527),
.B(n_1486),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1507),
.Y(n_1545)
);

NOR2xp67_ASAP7_75t_L g1546 ( 
.A(n_1523),
.B(n_1504),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1520),
.B(n_1476),
.Y(n_1547)
);

AOI221xp5_ASAP7_75t_L g1548 ( 
.A1(n_1511),
.A2(n_1496),
.B1(n_1501),
.B2(n_1477),
.C(n_1495),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1507),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1520),
.B(n_1465),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1518),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1519),
.B(n_1494),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1528),
.B(n_1488),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1519),
.B(n_1495),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1518),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1486),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1505),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1517),
.A2(n_1488),
.B(n_1474),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1506),
.B(n_1470),
.Y(n_1560)
);

OAI31xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1515),
.A2(n_1498),
.A3(n_1454),
.B(n_1453),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1505),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1506),
.B(n_1497),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1509),
.B(n_1497),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1517),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1525),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1516),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1509),
.B(n_1487),
.Y(n_1568)
);

OAI222xp33_ASAP7_75t_L g1569 ( 
.A1(n_1512),
.A2(n_1467),
.B1(n_1471),
.B2(n_1472),
.C1(n_1429),
.C2(n_1439),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1516),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1509),
.B(n_1487),
.Y(n_1571)
);

NOR2xp67_ASAP7_75t_L g1572 ( 
.A(n_1523),
.B(n_1484),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1519),
.B(n_1467),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1515),
.B(n_1492),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1558),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1560),
.B(n_1521),
.Y(n_1576)
);

NOR3xp33_ASAP7_75t_L g1577 ( 
.A(n_1540),
.B(n_1531),
.C(n_1512),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1548),
.B(n_1529),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1541),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1560),
.B(n_1519),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1541),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1558),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1562),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1541),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1538),
.B(n_1521),
.Y(n_1585)
);

OAI211xp5_ASAP7_75t_L g1586 ( 
.A1(n_1561),
.A2(n_1531),
.B(n_1532),
.C(n_1504),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1543),
.Y(n_1587)
);

NAND3x1_ASAP7_75t_L g1588 ( 
.A(n_1559),
.B(n_1504),
.C(n_1530),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1565),
.A2(n_1555),
.B1(n_1554),
.B2(n_1536),
.Y(n_1589)
);

AND2x4_ASAP7_75t_SL g1590 ( 
.A(n_1537),
.B(n_1353),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_1539),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1562),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1567),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1537),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1535),
.B(n_1522),
.Y(n_1595)
);

AOI21xp33_ASAP7_75t_L g1596 ( 
.A1(n_1538),
.A2(n_1532),
.B(n_1513),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1567),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1570),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1536),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1570),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1533),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1533),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1534),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1542),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1542),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1545),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1545),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1534),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1543),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1599),
.B(n_1564),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1590),
.B(n_1534),
.Y(n_1611)
);

CKINVDCx16_ASAP7_75t_R g1612 ( 
.A(n_1589),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1575),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1590),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1576),
.B(n_1564),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1588),
.A2(n_1574),
.B1(n_1544),
.B2(n_1535),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1585),
.B(n_1551),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1585),
.B(n_1551),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1575),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1579),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1582),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1608),
.B(n_1353),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1608),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1578),
.B(n_1574),
.Y(n_1624)
);

INVx3_ASAP7_75t_SL g1625 ( 
.A(n_1603),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1582),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1603),
.B(n_1591),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1576),
.B(n_1568),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1595),
.B(n_1568),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1571),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1601),
.B(n_1547),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1580),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1583),
.Y(n_1633)
);

INVx3_ASAP7_75t_SL g1634 ( 
.A(n_1580),
.Y(n_1634)
);

O2A1O1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1624),
.A2(n_1577),
.B(n_1586),
.C(n_1606),
.Y(n_1635)
);

OAI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1624),
.A2(n_1588),
.B(n_1546),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1623),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1617),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1622),
.A2(n_1580),
.B(n_1546),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1634),
.B(n_1594),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1622),
.A2(n_1594),
.B(n_1555),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1618),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1613),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1634),
.B(n_1594),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1623),
.B(n_1604),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1612),
.A2(n_1555),
.B1(n_1587),
.B2(n_1581),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1619),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.B(n_1544),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1621),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1626),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1616),
.A2(n_1596),
.B1(n_1587),
.B2(n_1584),
.C(n_1581),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1633),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1632),
.A2(n_1572),
.B1(n_1555),
.B2(n_1532),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1638),
.B(n_1628),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1648),
.B(n_1611),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1636),
.B(n_1611),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1637),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1644),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1642),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1644),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1648),
.B(n_1630),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_SL g1665 ( 
.A(n_1661),
.B(n_1640),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1654),
.A2(n_1635),
.B1(n_1651),
.B2(n_1646),
.C(n_1650),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1658),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_SL g1668 ( 
.A(n_1654),
.B(n_1641),
.C(n_1639),
.Y(n_1668)
);

NAND3xp33_ASAP7_75t_L g1669 ( 
.A(n_1659),
.B(n_1627),
.C(n_1643),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1656),
.B(n_1614),
.Y(n_1670)
);

OAI211xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1657),
.A2(n_1653),
.B(n_1627),
.C(n_1649),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1660),
.A2(n_1620),
.B1(n_1584),
.B2(n_1609),
.Y(n_1672)
);

OAI21xp33_ASAP7_75t_L g1673 ( 
.A1(n_1662),
.A2(n_1629),
.B(n_1631),
.Y(n_1673)
);

OAI322xp33_ASAP7_75t_SL g1674 ( 
.A1(n_1663),
.A2(n_1652),
.A3(n_1647),
.B1(n_1605),
.B2(n_1607),
.C1(n_1606),
.C2(n_1602),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1665),
.B(n_1655),
.Y(n_1675)
);

NAND4xp25_ASAP7_75t_L g1676 ( 
.A(n_1670),
.B(n_1664),
.C(n_1607),
.D(n_1602),
.Y(n_1676)
);

AOI222xp33_ASAP7_75t_L g1677 ( 
.A1(n_1666),
.A2(n_1620),
.B1(n_1609),
.B2(n_1579),
.C1(n_1598),
.C2(n_1583),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1673),
.A2(n_1598),
.B1(n_1592),
.B2(n_1597),
.C(n_1593),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1672),
.A2(n_1592),
.B(n_1537),
.C(n_1553),
.Y(n_1679)
);

XNOR2x1_ASAP7_75t_L g1680 ( 
.A(n_1669),
.B(n_1537),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1667),
.A2(n_1674),
.B(n_1600),
.Y(n_1681)
);

OAI21xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1675),
.A2(n_1552),
.B(n_1550),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1680),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1677),
.B(n_1668),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1681),
.B(n_1550),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1676),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1679),
.B(n_1671),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_SL g1688 ( 
.A(n_1678),
.B(n_1553),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1687),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1684),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1682),
.Y(n_1691)
);

AO22x2_ASAP7_75t_L g1692 ( 
.A1(n_1683),
.A2(n_1685),
.B1(n_1686),
.B2(n_1688),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1683),
.A2(n_1553),
.B1(n_1572),
.B2(n_1557),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1689),
.B(n_1557),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1692),
.Y(n_1695)
);

NOR4xp25_ASAP7_75t_L g1696 ( 
.A(n_1691),
.B(n_1552),
.C(n_1556),
.D(n_1549),
.Y(n_1696)
);

NOR3xp33_ASAP7_75t_L g1697 ( 
.A(n_1695),
.B(n_1690),
.C(n_1693),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1697),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1695),
.B(n_1696),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1698),
.Y(n_1700)
);

OAI22xp33_ASAP7_75t_SL g1701 ( 
.A1(n_1700),
.A2(n_1694),
.B1(n_1549),
.B2(n_1543),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1699),
.A2(n_1556),
.B1(n_1563),
.B2(n_1566),
.Y(n_1702)
);

AO22x2_ASAP7_75t_L g1703 ( 
.A1(n_1702),
.A2(n_1566),
.B1(n_1549),
.B2(n_1553),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1701),
.A2(n_1566),
.B(n_1563),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1703),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1705),
.A2(n_1704),
.B1(n_1573),
.B2(n_1504),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1573),
.B(n_1524),
.Y(n_1707)
);

OAI31xp33_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1573),
.A3(n_1569),
.B(n_1530),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1573),
.B1(n_1526),
.B2(n_1522),
.Y(n_1709)
);

AOI211xp5_ASAP7_75t_L g1710 ( 
.A1(n_1709),
.A2(n_1508),
.B(n_1530),
.C(n_1504),
.Y(n_1710)
);


endmodule