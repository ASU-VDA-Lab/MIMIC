module fake_jpeg_11443_n_133 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_0),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_13),
.B1(n_25),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_57),
.B1(n_19),
.B2(n_29),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_17),
.B(n_24),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_52),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_56),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_15),
.B1(n_18),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_58),
.B1(n_17),
.B2(n_19),
.Y(n_61)
);

NOR3xp33_ASAP7_75t_SL g52 ( 
.A(n_29),
.B(n_18),
.C(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_18),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_31),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_20),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_32),
.B1(n_36),
.B2(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_26),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_26),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_36),
.B1(n_41),
.B2(n_33),
.Y(n_70)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_74),
.B(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_14),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_14),
.Y(n_77)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_52),
.A3(n_60),
.B1(n_44),
.B2(n_45),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_81),
.A2(n_86),
.B(n_73),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_48),
.C(n_53),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_87),
.C(n_37),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_58),
.B1(n_43),
.B2(n_52),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_84),
.A2(n_91),
.B1(n_70),
.B2(n_63),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_55),
.B(n_53),
.C(n_37),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_46),
.B1(n_41),
.B2(n_37),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_94),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_65),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_67),
.B1(n_71),
.B2(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_74),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_98),
.B(n_91),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_66),
.B(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_46),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_86),
.C(n_82),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_85),
.B1(n_86),
.B2(n_84),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_97),
.B1(n_101),
.B2(n_93),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_79),
.C(n_86),
.Y(n_107)
);

OAI321xp33_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_80),
.A3(n_11),
.B1(n_46),
.B2(n_41),
.C(n_6),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_115),
.B(n_104),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_98),
.B(n_42),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_2),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_111),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_121),
.C(n_122),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_111),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_104),
.B(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_113),
.B1(n_37),
.B2(n_42),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_41),
.C(n_8),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_3),
.B(n_5),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_129),
.C(n_3),
.Y(n_131)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_9),
.Y(n_133)
);


endmodule