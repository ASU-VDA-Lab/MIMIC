module fake_jpeg_14163_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_5),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_48),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

INVx5_ASAP7_75t_SL g108 ( 
.A(n_47),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_56),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_25),
.B(n_0),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_25),
.C(n_38),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_60),
.B(n_67),
.Y(n_103)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_62),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_32),
.B(n_7),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_14),
.Y(n_88)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_74),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_30),
.Y(n_104)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_76),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_27),
.B1(n_58),
.B2(n_37),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_79),
.A2(n_91),
.B1(n_113),
.B2(n_47),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_83),
.B(n_119),
.C(n_3),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_37),
.B1(n_36),
.B2(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_90),
.B1(n_102),
.B2(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_88),
.B(n_112),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_42),
.A2(n_27),
.B1(n_38),
.B2(n_28),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_35),
.B1(n_26),
.B2(n_33),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_54),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_55),
.A2(n_35),
.B1(n_40),
.B2(n_22),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_54),
.A2(n_40),
.B1(n_22),
.B2(n_16),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_106),
.A2(n_107),
.B1(n_111),
.B2(n_116),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_7),
.B1(n_13),
.B2(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_49),
.B(n_8),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_6),
.B1(n_13),
.B2(n_4),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_115),
.B1(n_81),
.B2(n_123),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_6),
.C(n_10),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_41),
.B(n_12),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_12),
.Y(n_121)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_127),
.B(n_128),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_75),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_108),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_82),
.A2(n_70),
.B1(n_68),
.B2(n_59),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_92),
.B1(n_95),
.B2(n_109),
.Y(n_168)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_63),
.B1(n_62),
.B2(n_65),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_155),
.B1(n_166),
.B2(n_125),
.Y(n_182)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_12),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_137),
.B(n_142),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_61),
.B1(n_44),
.B2(n_64),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_140),
.B1(n_131),
.B2(n_130),
.Y(n_192)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_84),
.A2(n_57),
.B1(n_43),
.B2(n_46),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_1),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_78),
.B(n_14),
.Y(n_142)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_149),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

BUFx16f_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_105),
.Y(n_150)
);

CKINVDCx10_ASAP7_75t_R g151 ( 
.A(n_80),
.Y(n_151)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx6_ASAP7_75t_SL g189 ( 
.A(n_152),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_96),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_156),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_93),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_159),
.Y(n_173)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_85),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_101),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_162),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_94),
.B(n_101),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_164),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_100),
.B(n_77),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_140),
.C(n_151),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_118),
.A2(n_109),
.B1(n_92),
.B2(n_95),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_181),
.B1(n_136),
.B2(n_148),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_93),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_188),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_192),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_126),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_198),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_129),
.A2(n_110),
.B1(n_118),
.B2(n_143),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_199),
.B1(n_169),
.B2(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_132),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_143),
.B(n_140),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_194),
.A2(n_200),
.B(n_178),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_134),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_135),
.B1(n_166),
.B2(n_163),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_140),
.A2(n_157),
.B(n_144),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_145),
.B(n_139),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_203),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_148),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_172),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_154),
.B(n_146),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_209),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_182),
.A2(n_152),
.B1(n_167),
.B2(n_133),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_221),
.B1(n_202),
.B2(n_216),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_159),
.C(n_158),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_175),
.C(n_174),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_213),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_210),
.A2(n_219),
.B(n_222),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_170),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_220),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_218),
.Y(n_244)
);

NAND2x1_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_176),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_190),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_187),
.B(n_176),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_176),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_223),
.B(n_230),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_227),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_172),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_177),
.B(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_233),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_192),
.A2(n_168),
.B1(n_189),
.B2(n_184),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_231),
.A2(n_213),
.B(n_209),
.Y(n_262)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_192),
.B(n_189),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_175),
.B(n_184),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_185),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_235),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_185),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_232),
.A2(n_192),
.B1(n_174),
.B2(n_193),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_257),
.B1(n_212),
.B2(n_223),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_245),
.A2(n_212),
.B(n_218),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_253),
.C(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_197),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_250),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_197),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_230),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_256),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_211),
.C(n_219),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_232),
.A2(n_202),
.B1(n_223),
.B2(n_210),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_202),
.B1(n_212),
.B2(n_206),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_256),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_260),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_222),
.B1(n_208),
.B2(n_205),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_269),
.B1(n_244),
.B2(n_251),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_220),
.C(n_228),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_273),
.C(n_276),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_219),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_278),
.C(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_270),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_274),
.Y(n_291)
);

A2O1A1O1Ixp25_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_217),
.B(n_215),
.C(n_236),
.D(n_235),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_233),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_279),
.Y(n_298)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_249),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_280),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_252),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_246),
.C(n_243),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_244),
.C(n_250),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_284),
.A2(n_258),
.B1(n_243),
.B2(n_248),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_278),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_287),
.B(n_292),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_295),
.B1(n_238),
.B2(n_245),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_257),
.C(n_251),
.Y(n_294)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_294),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_247),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_274),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_299),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_241),
.B1(n_239),
.B2(n_275),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_301),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_290),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_304),
.Y(n_316)
);

AO221x1_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_261),
.B1(n_240),
.B2(n_271),
.C(n_266),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_242),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_251),
.B(n_284),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_310),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_288),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_262),
.B(n_272),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_289),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_287),
.C(n_285),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_318),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_317),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_313),
.A2(n_241),
.B1(n_296),
.B2(n_242),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_294),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_285),
.C(n_292),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_295),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_323),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_326),
.B(n_329),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_319),
.A2(n_308),
.B(n_311),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_308),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_314),
.A2(n_313),
.B1(n_305),
.B2(n_309),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_323),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_332),
.A2(n_334),
.B1(n_330),
.B2(n_245),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_245),
.B1(n_272),
.B2(n_315),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_328),
.A2(n_316),
.B(n_324),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_325),
.B(n_331),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_297),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_336),
.A2(n_286),
.B(n_264),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_334),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_338),
.A2(n_339),
.B(n_333),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_340),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_341),
.C(n_321),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_279),
.B(n_263),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_263),
.Y(n_345)
);


endmodule