module fake_jpeg_23766_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_0),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_20),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_26),
.C(n_31),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_63),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_19),
.B1(n_30),
.B2(n_27),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_68),
.B1(n_27),
.B2(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_45),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_19),
.B1(n_29),
.B2(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_70),
.B(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_71),
.B(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_49),
.B(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_36),
.B1(n_37),
.B2(n_35),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_75),
.A2(n_79),
.B1(n_21),
.B2(n_29),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_34),
.B1(n_39),
.B2(n_38),
.Y(n_79)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_45),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_34),
.C(n_43),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_58),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_45),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_0),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_64),
.B(n_32),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_42),
.B(n_32),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_38),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_1),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_103),
.B(n_117),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_46),
.B1(n_60),
.B2(n_50),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_71),
.B1(n_78),
.B2(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_56),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_102),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_20),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_110),
.B1(n_75),
.B2(n_70),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_24),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_115),
.C(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_16),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_17),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_73),
.B(n_25),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_21),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_74),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_127),
.C(n_137),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_122),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_72),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_128),
.A2(n_135),
.B1(n_115),
.B2(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_101),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_82),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_79),
.B(n_88),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_77),
.B1(n_85),
.B2(n_76),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_95),
.C(n_83),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_100),
.C(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_148),
.Y(n_162)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_144),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_143),
.B1(n_146),
.B2(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_108),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_147),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_107),
.B1(n_109),
.B2(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_107),
.B1(n_115),
.B2(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_108),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_103),
.C(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_98),
.Y(n_168)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_145),
.A2(n_127),
.B(n_136),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_118),
.B(n_123),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_120),
.B1(n_132),
.B2(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_167),
.B1(n_168),
.B2(n_141),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_137),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_165),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_119),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_169),
.A2(n_170),
.B(n_176),
.Y(n_181)
);

AOI321xp33_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_154),
.A3(n_145),
.B1(n_148),
.B2(n_150),
.C(n_151),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_154),
.B(n_146),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_171),
.A2(n_2),
.B(n_6),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_126),
.C(n_143),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_159),
.C(n_166),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_126),
.C(n_125),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_12),
.Y(n_183)
);

OAI321xp33_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_118),
.A3(n_95),
.B1(n_25),
.B2(n_129),
.C(n_8),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_80),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_129),
.B(n_3),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_178),
.A2(n_161),
.B(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_185),
.C(n_7),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_9),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_171),
.A2(n_156),
.B1(n_175),
.B2(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_7),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_81),
.C(n_80),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_2),
.Y(n_188)
);

NAND4xp25_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_175),
.C(n_11),
.D(n_8),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_187),
.A2(n_12),
.B(n_14),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_188),
.B(n_191),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_181),
.B(n_180),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_188),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_189),
.B(n_192),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);


endmodule