module fake_jpeg_29301_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_39),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_63),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_14),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_12),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_53),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_22),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_57),
.Y(n_65)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_28),
.A2(n_0),
.B(n_2),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_62),
.B(n_4),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_0),
.C(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_4),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_29),
.B1(n_35),
.B2(n_26),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_81),
.B1(n_88),
.B2(n_27),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_11),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_73),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_54),
.B1(n_40),
.B2(n_43),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_75),
.A2(n_87),
.B1(n_53),
.B2(n_51),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_38),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_32),
.B1(n_35),
.B2(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_23),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_85),
.B(n_90),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_32),
.B1(n_18),
.B2(n_25),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_32),
.B1(n_26),
.B2(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_39),
.B(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_97),
.Y(n_129)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_94),
.Y(n_107)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_21),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_31),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_101),
.C(n_31),
.Y(n_118)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_117),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx5_ASAP7_75t_SL g153 ( 
.A(n_112),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_64),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_34),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_116),
.Y(n_139)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_121),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_25),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_87),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_126),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_98),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_67),
.A2(n_55),
.B1(n_61),
.B2(n_27),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_88),
.B1(n_81),
.B2(n_75),
.Y(n_136)
);

BUFx4f_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_36),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_127),
.B(n_128),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_36),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_131),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_76),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_158),
.B(n_78),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_87),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_144),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_8),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_89),
.B1(n_95),
.B2(n_101),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_145),
.B1(n_9),
.B2(n_6),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_101),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_131),
.B1(n_109),
.B2(n_105),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_8),
.B(n_9),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_124),
.A2(n_59),
.B1(n_77),
.B2(n_82),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_107),
.B1(n_94),
.B2(n_104),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_34),
.CI(n_21),
.CON(n_152),
.SN(n_152)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_5),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_82),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_157),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_120),
.B(n_113),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_107),
.A2(n_77),
.B(n_93),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_169),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_120),
.C(n_117),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_148),
.C(n_154),
.Y(n_193)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_162),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_164),
.B1(n_134),
.B2(n_133),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_132),
.B1(n_122),
.B2(n_110),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_172),
.Y(n_191)
);

AOI22x1_ASAP7_75t_SL g166 ( 
.A1(n_139),
.A2(n_126),
.B1(n_74),
.B2(n_78),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_177),
.B1(n_150),
.B2(n_135),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_SL g172 ( 
.A(n_150),
.B(n_126),
.C(n_102),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_5),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_174),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_108),
.B(n_7),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_6),
.Y(n_178)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_144),
.B(n_172),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_152),
.C(n_178),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_180),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_152),
.B(n_150),
.C(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_170),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_136),
.B1(n_149),
.B2(n_142),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_192),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_153),
.B1(n_135),
.B2(n_154),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_160),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_143),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_202),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_209),
.C(n_213),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_193),
.C(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_210),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_167),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_176),
.B(n_164),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_221),
.C(n_190),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_195),
.B1(n_188),
.B2(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_212),
.B1(n_201),
.B2(n_207),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_222),
.B(n_184),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_208),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

AOI31xp67_ASAP7_75t_SL g236 ( 
.A1(n_227),
.A2(n_223),
.A3(n_218),
.B(n_182),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_230),
.C(n_221),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_201),
.B(n_217),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_201),
.C(n_190),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_220),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_236),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_234),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_228),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_237),
.A2(n_233),
.B1(n_214),
.B2(n_194),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_177),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_241),
.A2(n_243),
.B1(n_238),
.B2(n_194),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_242),
.A2(n_243),
.B(n_176),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_239),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_245),
.A3(n_179),
.B1(n_162),
.B2(n_171),
.C1(n_175),
.C2(n_163),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_134),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_8),
.Y(n_248)
);


endmodule