module fake_jpeg_11114_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx2_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_57),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_60),
.B(n_74),
.Y(n_164)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_61),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_68),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_21),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_72),
.B(n_93),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_17),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_23),
.B(n_15),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_76),
.B(n_79),
.Y(n_165)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_30),
.B(n_44),
.Y(n_79)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g210 ( 
.A(n_80),
.Y(n_210)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_14),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_83),
.B(n_111),
.Y(n_186)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_39),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_87),
.Y(n_131)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_92),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_48),
.B(n_0),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_96),
.B(n_114),
.Y(n_160)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_97),
.B(n_110),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_104),
.Y(n_154)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_106),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_45),
.B(n_14),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_112),
.B(n_113),
.Y(n_172)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_48),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_119),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_48),
.B(n_1),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_46),
.B(n_13),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_123),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_121),
.B(n_37),
.C(n_2),
.Y(n_203)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_122),
.B(n_5),
.Y(n_208)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_37),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_37),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_79),
.B(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_126),
.B(n_146),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_25),
.B(n_33),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_128),
.B(n_10),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_60),
.B(n_46),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_139),
.B(n_143),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_58),
.A2(n_35),
.B1(n_33),
.B2(n_54),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_141),
.A2(n_152),
.B1(n_153),
.B2(n_177),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_76),
.B(n_35),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_83),
.A2(n_35),
.B(n_33),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_26),
.B1(n_27),
.B2(n_31),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_109),
.A2(n_55),
.B1(n_54),
.B2(n_56),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_55),
.B1(n_51),
.B2(n_50),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_155),
.A2(n_130),
.B1(n_128),
.B2(n_172),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_161),
.B(n_162),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_87),
.B(n_55),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_119),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_163),
.B(n_166),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_67),
.B(n_51),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_71),
.B(n_22),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_171),
.B(n_178),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_110),
.B(n_32),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_173),
.B(n_184),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_63),
.A2(n_25),
.B1(n_50),
.B2(n_22),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_19),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_68),
.A2(n_25),
.B1(n_47),
.B2(n_19),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_182),
.A2(n_190),
.B1(n_204),
.B2(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_69),
.B(n_47),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_124),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_200),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_101),
.A2(n_41),
.B1(n_32),
.B2(n_31),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_70),
.B(n_41),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_192),
.B(n_199),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_73),
.B(n_27),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_75),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_91),
.B(n_26),
.C(n_37),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_5),
.C(n_7),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_98),
.B(n_1),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_202),
.B(n_188),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_100),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_72),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_112),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_8),
.B1(n_10),
.B2(n_204),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_211),
.B(n_240),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_212),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_214),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_215),
.Y(n_295)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_216),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_217),
.A2(n_271),
.B1(n_272),
.B2(n_256),
.Y(n_312)
);

BUFx2_ASAP7_75t_SL g218 ( 
.A(n_210),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_218),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_219),
.A2(n_258),
.B(n_179),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_210),
.Y(n_220)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_150),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_222),
.B(n_232),
.Y(n_283)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_223),
.Y(n_309)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_225),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_227),
.Y(n_316)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_228),
.Y(n_318)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_231),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_165),
.B(n_7),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_233),
.A2(n_267),
.B1(n_248),
.B2(n_246),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_150),
.A2(n_8),
.B1(n_147),
.B2(n_136),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_125),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_238),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_160),
.B(n_8),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_237),
.B(n_247),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_164),
.B(n_186),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_239),
.B(n_263),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_210),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_147),
.A2(n_136),
.B1(n_183),
.B2(n_151),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_243),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_175),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_250),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_131),
.B(n_172),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_246),
.B(n_248),
.C(n_264),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_170),
.B(n_159),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_131),
.B(n_137),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_249),
.Y(n_303)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_134),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_251),
.B(n_255),
.Y(n_314)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_253),
.Y(n_301)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_257),
.B(n_260),
.Y(n_317)
);

AO22x1_ASAP7_75t_L g258 ( 
.A1(n_154),
.A2(n_209),
.B1(n_177),
.B2(n_156),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_137),
.B(n_156),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_261),
.Y(n_300)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

AO22x2_ASAP7_75t_L g261 ( 
.A1(n_132),
.A2(n_158),
.B1(n_197),
.B2(n_134),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_127),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_268),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_127),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_207),
.B(n_182),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_175),
.A2(n_153),
.B(n_140),
.C(n_205),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_266),
.A2(n_144),
.B(n_181),
.C(n_246),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_169),
.A2(n_174),
.B1(n_180),
.B2(n_135),
.Y(n_267)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_133),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_140),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_269),
.B(n_270),
.Y(n_332)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_197),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_195),
.A2(n_135),
.B1(n_180),
.B2(n_174),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_133),
.A2(n_193),
.B1(n_149),
.B2(n_196),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g273 ( 
.A(n_138),
.B(n_179),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_273),
.B(n_277),
.C(n_220),
.Y(n_331)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_196),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_275),
.A2(n_276),
.B1(n_257),
.B2(n_268),
.Y(n_325)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_149),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_168),
.B(n_191),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_279),
.C(n_280),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_132),
.B(n_158),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_138),
.B(n_179),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_193),
.B(n_188),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_181),
.Y(n_305)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_288),
.B(n_215),
.C(n_249),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_247),
.B(n_181),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_289),
.B(n_327),
.C(n_302),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_264),
.A2(n_168),
.B(n_144),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_293),
.A2(n_299),
.B(n_326),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_230),
.A2(n_188),
.B1(n_142),
.B2(n_144),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_294),
.A2(n_308),
.B1(n_323),
.B2(n_313),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_305),
.B(n_331),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_237),
.B(n_219),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_311),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_241),
.A2(n_221),
.B1(n_230),
.B2(n_259),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_219),
.B(n_265),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_256),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_329),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_321),
.A2(n_322),
.B1(n_313),
.B2(n_299),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_229),
.A2(n_258),
.B1(n_248),
.B2(n_211),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_325),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_266),
.A2(n_240),
.B(n_277),
.Y(n_326)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_231),
.B(n_281),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_252),
.B(n_224),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_245),
.B(n_225),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_333),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_223),
.B(n_273),
.Y(n_333)
);

AOI32xp33_ASAP7_75t_L g334 ( 
.A1(n_282),
.A2(n_274),
.A3(n_273),
.B1(n_261),
.B2(n_277),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_334),
.B(n_235),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_285),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_336),
.B(n_357),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_337),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_322),
.A2(n_261),
.B1(n_251),
.B2(n_276),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_338),
.A2(n_346),
.B1(n_348),
.B2(n_358),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_315),
.B(n_213),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_339),
.B(n_345),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_341),
.A2(n_351),
.B(n_352),
.Y(n_379)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_284),
.Y(n_342)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_311),
.B(n_255),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_300),
.A2(n_261),
.B1(n_275),
.B2(n_226),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_347),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_300),
.A2(n_227),
.B1(n_228),
.B2(n_253),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_284),
.Y(n_350)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_326),
.A2(n_293),
.B(n_308),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_307),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_353),
.B(n_365),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

INVx8_ASAP7_75t_L g398 ( 
.A(n_355),
.Y(n_398)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_328),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_321),
.A2(n_304),
.B1(n_286),
.B2(n_330),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_304),
.A2(n_288),
.B(n_298),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_324),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_327),
.A2(n_302),
.B1(n_323),
.B2(n_286),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_303),
.B1(n_301),
.B2(n_319),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_363),
.B(n_324),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_364),
.B(n_309),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_283),
.B(n_332),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_289),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_369),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_297),
.B(n_292),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_368),
.B(n_375),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_306),
.B(n_305),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_302),
.B(n_333),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_319),
.C(n_291),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_371),
.A2(n_301),
.B1(n_318),
.B2(n_316),
.Y(n_395)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_374),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_317),
.A2(n_290),
.B(n_296),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_314),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_292),
.B(n_291),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_397),
.C(n_403),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_378),
.A2(n_400),
.B1(n_408),
.B2(n_338),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_382),
.B(n_391),
.Y(n_409)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_347),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_386),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_368),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_406),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_395),
.A2(n_342),
.B1(n_344),
.B2(n_350),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_320),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_405),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_336),
.B(n_318),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_399),
.B(n_404),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_343),
.A2(n_310),
.B1(n_309),
.B2(n_320),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_361),
.B(n_316),
.C(n_295),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_287),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_374),
.B(n_287),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_375),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_407),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_343),
.A2(n_290),
.B1(n_295),
.B2(n_352),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_414),
.B1(n_415),
.B2(n_387),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_358),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_420),
.C(n_422),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_408),
.A2(n_371),
.B1(n_337),
.B2(n_346),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_402),
.A2(n_354),
.B1(n_348),
.B2(n_345),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_379),
.A2(n_367),
.B(n_341),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_418),
.A2(n_427),
.B(n_430),
.Y(n_455)
);

INVx6_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_419),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_382),
.B(n_394),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_364),
.Y(n_422)
);

OAI32xp33_ASAP7_75t_L g423 ( 
.A1(n_396),
.A2(n_349),
.A3(n_360),
.B1(n_339),
.B2(n_369),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_424),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_403),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_377),
.B(n_370),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_405),
.C(n_404),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_393),
.B(n_360),
.Y(n_426)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_379),
.A2(n_367),
.B(n_351),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_428),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_385),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_429),
.B(n_380),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_395),
.A2(n_362),
.B(n_385),
.Y(n_430)
);

XNOR2x2_ASAP7_75t_SL g431 ( 
.A(n_391),
.B(n_370),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_431),
.B(n_353),
.Y(n_447)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_376),
.Y(n_432)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_433),
.A2(n_434),
.B1(n_378),
.B2(n_381),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_392),
.A2(n_366),
.B1(n_363),
.B2(n_359),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_340),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_436),
.B(n_383),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_439),
.A2(n_415),
.B1(n_424),
.B2(n_427),
.Y(n_462)
);

OAI22x1_ASAP7_75t_L g441 ( 
.A1(n_414),
.A2(n_392),
.B1(n_388),
.B2(n_381),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_441),
.B(n_418),
.Y(n_470)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_442),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_456),
.B1(n_417),
.B2(n_400),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_340),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_450),
.C(n_452),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_413),
.B(n_380),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_417),
.Y(n_464)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_457),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_383),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_453),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_373),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_435),
.B(n_365),
.C(n_387),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_436),
.B(n_356),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_458),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_411),
.A2(n_389),
.B1(n_384),
.B2(n_401),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_412),
.B(n_401),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_426),
.B(n_372),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_389),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_420),
.C(n_409),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_462),
.B(n_463),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_456),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_464),
.B(n_437),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_434),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_471),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_470),
.A2(n_477),
.B(n_455),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_409),
.C(n_431),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_474),
.C(n_478),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_473),
.A2(n_439),
.B1(n_451),
.B2(n_448),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_430),
.C(n_384),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_438),
.B(n_452),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_457),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_455),
.A2(n_423),
.B(n_390),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_390),
.C(n_347),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_410),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_460),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_482),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_473),
.B1(n_474),
.B2(n_472),
.Y(n_500)
);

XNOR2x1_ASAP7_75t_L g482 ( 
.A(n_462),
.B(n_478),
.Y(n_482)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_484),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_476),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_489),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_448),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_491),
.Y(n_502)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_466),
.A2(n_441),
.B1(n_460),
.B2(n_440),
.Y(n_490)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_490),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_447),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_440),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_461),
.C(n_416),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g498 ( 
.A(n_480),
.B(n_477),
.CI(n_470),
.CON(n_498),
.SN(n_498)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_489),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_468),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_499),
.B(n_501),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_500),
.A2(n_416),
.B1(n_419),
.B2(n_407),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_469),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_482),
.A2(n_492),
.B1(n_469),
.B2(n_461),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_503),
.A2(n_386),
.B1(n_398),
.B2(n_505),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_505),
.B(n_493),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_492),
.C(n_487),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g519 ( 
.A(n_506),
.B(n_508),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_487),
.C(n_491),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_SL g515 ( 
.A(n_509),
.B(n_511),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_510),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_496),
.B(n_355),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_512),
.B(n_514),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_495),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_504),
.A2(n_386),
.B1(n_398),
.B2(n_497),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_507),
.B(n_494),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_518),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_520),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_509),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_503),
.C(n_502),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_506),
.B(n_513),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_523),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_519),
.B(n_514),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g527 ( 
.A1(n_524),
.A2(n_517),
.B(n_516),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_525),
.B(n_502),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_527),
.B(n_529),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_526),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_522),
.B(n_516),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_530),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_522),
.Y(n_534)
);


endmodule