module fake_jpeg_2583_n_226 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_22),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_15),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_15),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

CKINVDCx6p67_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_87),
.Y(n_99)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_66),
.B1(n_73),
.B2(n_55),
.Y(n_91)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_74),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_77),
.B1(n_71),
.B2(n_55),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_94),
.B1(n_81),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_73),
.B1(n_66),
.B2(n_71),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_73),
.B1(n_67),
.B2(n_78),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_79),
.B1(n_57),
.B2(n_54),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_74),
.B1(n_76),
.B2(n_72),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_76),
.B1(n_72),
.B2(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_101),
.B1(n_81),
.B2(n_60),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_70),
.B1(n_69),
.B2(n_59),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_105),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_104),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_63),
.C(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_64),
.Y(n_105)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_108),
.B(n_88),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_14),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_113),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_60),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_2),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_115),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_120),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_88),
.B1(n_9),
.B2(n_10),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_11),
.B(n_12),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_29),
.A3(n_51),
.B1(n_47),
.B2(n_43),
.Y(n_119)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_32),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_6),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_28),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_128),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_25),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_140),
.B1(n_107),
.B2(n_24),
.Y(n_150)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_134),
.B(n_130),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_13),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_136),
.B(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_14),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_17),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_145),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_19),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_149),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_150),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_20),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_152),
.B(n_163),
.Y(n_182)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_161),
.Y(n_179)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_21),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_153),
.B(n_144),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_35),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_139),
.B(n_34),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_166),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_170),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_125),
.C(n_39),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_178),
.C(n_185),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_154),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_175),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_53),
.C(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_184),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_156),
.B(n_164),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_160),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_185),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_193),
.Y(n_201)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_196),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_168),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_177),
.B1(n_171),
.B2(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_190),
.B1(n_193),
.B2(n_188),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_179),
.C(n_172),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_207),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_180),
.C(n_173),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_205),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_209),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_189),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_187),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_210),
.B(n_201),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_214),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_222),
.B(n_216),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_216),
.C(n_213),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_224),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_170),
.Y(n_226)
);


endmodule