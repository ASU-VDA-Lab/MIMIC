module fake_jpeg_25786_n_19 (n_3, n_2, n_1, n_0, n_4, n_19);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_19;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_18;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g5 ( 
.A(n_2),
.B(n_0),
.Y(n_5)
);

OAI22xp33_ASAP7_75t_L g6 ( 
.A1(n_4),
.A2(n_2),
.B1(n_3),
.B2(n_1),
.Y(n_6)
);

INVx13_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

AOI22xp33_ASAP7_75t_SL g8 ( 
.A1(n_1),
.A2(n_3),
.B1(n_2),
.B2(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_9),
.B(n_10),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_0),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_1),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_11),
.Y(n_17)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_9),
.CI(n_14),
.CON(n_16),
.SN(n_16)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_17),
.B(n_15),
.Y(n_18)
);

AOI322xp5_ASAP7_75t_L g19 ( 
.A1(n_18),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_16),
.C1(n_17),
.C2(n_13),
.Y(n_19)
);


endmodule