module fake_jpeg_3099_n_534 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_378;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_59),
.Y(n_101)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_50),
.Y(n_147)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_53),
.Y(n_113)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_56),
.Y(n_162)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_58),
.B(n_60),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_69),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_15),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_6),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_76),
.B(n_36),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_98),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_99),
.B(n_42),
.Y(n_141)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_100),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_109),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_43),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_18),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_121),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_53),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_18),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_132),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_92),
.Y(n_132)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_15),
.B1(n_42),
.B2(n_43),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_152),
.B1(n_33),
.B2(n_29),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_51),
.B(n_46),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_138),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_38),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_91),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_66),
.B(n_46),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_150),
.B(n_155),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_48),
.A2(n_45),
.B1(n_40),
.B2(n_36),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_71),
.B(n_45),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_159),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_75),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_164),
.B(n_177),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_62),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_165),
.Y(n_247)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_114),
.A2(n_40),
.B1(n_33),
.B2(n_29),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_170),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_172),
.A2(n_139),
.B1(n_115),
.B2(n_126),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_28),
.B1(n_85),
.B2(n_63),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_173),
.A2(n_197),
.B1(n_134),
.B2(n_84),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_117),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_174),
.B(n_188),
.Y(n_225)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_127),
.B(n_28),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g180 ( 
.A(n_101),
.Y(n_180)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_109),
.B(n_50),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g243 ( 
.A(n_183),
.B(n_201),
.Y(n_243)
);

CKINVDCx12_ASAP7_75t_R g184 ( 
.A(n_107),
.Y(n_184)
);

INVxp33_ASAP7_75t_SL g223 ( 
.A(n_184),
.Y(n_223)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

OR2x4_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_79),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_187),
.A2(n_183),
.B(n_165),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_103),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_191),
.Y(n_234)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_111),
.B(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_192),
.B(n_194),
.Y(n_232)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_195),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_0),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_198),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_146),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_147),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_202),
.Y(n_215)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_200),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_94),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_120),
.A2(n_88),
.B1(n_73),
.B2(n_82),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_203),
.A2(n_205),
.B1(n_161),
.B2(n_160),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_77),
.B1(n_68),
.B2(n_65),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_209),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_129),
.B(n_0),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_116),
.Y(n_213)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_112),
.B(n_55),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_210),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_211),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_213),
.B(n_216),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_162),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_187),
.A2(n_130),
.B1(n_123),
.B2(n_142),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_229),
.A2(n_238),
.B1(n_203),
.B2(n_131),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_176),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_235),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_168),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_237),
.A2(n_201),
.B(n_188),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_165),
.A2(n_102),
.B1(n_64),
.B2(n_81),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_183),
.A2(n_126),
.B(n_142),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_164),
.B(n_201),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_248),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_164),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_249),
.Y(n_305)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_194),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_253),
.B(n_261),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_204),
.B1(n_179),
.B2(n_163),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_258),
.A2(n_262),
.B1(n_246),
.B2(n_247),
.Y(n_280)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_260),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_174),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_208),
.B1(n_207),
.B2(n_199),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_213),
.B(n_208),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_272),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_248),
.B1(n_227),
.B2(n_228),
.Y(n_282)
);

AO21x1_ASAP7_75t_L g306 ( 
.A1(n_267),
.A2(n_222),
.B(n_239),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_177),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_197),
.B1(n_206),
.B2(n_190),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_277),
.B(n_171),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_216),
.B(n_209),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_276),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_236),
.B(n_196),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_271),
.B(n_278),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_240),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_243),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_275),
.Y(n_297)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_198),
.Y(n_276)
);

O2A1O1Ixp33_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_182),
.B(n_202),
.C(n_181),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_186),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_224),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_283),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_261),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_220),
.B(n_215),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_285),
.A2(n_286),
.B(n_306),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_254),
.A2(n_246),
.B1(n_248),
.B2(n_238),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_289),
.A2(n_299),
.B1(n_309),
.B2(n_278),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_254),
.A2(n_248),
.B1(n_225),
.B2(n_226),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_290),
.Y(n_342)
);

AO22x1_ASAP7_75t_SL g293 ( 
.A1(n_249),
.A2(n_243),
.B1(n_226),
.B2(n_218),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_302),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_243),
.C(n_234),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_294),
.B(n_295),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_234),
.C(n_218),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_233),
.B1(n_222),
.B2(n_211),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_256),
.Y(n_300)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_300),
.Y(n_317)
);

OAI32xp33_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_224),
.A3(n_230),
.B1(n_193),
.B2(n_195),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_264),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_256),
.Y(n_304)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_197),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_SL g323 ( 
.A1(n_308),
.A2(n_267),
.B(n_279),
.C(n_272),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_249),
.A2(n_230),
.B1(n_143),
.B2(n_156),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_276),
.Y(n_310)
);

INVx13_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_263),
.B(n_223),
.C(n_130),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_255),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_259),
.B1(n_250),
.B2(n_249),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_313),
.A2(n_316),
.B1(n_325),
.B2(n_331),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_300),
.A2(n_250),
.B1(n_249),
.B2(n_275),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_327),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_319),
.A2(n_292),
.B1(n_298),
.B2(n_293),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_294),
.Y(n_345)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_323),
.A2(n_305),
.B(n_306),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_271),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_324),
.B(n_340),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_252),
.B1(n_250),
.B2(n_266),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_287),
.B(n_253),
.Y(n_326)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_281),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_287),
.B(n_270),
.Y(n_329)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_329),
.Y(n_361)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_308),
.A2(n_268),
.B1(n_251),
.B2(n_265),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_308),
.A2(n_268),
.B1(n_251),
.B2(n_258),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_333),
.A2(n_343),
.B1(n_299),
.B2(n_297),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_301),
.A2(n_269),
.B(n_277),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_335),
.A2(n_344),
.B(n_309),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_306),
.Y(n_336)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_303),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_337),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_212),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_285),
.Y(n_351)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_242),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_280),
.A2(n_260),
.B1(n_277),
.B2(n_244),
.Y(n_343)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_293),
.A2(n_260),
.B(n_219),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_345),
.B(n_329),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_346),
.A2(n_349),
.B1(n_374),
.B2(n_344),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_347),
.A2(n_359),
.B(n_360),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_333),
.A2(n_288),
.B1(n_286),
.B2(n_298),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_295),
.C(n_297),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_373),
.C(n_337),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_351),
.A2(n_363),
.B1(n_375),
.B2(n_336),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_328),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_352),
.B(n_367),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_291),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_354),
.B(n_239),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_342),
.A2(n_305),
.B1(n_292),
.B2(n_293),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_326),
.B(n_212),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_318),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_372),
.Y(n_379)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_369),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_341),
.B(n_212),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_378),
.Y(n_385)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_371),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_320),
.B(n_311),
.C(n_316),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_331),
.A2(n_284),
.B1(n_307),
.B2(n_302),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_319),
.A2(n_315),
.B1(n_325),
.B2(n_314),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_332),
.Y(n_376)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_376),
.Y(n_391)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_327),
.B(n_307),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_381),
.B(n_398),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_313),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_387),
.Y(n_413)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_338),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_384),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_358),
.C(n_364),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_314),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_388),
.A2(n_404),
.B1(n_362),
.B2(n_376),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_390),
.A2(n_156),
.B1(n_143),
.B2(n_128),
.Y(n_432)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_392),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_334),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_401),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_347),
.A2(n_344),
.B(n_335),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_394),
.A2(n_365),
.B(n_366),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_357),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_395),
.B(n_407),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_343),
.Y(n_396)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_396),
.Y(n_416)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_397),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_361),
.B(n_323),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_323),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_361),
.B(n_323),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_403),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_323),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_346),
.A2(n_328),
.B1(n_322),
.B2(n_317),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_322),
.B1(n_317),
.B2(n_244),
.Y(n_405)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_406),
.Y(n_433)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_356),
.A2(n_185),
.B1(n_219),
.B2(n_242),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_408),
.A2(n_374),
.B1(n_349),
.B2(n_371),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_358),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_409),
.B(n_417),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_411),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_414),
.B(n_423),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_415),
.A2(n_432),
.B1(n_404),
.B2(n_399),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_387),
.C(n_393),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_369),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_421),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_364),
.C(n_362),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_363),
.C(n_348),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_368),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_425),
.B(n_166),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_388),
.A2(n_365),
.B1(n_360),
.B2(n_377),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_178),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_428),
.A2(n_189),
.B(n_175),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_379),
.B(n_366),
.C(n_239),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_429),
.B(n_430),
.C(n_394),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_379),
.B(n_170),
.C(n_191),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_396),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_434),
.A2(n_106),
.B1(n_131),
.B2(n_178),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_403),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_440),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_431),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_444),
.B1(n_447),
.B2(n_454),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_437),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_439),
.A2(n_446),
.B1(n_136),
.B2(n_102),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_389),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_389),
.C(n_401),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_445),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_428),
.A2(n_384),
.B(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_443),
.Y(n_469)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_402),
.C(n_391),
.Y(n_445)
);

AOI321xp33_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_383),
.A3(n_380),
.B1(n_178),
.B2(n_122),
.C(n_133),
.Y(n_446)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_171),
.C(n_123),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_452),
.C(n_412),
.Y(n_459)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_115),
.C(n_128),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_200),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_122),
.Y(n_471)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_433),
.Y(n_454)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_455),
.Y(n_475)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_457),
.B(n_456),
.Y(n_458)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_458),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_471),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_451),
.B(n_423),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_461),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_422),
.C(n_427),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_441),
.A2(n_427),
.B1(n_416),
.B2(n_424),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_443),
.B1(n_439),
.B2(n_447),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_422),
.C(n_411),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_465),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_426),
.C(n_412),
.Y(n_465)
);

FAx1_ASAP7_75t_SL g467 ( 
.A(n_445),
.B(n_430),
.CI(n_432),
.CON(n_467),
.SN(n_467)
);

MAJx2_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_157),
.C(n_124),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_106),
.C(n_169),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_435),
.C(n_453),
.Y(n_482)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_476),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_441),
.B(n_12),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_477),
.B(n_11),
.Y(n_489)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_469),
.A2(n_448),
.B(n_449),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_483),
.A2(n_3),
.B(n_4),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_452),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_487),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_462),
.C(n_464),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_446),
.B(n_133),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_488),
.A2(n_494),
.B1(n_471),
.B2(n_467),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_490),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_462),
.B(n_161),
.C(n_160),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_474),
.B(n_157),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_491),
.B(n_493),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_492),
.B(n_490),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_124),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_476),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_486),
.A2(n_470),
.B1(n_475),
.B2(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_459),
.C(n_472),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_501),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_500),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_SL g503 ( 
.A(n_478),
.B(n_485),
.C(n_481),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_503),
.B(n_4),
.C(n_9),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_481),
.B(n_467),
.C(n_146),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_504),
.B(n_506),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_479),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_483),
.A2(n_5),
.B(n_1),
.C(n_3),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_507),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_508),
.B(n_0),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_511),
.A2(n_516),
.B(n_517),
.Y(n_522)
);

OA21x2_ASAP7_75t_SL g513 ( 
.A1(n_497),
.A2(n_492),
.B(n_482),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_504),
.C(n_498),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_515),
.A2(n_9),
.B(n_10),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_496),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_499),
.B(n_9),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_512),
.A2(n_495),
.B(n_508),
.Y(n_519)
);

A2O1A1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_519),
.A2(n_524),
.B(n_510),
.C(n_513),
.Y(n_527)
);

AOI21xp33_ASAP7_75t_L g520 ( 
.A1(n_509),
.A2(n_507),
.B(n_502),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_521),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_523),
.B(n_10),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_514),
.A2(n_10),
.B(n_11),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_522),
.B(n_518),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_525),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_527),
.B(n_528),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_526),
.C(n_13),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_SL g532 ( 
.A1(n_531),
.A2(n_529),
.B1(n_13),
.B2(n_0),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_13),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_13),
.Y(n_534)
);


endmodule