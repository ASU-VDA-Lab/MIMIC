module real_jpeg_23006_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_288;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_249;
wire n_286;
wire n_292;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_271;
wire n_131;
wire n_47;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_173;
wire n_40;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_306;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_80;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_1),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_1),
.B(n_78),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_167),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_1),
.A2(n_28),
.B(n_48),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_1),
.B(n_121),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_1),
.A2(n_91),
.B1(n_255),
.B2(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_1),
.A2(n_61),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_36),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_2),
.A2(n_36),
.B1(n_61),
.B2(n_62),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_2),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_5),
.A2(n_68),
.B1(n_70),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_176),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_176),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_176),
.Y(n_255)
);

INVx8_ASAP7_75t_SL g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_53),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_7),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_27),
.B1(n_61),
.B2(n_62),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_8),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_8),
.A2(n_27),
.B1(n_70),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_44),
.B1(n_61),
.B2(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_44),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_10),
.A2(n_68),
.B1(n_70),
.B2(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_73),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_73),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_73),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_13),
.A2(n_66),
.B1(n_70),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_116),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_116),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_116),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_15),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_150),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_148),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_20),
.B(n_122),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_89),
.C(n_102),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_21),
.B(n_89),
.CI(n_102),
.CON(n_179),
.SN(n_179)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_54),
.B2(n_88),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_22),
.B(n_55),
.C(n_79),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_24),
.B(n_39),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_25),
.A2(n_172),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_26),
.B(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_30),
.B1(n_48),
.B2(n_50),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_30),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_31),
.A2(n_107),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_31),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_34),
.A2(n_91),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_38),
.B(n_167),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_40),
.A2(n_51),
.B(n_112),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_41),
.A2(n_42),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_41),
.B(n_82),
.Y(n_278)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_42),
.A2(n_50),
.B(n_167),
.C(n_231),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_42),
.A2(n_61),
.A3(n_81),
.B1(n_271),
.B2(n_278),
.Y(n_277)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_45),
.A2(n_52),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_45),
.A2(n_51),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_45),
.A2(n_129),
.B(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_46),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_46),
.A2(n_99),
.B(n_130),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_46),
.A2(n_131),
.B1(n_229),
.B2(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_46),
.A2(n_131),
.B1(n_237),
.B2(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_51),
.B(n_167),
.Y(n_253)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_79),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_69),
.B(n_74),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_56),
.A2(n_57),
.B1(n_69),
.B2(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_56),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_56),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_65),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_58),
.A2(n_62),
.A3(n_71),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_59),
.B(n_61),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_61),
.A2(n_62),
.B1(n_81),
.B2(n_82),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_62),
.B(n_167),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_70),
.A2(n_166),
.B(n_167),
.Y(n_191)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_75),
.Y(n_139)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_76),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_78),
.B(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_78),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_78),
.A2(n_175),
.B1(n_177),
.B2(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_84),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_80),
.B(n_119),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_80),
.A2(n_118),
.B1(n_211),
.B2(n_269),
.Y(n_268)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_85),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_85),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_85),
.A2(n_121),
.B1(n_162),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_85),
.A2(n_121),
.B1(n_193),
.B2(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_96),
.B1(n_97),
.B2(n_101),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_97),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_101),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B(n_95),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_91),
.A2(n_92),
.B1(n_245),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_91),
.A2(n_95),
.B(n_108),
.Y(n_279)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_94),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_100),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.C(n_117),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_104),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_111),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_105),
.B(n_111),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_114),
.B(n_117),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_147),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_133),
.B1(n_145),
.B2(n_146),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_128),
.B(n_132),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_144),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_180),
.B(n_306),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_179),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_152),
.B(n_179),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.C(n_159),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_159),
.A2(n_160),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_174),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_174),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_169),
.B1(n_170),
.B2(n_206),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_179),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_218),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_198),
.B(n_217),
.Y(n_182)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_183),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_195),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_184),
.B(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_194),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_186),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_194),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.C(n_192),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_192),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_199),
.B(n_202),
.Y(n_305)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.C(n_207),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_203),
.B(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_209),
.B(n_288),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_304),
.C(n_305),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_298),
.B(n_303),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_283),
.B(n_297),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_264),
.B(n_282),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_241),
.B(n_263),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_232),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_224),
.B(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_225),
.A2(n_226),
.B1(n_230),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_238),
.C(n_239),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_236),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_240),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_251),
.B(n_262),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_249),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_243),
.B(n_249),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_256),
.B(n_261),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_254),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_266),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_276),
.B1(n_280),
.B2(n_281),
.Y(n_266)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_275),
.C(n_280),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_279),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_284),
.B(n_285),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_290),
.B2(n_291),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_293),
.C(n_295),
.Y(n_299)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);


endmodule