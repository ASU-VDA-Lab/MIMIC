module real_aes_15851_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_1787;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_1712;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_1802;
wire n_397;
wire n_727;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1777;
wire n_444;
wire n_1200;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1280;
wire n_729;
wire n_394;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_1705;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_0), .A2(n_57), .B1(n_575), .B2(n_576), .Y(n_574) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_0), .Y(n_606) );
INVx1_ASAP7_75t_L g783 ( .A(n_1), .Y(n_783) );
XNOR2xp5_ASAP7_75t_L g1120 ( .A(n_2), .B(n_1121), .Y(n_1120) );
INVx1_ASAP7_75t_L g1775 ( .A(n_3), .Y(n_1775) );
INVx1_ASAP7_75t_L g401 ( .A(n_4), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_4), .B(n_362), .Y(n_467) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_4), .B(n_366), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_4), .B(n_250), .Y(n_1673) );
CKINVDCx5p33_ASAP7_75t_R g640 ( .A(n_5), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_6), .A2(n_254), .B1(n_963), .B2(n_1387), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_6), .A2(n_195), .B1(n_939), .B2(n_953), .Y(n_1403) );
INVx1_ASAP7_75t_L g469 ( .A(n_7), .Y(n_469) );
INVx1_ASAP7_75t_L g1698 ( .A(n_8), .Y(n_1698) );
OAI22xp5_ASAP7_75t_L g1711 ( .A1(n_8), .A2(n_81), .B1(n_1712), .B2(n_1717), .Y(n_1711) );
INVx1_ASAP7_75t_L g1350 ( .A(n_9), .Y(n_1350) );
OAI22xp33_ASAP7_75t_SL g672 ( .A1(n_10), .A2(n_331), .B1(n_585), .B2(n_673), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_10), .A2(n_176), .B1(n_446), .B2(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g1379 ( .A(n_11), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_11), .A2(n_254), .B1(n_953), .B2(n_1173), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g1351 ( .A1(n_12), .A2(n_147), .B1(n_354), .B2(n_363), .Y(n_1351) );
OAI22xp5_ASAP7_75t_L g1353 ( .A1(n_12), .A2(n_147), .B1(n_690), .B2(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g793 ( .A(n_13), .Y(n_793) );
INVx1_ASAP7_75t_L g1661 ( .A(n_14), .Y(n_1661) );
INVx1_ASAP7_75t_L g545 ( .A(n_15), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_16), .A2(n_42), .B1(n_775), .B2(n_777), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_16), .A2(n_42), .B1(n_354), .B2(n_363), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_17), .Y(n_701) );
INVx2_ASAP7_75t_L g412 ( .A(n_18), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g1486 ( .A1(n_19), .A2(n_22), .B1(n_1432), .B2(n_1440), .Y(n_1486) );
INVx1_ASAP7_75t_L g1189 ( .A(n_20), .Y(n_1189) );
INVx1_ASAP7_75t_L g1187 ( .A(n_21), .Y(n_1187) );
XNOR2xp5_ASAP7_75t_L g532 ( .A(n_22), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g1247 ( .A(n_23), .Y(n_1247) );
INVx1_ASAP7_75t_L g1300 ( .A(n_24), .Y(n_1300) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_25), .A2(n_175), .B1(n_945), .B2(n_948), .Y(n_944) );
AOI22xp33_ASAP7_75t_SL g972 ( .A1(n_25), .A2(n_133), .B1(n_973), .B2(n_974), .Y(n_972) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_26), .A2(n_87), .B1(n_808), .B2(n_956), .C(n_1176), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_26), .A2(n_40), .B1(n_974), .B2(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g835 ( .A(n_27), .Y(n_835) );
AOI22xp33_ASAP7_75t_SL g1326 ( .A1(n_28), .A2(n_158), .B1(n_603), .B2(n_963), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_28), .A2(n_203), .B1(n_516), .B2(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g1078 ( .A(n_29), .Y(n_1078) );
INVx1_ASAP7_75t_L g986 ( .A(n_30), .Y(n_986) );
OAI221xp5_ASAP7_75t_L g1786 ( .A1(n_31), .A2(n_86), .B1(n_409), .B2(n_690), .C(n_1787), .Y(n_1786) );
INVx1_ASAP7_75t_L g1799 ( .A(n_31), .Y(n_1799) );
HB1xp67_ASAP7_75t_L g1420 ( .A(n_32), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_32), .B(n_1418), .Y(n_1433) );
AOI22xp33_ASAP7_75t_L g1566 ( .A1(n_33), .A2(n_190), .B1(n_1440), .B2(n_1461), .Y(n_1566) );
INVx1_ASAP7_75t_L g1134 ( .A(n_34), .Y(n_1134) );
OAI22xp33_ASAP7_75t_SL g389 ( .A1(n_35), .A2(n_163), .B1(n_390), .B2(n_392), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_35), .A2(n_163), .B1(n_408), .B2(n_417), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g929 ( .A1(n_36), .A2(n_201), .B1(n_330), .B2(n_609), .C1(n_610), .C2(n_930), .Y(n_929) );
OAI222xp33_ASAP7_75t_L g980 ( .A1(n_36), .A2(n_201), .B1(n_330), .B2(n_483), .C1(n_575), .C2(n_576), .Y(n_980) );
CKINVDCx5p33_ASAP7_75t_R g1038 ( .A(n_37), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_38), .A2(n_181), .B1(n_844), .B2(n_845), .Y(n_843) );
OAI22xp33_ASAP7_75t_L g855 ( .A1(n_38), .A2(n_181), .B1(n_354), .B2(n_856), .Y(n_855) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_39), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_39), .A2(n_57), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g1177 ( .A1(n_40), .A2(n_70), .B1(n_808), .B2(n_956), .C(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1289 ( .A(n_41), .Y(n_1289) );
INVx1_ASAP7_75t_L g1104 ( .A(n_43), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_43), .A2(n_336), .B1(n_759), .B2(n_1112), .Y(n_1111) );
INVx1_ASAP7_75t_L g890 ( .A(n_44), .Y(n_890) );
INVx1_ASAP7_75t_L g852 ( .A(n_45), .Y(n_852) );
OAI211xp5_ASAP7_75t_L g857 ( .A1(n_45), .A2(n_375), .B(n_750), .C(n_858), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g1459 ( .A1(n_46), .A2(n_207), .B1(n_1432), .B2(n_1437), .Y(n_1459) );
AOI22xp5_ASAP7_75t_L g1447 ( .A1(n_47), .A2(n_325), .B1(n_1440), .B2(n_1448), .Y(n_1447) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_48), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g1377 ( .A(n_49), .Y(n_1377) );
INVx1_ASAP7_75t_L g1137 ( .A(n_50), .Y(n_1137) );
AOI22xp33_ASAP7_75t_SL g1317 ( .A1(n_51), .A2(n_203), .B1(n_1318), .B2(n_1321), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_51), .A2(n_158), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
INVx1_ASAP7_75t_L g1181 ( .A(n_52), .Y(n_1181) );
AOI22xp33_ASAP7_75t_SL g1211 ( .A1(n_52), .A2(n_258), .B1(n_963), .B2(n_1212), .Y(n_1211) );
INVx1_ASAP7_75t_L g1778 ( .A(n_53), .Y(n_1778) );
AOI22xp5_ASAP7_75t_L g1460 ( .A1(n_54), .A2(n_302), .B1(n_1440), .B2(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1071 ( .A(n_55), .Y(n_1071) );
XNOR2xp5_ASAP7_75t_L g746 ( .A(n_56), .B(n_747), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g1466 ( .A1(n_56), .A2(n_119), .B1(n_1432), .B2(n_1437), .Y(n_1466) );
INVx1_ASAP7_75t_L g1254 ( .A(n_58), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_59), .B(n_438), .Y(n_1789) );
INVxp67_ASAP7_75t_SL g1796 ( .A(n_59), .Y(n_1796) );
OAI211xp5_ASAP7_75t_SL g868 ( .A1(n_60), .A2(n_688), .B(n_768), .C(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g880 ( .A(n_60), .Y(n_880) );
OAI211xp5_ASAP7_75t_L g1271 ( .A1(n_61), .A2(n_431), .B(n_1272), .C(n_1274), .Y(n_1271) );
INVx1_ASAP7_75t_L g1281 ( .A(n_61), .Y(n_1281) );
OAI211xp5_ASAP7_75t_L g660 ( .A1(n_62), .A2(n_661), .B(n_662), .C(n_666), .Y(n_660) );
INVx1_ASAP7_75t_L g687 ( .A(n_62), .Y(n_687) );
INVx1_ASAP7_75t_L g833 ( .A(n_63), .Y(n_833) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_64), .A2(n_170), .B1(n_408), .B2(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_64), .A2(n_170), .B1(n_390), .B2(n_882), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_65), .Y(n_629) );
INVx1_ASAP7_75t_L g578 ( .A(n_66), .Y(n_578) );
OAI222xp33_ASAP7_75t_L g1366 ( .A1(n_67), .A2(n_178), .B1(n_671), .B2(n_674), .C1(n_1367), .C2(n_1368), .Y(n_1366) );
OAI222xp33_ASAP7_75t_L g1393 ( .A1(n_67), .A2(n_178), .B1(n_222), .B2(n_1394), .C1(n_1395), .C2(n_1396), .Y(n_1393) );
XOR2xp5_ASAP7_75t_L g1761 ( .A(n_68), .B(n_1762), .Y(n_1761) );
OAI22xp33_ASAP7_75t_L g1792 ( .A1(n_69), .A2(n_182), .B1(n_446), .B2(n_928), .Y(n_1792) );
INVxp67_ASAP7_75t_SL g1798 ( .A(n_69), .Y(n_1798) );
AOI22xp33_ASAP7_75t_L g1213 ( .A1(n_70), .A2(n_87), .B1(n_1214), .B2(n_1216), .Y(n_1213) );
INVx1_ASAP7_75t_L g1345 ( .A(n_71), .Y(n_1345) );
INVx1_ASAP7_75t_L g1299 ( .A(n_72), .Y(n_1299) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_73), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_74), .A2(n_167), .B1(n_408), .B2(n_417), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_74), .A2(n_167), .B1(n_392), .B2(n_759), .Y(n_860) );
INVx1_ASAP7_75t_L g583 ( .A(n_75), .Y(n_583) );
INVx1_ASAP7_75t_L g1295 ( .A(n_76), .Y(n_1295) );
INVx1_ASAP7_75t_L g900 ( .A(n_77), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_78), .Y(n_1000) );
INVx1_ASAP7_75t_L g568 ( .A(n_79), .Y(n_568) );
INVx1_ASAP7_75t_L g757 ( .A(n_80), .Y(n_757) );
OAI211xp5_ASAP7_75t_L g767 ( .A1(n_80), .A2(n_688), .B(n_768), .C(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g1680 ( .A(n_81), .Y(n_1680) );
INVx1_ASAP7_75t_L g1777 ( .A(n_82), .Y(n_1777) );
INVx1_ASAP7_75t_L g502 ( .A(n_83), .Y(n_502) );
INVx1_ASAP7_75t_L g1131 ( .A(n_84), .Y(n_1131) );
XNOR2xp5_ASAP7_75t_L g1026 ( .A(n_85), .B(n_1027), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g1451 ( .A1(n_85), .A2(n_335), .B1(n_1432), .B2(n_1437), .Y(n_1451) );
OAI22xp33_ASAP7_75t_L g1801 ( .A1(n_86), .A2(n_182), .B1(n_673), .B2(n_734), .Y(n_1801) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_88), .A2(n_192), .B1(n_409), .B2(n_446), .Y(n_1184) );
INVx1_ASAP7_75t_L g1195 ( .A(n_88), .Y(n_1195) );
INVx1_ASAP7_75t_L g1017 ( .A(n_89), .Y(n_1017) );
OAI211xp5_ASAP7_75t_L g1022 ( .A1(n_89), .A2(n_431), .B(n_511), .C(n_1023), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_90), .A2(n_266), .B1(n_673), .B2(n_726), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_90), .A2(n_127), .B1(n_419), .B2(n_446), .Y(n_737) );
INVx1_ASAP7_75t_L g899 ( .A(n_91), .Y(n_899) );
INVx1_ASAP7_75t_L g1791 ( .A(n_92), .Y(n_1791) );
CKINVDCx5p33_ASAP7_75t_R g729 ( .A(n_93), .Y(n_729) );
INVx1_ASAP7_75t_L g1276 ( .A(n_94), .Y(n_1276) );
OAI211xp5_ASAP7_75t_L g1279 ( .A1(n_94), .A2(n_753), .B(n_1090), .C(n_1280), .Y(n_1279) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_95), .Y(n_698) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_96), .Y(n_627) );
INVx1_ASAP7_75t_L g1190 ( .A(n_97), .Y(n_1190) );
AOI22xp33_ASAP7_75t_SL g1327 ( .A1(n_98), .A2(n_341), .B1(n_1318), .B2(n_1321), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_98), .A2(n_99), .B1(n_1333), .B2(n_1336), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_99), .A2(n_311), .B1(n_963), .B2(n_1323), .Y(n_1322) );
AOI22xp5_ASAP7_75t_SL g1452 ( .A1(n_100), .A2(n_218), .B1(n_1440), .B2(n_1448), .Y(n_1452) );
XOR2xp5_ASAP7_75t_L g622 ( .A(n_101), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g1135 ( .A(n_102), .Y(n_1135) );
INVx1_ASAP7_75t_L g547 ( .A(n_103), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_103), .A2(n_288), .B1(n_596), .B2(n_603), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_104), .Y(n_1042) );
INVx1_ASAP7_75t_L g1294 ( .A(n_105), .Y(n_1294) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_106), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g1158 ( .A1(n_107), .A2(n_139), .B1(n_363), .B2(n_673), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_107), .A2(n_125), .B1(n_408), .B2(n_446), .Y(n_1160) );
INVx1_ASAP7_75t_L g1127 ( .A(n_108), .Y(n_1127) );
INVx1_ASAP7_75t_L g1139 ( .A(n_109), .Y(n_1139) );
OAI211xp5_ASAP7_75t_L g1013 ( .A1(n_110), .A2(n_662), .B(n_915), .C(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1024 ( .A(n_110), .Y(n_1024) );
INVx1_ASAP7_75t_L g1418 ( .A(n_111), .Y(n_1418) );
INVx1_ASAP7_75t_L g563 ( .A(n_112), .Y(n_563) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_113), .A2(n_291), .B1(n_363), .B2(n_391), .Y(n_1019) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_113), .A2(n_153), .B1(n_409), .B2(n_419), .Y(n_1025) );
XOR2xp5_ASAP7_75t_L g1360 ( .A(n_114), .B(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g788 ( .A(n_115), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_116), .A2(n_314), .B1(n_1437), .B2(n_1448), .Y(n_1454) );
INVx1_ASAP7_75t_L g384 ( .A(n_117), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_118), .Y(n_1154) );
INVx1_ASAP7_75t_L g542 ( .A(n_120), .Y(n_542) );
INVx1_ASAP7_75t_L g476 ( .A(n_121), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_122), .A2(n_252), .B1(n_927), .B2(n_928), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g979 ( .A1(n_122), .A2(n_252), .B1(n_585), .B2(n_759), .Y(n_979) );
INVx1_ASAP7_75t_L g1275 ( .A(n_123), .Y(n_1275) );
INVx1_ASAP7_75t_L g1250 ( .A(n_124), .Y(n_1250) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_125), .A2(n_216), .B1(n_759), .B2(n_1157), .Y(n_1156) );
OAI22xp33_ASAP7_75t_SL g732 ( .A1(n_126), .A2(n_127), .B1(n_733), .B2(n_734), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_126), .A2(n_131), .B1(n_684), .B2(n_685), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g1686 ( .A1(n_128), .A2(n_260), .B1(n_603), .B2(n_1687), .Y(n_1686) );
AOI221xp5_ASAP7_75t_L g1728 ( .A1(n_128), .A2(n_324), .B1(n_607), .B2(n_1724), .C(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g903 ( .A(n_129), .Y(n_903) );
INVx1_ASAP7_75t_L g1253 ( .A(n_130), .Y(n_1253) );
INVx1_ASAP7_75t_L g730 ( .A(n_131), .Y(n_730) );
INVx1_ASAP7_75t_L g831 ( .A(n_132), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_133), .A2(n_286), .B1(n_955), .B2(n_956), .Y(n_954) );
INVx1_ASAP7_75t_L g1292 ( .A(n_134), .Y(n_1292) );
INVx1_ASAP7_75t_L g1251 ( .A(n_135), .Y(n_1251) );
AOI31xp33_ASAP7_75t_L g1170 ( .A1(n_136), .A2(n_1171), .A3(n_1183), .B(n_1193), .Y(n_1170) );
NAND2xp33_ASAP7_75t_SL g1209 ( .A(n_136), .B(n_1210), .Y(n_1209) );
INVxp67_ASAP7_75t_SL g1222 ( .A(n_136), .Y(n_1222) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_137), .A2(n_183), .B1(n_363), .B2(n_733), .Y(n_1055) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_137), .A2(n_174), .B1(n_409), .B2(n_419), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g1040 ( .A(n_138), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_139), .A2(n_216), .B1(n_777), .B2(n_1166), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_140), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_141), .Y(n_1031) );
OAI211xp5_ASAP7_75t_L g369 ( .A1(n_142), .A2(n_370), .B(n_375), .C(n_380), .Y(n_369) );
INVx1_ASAP7_75t_L g440 ( .A(n_142), .Y(n_440) );
OAI22xp33_ASAP7_75t_L g1277 ( .A1(n_143), .A2(n_156), .B1(n_444), .B2(n_447), .Y(n_1277) );
OAI22xp33_ASAP7_75t_L g1284 ( .A1(n_143), .A2(n_156), .B1(n_363), .B2(n_673), .Y(n_1284) );
INVx1_ASAP7_75t_L g388 ( .A(n_144), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_144), .A2(n_424), .B(n_431), .C(n_435), .Y(n_423) );
INVx1_ASAP7_75t_L g894 ( .A(n_145), .Y(n_894) );
INVx1_ASAP7_75t_L g870 ( .A(n_146), .Y(n_870) );
INVx1_ASAP7_75t_L g471 ( .A(n_148), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_149), .Y(n_631) );
INVx1_ASAP7_75t_L g1129 ( .A(n_150), .Y(n_1129) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_151), .Y(n_800) );
INVx1_ASAP7_75t_L g1349 ( .A(n_152), .Y(n_1349) );
OAI22xp33_ASAP7_75t_L g1018 ( .A1(n_153), .A2(n_268), .B1(n_673), .B2(n_761), .Y(n_1018) );
INVx1_ASAP7_75t_L g1053 ( .A(n_154), .Y(n_1053) );
OAI211xp5_ASAP7_75t_L g1058 ( .A1(n_154), .A2(n_431), .B(n_511), .C(n_1059), .Y(n_1058) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_155), .Y(n_991) );
INVx1_ASAP7_75t_L g1774 ( .A(n_157), .Y(n_1774) );
INVx1_ASAP7_75t_L g1248 ( .A(n_159), .Y(n_1248) );
INVx1_ASAP7_75t_L g756 ( .A(n_160), .Y(n_756) );
OAI211xp5_ASAP7_75t_L g1050 ( .A1(n_161), .A2(n_662), .B(n_915), .C(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1060 ( .A(n_161), .Y(n_1060) );
INVx1_ASAP7_75t_L g1291 ( .A(n_162), .Y(n_1291) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_164), .Y(n_637) );
INVx1_ASAP7_75t_L g1563 ( .A(n_165), .Y(n_1563) );
AOI22xp5_ASAP7_75t_SL g1465 ( .A1(n_166), .A2(n_177), .B1(n_1440), .B2(n_1448), .Y(n_1465) );
INVx1_ASAP7_75t_L g501 ( .A(n_168), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_169), .A2(n_251), .B1(n_759), .B2(n_760), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_169), .A2(n_251), .B1(n_765), .B2(n_766), .Y(n_764) );
OAI22xp33_ASAP7_75t_L g1054 ( .A1(n_171), .A2(n_174), .B1(n_673), .B2(n_761), .Y(n_1054) );
OAI22xp33_ASAP7_75t_L g1057 ( .A1(n_171), .A2(n_183), .B1(n_446), .B2(n_690), .Y(n_1057) );
INVx1_ASAP7_75t_L g871 ( .A(n_172), .Y(n_871) );
OAI211xp5_ASAP7_75t_L g877 ( .A1(n_172), .A2(n_370), .B(n_375), .C(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g797 ( .A(n_173), .Y(n_797) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_175), .A2(n_286), .B1(n_965), .B2(n_969), .Y(n_964) );
OAI22xp33_ASAP7_75t_SL g675 ( .A1(n_176), .A2(n_296), .B1(n_363), .B2(n_391), .Y(n_675) );
INVx1_ASAP7_75t_L g1244 ( .A(n_179), .Y(n_1244) );
INVx2_ASAP7_75t_L g1435 ( .A(n_180), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_180), .B(n_1436), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_180), .B(n_293), .Y(n_1443) );
AOI22xp5_ASAP7_75t_SL g1485 ( .A1(n_184), .A2(n_259), .B1(n_1437), .B2(n_1442), .Y(n_1485) );
CKINVDCx5p33_ASAP7_75t_R g1036 ( .A(n_185), .Y(n_1036) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_186), .Y(n_708) );
INVx1_ASAP7_75t_L g792 ( .A(n_187), .Y(n_792) );
INVx1_ASAP7_75t_L g891 ( .A(n_188), .Y(n_891) );
INVx1_ASAP7_75t_L g825 ( .A(n_189), .Y(n_825) );
OAI21xp33_ASAP7_75t_L g1667 ( .A1(n_191), .A2(n_1668), .B(n_1674), .Y(n_1667) );
OAI221xp5_ASAP7_75t_L g1738 ( .A1(n_191), .A2(n_282), .B1(n_522), .B2(n_1147), .C(n_1739), .Y(n_1738) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_192), .A2(n_276), .B1(n_726), .B2(n_733), .Y(n_1199) );
AOI22xp5_ASAP7_75t_L g1439 ( .A1(n_193), .A2(n_309), .B1(n_1440), .B2(n_1442), .Y(n_1439) );
INVx1_ASAP7_75t_L g1155 ( .A(n_194), .Y(n_1155) );
OAI211xp5_ASAP7_75t_L g1161 ( .A1(n_194), .A2(n_431), .B(n_1162), .C(n_1163), .Y(n_1161) );
INVx1_ASAP7_75t_L g1380 ( .A(n_195), .Y(n_1380) );
AOI22xp5_ASAP7_75t_L g1446 ( .A1(n_196), .A2(n_261), .B1(n_1432), .B2(n_1437), .Y(n_1446) );
INVx1_ASAP7_75t_L g1106 ( .A(n_197), .Y(n_1106) );
OAI22xp33_ASAP7_75t_L g1116 ( .A1(n_197), .A2(n_228), .B1(n_363), .B2(n_673), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_198), .A2(n_321), .B1(n_936), .B2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_198), .A2(n_245), .B1(n_965), .B2(n_969), .Y(n_971) );
INVx1_ASAP7_75t_L g1768 ( .A(n_199), .Y(n_1768) );
INVx1_ASAP7_75t_L g1231 ( .A(n_200), .Y(n_1231) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_202), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g1455 ( .A1(n_204), .A2(n_278), .B1(n_1432), .B2(n_1440), .Y(n_1455) );
INVx1_ASAP7_75t_L g822 ( .A(n_205), .Y(n_822) );
OAI211xp5_ASAP7_75t_L g1363 ( .A1(n_206), .A2(n_856), .B(n_1364), .C(n_1372), .Y(n_1363) );
INVx1_ASAP7_75t_L g1399 ( .A(n_206), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g1270 ( .A1(n_208), .A2(n_232), .B1(n_408), .B2(n_1166), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g1283 ( .A1(n_208), .A2(n_232), .B1(n_759), .B2(n_1112), .Y(n_1283) );
AOI22xp33_ASAP7_75t_SL g1685 ( .A1(n_209), .A2(n_313), .B1(n_967), .B2(n_1321), .Y(n_1685) );
AOI221xp5_ASAP7_75t_L g1725 ( .A1(n_209), .A2(n_231), .B1(n_607), .B2(n_1726), .C(n_1727), .Y(n_1725) );
INVx1_ASAP7_75t_L g1771 ( .A(n_210), .Y(n_1771) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_211), .A2(n_287), .B1(n_354), .B2(n_363), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g443 ( .A1(n_211), .A2(n_287), .B1(n_444), .B2(n_447), .Y(n_443) );
INVx2_ASAP7_75t_L g456 ( .A(n_212), .Y(n_456) );
INVx1_ASAP7_75t_L g530 ( .A(n_212), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g1737 ( .A(n_212), .B(n_412), .Y(n_1737) );
CKINVDCx5p33_ASAP7_75t_R g992 ( .A(n_213), .Y(n_992) );
XOR2xp5_ASAP7_75t_L g816 ( .A(n_214), .B(n_817), .Y(n_816) );
OAI22xp33_ASAP7_75t_L g1227 ( .A1(n_215), .A2(n_275), .B1(n_726), .B2(n_733), .Y(n_1227) );
OAI22xp5_ASAP7_75t_SL g1234 ( .A1(n_215), .A2(n_244), .B1(n_409), .B2(n_446), .Y(n_1234) );
INVx1_ASAP7_75t_L g1081 ( .A(n_217), .Y(n_1081) );
XOR2xp5_ASAP7_75t_L g919 ( .A(n_219), .B(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g1371 ( .A(n_220), .Y(n_1371) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_220), .A2(n_249), .B1(n_409), .B2(n_419), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1704 ( .A1(n_221), .A2(n_323), .B1(n_603), .B2(n_1705), .Y(n_1704) );
AOI22xp33_ASAP7_75t_L g1723 ( .A1(n_221), .A2(n_260), .B1(n_1339), .B2(n_1724), .Y(n_1723) );
INVx1_ASAP7_75t_L g1365 ( .A(n_222), .Y(n_1365) );
INVx1_ASAP7_75t_L g1099 ( .A(n_223), .Y(n_1099) );
OA211x2_ASAP7_75t_L g1113 ( .A1(n_223), .A2(n_483), .B(n_753), .C(n_1114), .Y(n_1113) );
BUFx3_ASAP7_75t_L g414 ( .A(n_224), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_225), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g1043 ( .A(n_226), .Y(n_1043) );
OAI22xp5_ASAP7_75t_SL g1065 ( .A1(n_227), .A2(n_1066), .B1(n_1109), .B2(n_1118), .Y(n_1065) );
NAND4xp25_ASAP7_75t_L g1066 ( .A(n_227), .B(n_1067), .C(n_1083), .D(n_1093), .Y(n_1066) );
INVx1_ASAP7_75t_L g1103 ( .A(n_228), .Y(n_1103) );
INVx1_ASAP7_75t_L g1675 ( .A(n_229), .Y(n_1675) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_230), .A2(n_245), .B1(n_936), .B2(n_942), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_230), .A2(n_321), .B1(n_961), .B2(n_962), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1707 ( .A1(n_231), .A2(n_324), .B1(n_965), .B2(n_969), .Y(n_1707) );
OA22x2_ASAP7_75t_L g1267 ( .A1(n_233), .A2(n_1268), .B1(n_1310), .B2(n_1311), .Y(n_1267) );
INVxp67_ASAP7_75t_L g1311 ( .A(n_233), .Y(n_1311) );
AOI22xp5_ASAP7_75t_L g1431 ( .A1(n_233), .A2(n_270), .B1(n_1432), .B2(n_1437), .Y(n_1431) );
INVx1_ASAP7_75t_L g552 ( .A(n_234), .Y(n_552) );
INVx1_ASAP7_75t_L g1348 ( .A(n_235), .Y(n_1348) );
INVx1_ASAP7_75t_L g1376 ( .A(n_236), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1404 ( .A(n_236), .B(n_1405), .Y(n_1404) );
CKINVDCx5p33_ASAP7_75t_R g1035 ( .A(n_237), .Y(n_1035) );
INVx1_ASAP7_75t_L g1073 ( .A(n_238), .Y(n_1073) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_239), .Y(n_994) );
INVx1_ASAP7_75t_L g829 ( .A(n_240), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_241), .A2(n_307), .B1(n_354), .B2(n_363), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g774 ( .A1(n_241), .A2(n_307), .B1(n_775), .B2(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g482 ( .A(n_242), .Y(n_482) );
INVx1_ASAP7_75t_L g1230 ( .A(n_243), .Y(n_1230) );
OAI22xp33_ASAP7_75t_L g1232 ( .A1(n_244), .A2(n_281), .B1(n_673), .B2(n_734), .Y(n_1232) );
INVx1_ASAP7_75t_L g560 ( .A(n_246), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_246), .A2(n_294), .B1(n_594), .B2(n_596), .Y(n_593) );
XOR2xp5_ASAP7_75t_L g693 ( .A(n_247), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g789 ( .A(n_248), .Y(n_789) );
INVx1_ASAP7_75t_L g1373 ( .A(n_249), .Y(n_1373) );
BUFx3_ASAP7_75t_L g362 ( .A(n_250), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_250), .Y(n_366) );
XOR2x2_ASAP7_75t_L g864 ( .A(n_253), .B(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g1098 ( .A(n_255), .Y(n_1098) );
INVx1_ASAP7_75t_L g1767 ( .A(n_256), .Y(n_1767) );
INVx1_ASAP7_75t_L g1082 ( .A(n_257), .Y(n_1082) );
AOI22xp5_ASAP7_75t_L g1172 ( .A1(n_258), .A2(n_283), .B1(n_1101), .B2(n_1173), .Y(n_1172) );
INVxp67_ASAP7_75t_SL g1657 ( .A(n_261), .Y(n_1657) );
AOI22xp33_ASAP7_75t_L g1754 ( .A1(n_261), .A2(n_1755), .B1(n_1760), .B2(n_1802), .Y(n_1754) );
INVx1_ASAP7_75t_L g924 ( .A(n_262), .Y(n_924) );
INVx1_ASAP7_75t_L g821 ( .A(n_263), .Y(n_821) );
OAI211xp5_ASAP7_75t_L g1228 ( .A1(n_264), .A2(n_483), .B(n_662), .C(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1239 ( .A(n_264), .Y(n_1239) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_265), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_266), .B(n_409), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_267), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g1021 ( .A1(n_268), .A2(n_291), .B1(n_446), .B2(n_690), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_269), .Y(n_638) );
INVx1_ASAP7_75t_L g1077 ( .A(n_271), .Y(n_1077) );
XOR2x2_ASAP7_75t_L g350 ( .A(n_272), .B(n_351), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_273), .Y(n_1033) );
XOR2x2_ASAP7_75t_L g1313 ( .A(n_274), .B(n_1314), .Y(n_1313) );
OAI22xp33_ASAP7_75t_L g1240 ( .A1(n_275), .A2(n_281), .B1(n_419), .B2(n_690), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1191 ( .A1(n_276), .A2(n_310), .B1(n_419), .B2(n_690), .Y(n_1191) );
INVx1_ASAP7_75t_L g1346 ( .A(n_277), .Y(n_1346) );
INVx1_ASAP7_75t_L g416 ( .A(n_279), .Y(n_416) );
INVx1_ASAP7_75t_L g422 ( .A(n_279), .Y(n_422) );
INVx1_ASAP7_75t_L g1702 ( .A(n_280), .Y(n_1702) );
INVxp67_ASAP7_75t_SL g1749 ( .A(n_282), .Y(n_1749) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_283), .A2(n_312), .B1(n_1214), .B2(n_1216), .Y(n_1217) );
INVx1_ASAP7_75t_L g1074 ( .A(n_284), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g846 ( .A1(n_285), .A2(n_688), .B(n_847), .C(n_849), .Y(n_846) );
INVx1_ASAP7_75t_L g859 ( .A(n_285), .Y(n_859) );
INVx1_ASAP7_75t_L g555 ( .A(n_288), .Y(n_555) );
INVx1_ASAP7_75t_L g667 ( .A(n_289), .Y(n_667) );
OAI211xp5_ASAP7_75t_SL g679 ( .A1(n_289), .A2(n_609), .B(n_680), .C(n_688), .Y(n_679) );
INVx1_ASAP7_75t_L g895 ( .A(n_290), .Y(n_895) );
INVx1_ASAP7_75t_L g1770 ( .A(n_292), .Y(n_1770) );
INVx1_ASAP7_75t_L g1436 ( .A(n_293), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_293), .B(n_1435), .Y(n_1441) );
INVx1_ASAP7_75t_L g538 ( .A(n_294), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g995 ( .A(n_295), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_296), .A2(n_331), .B1(n_409), .B2(n_419), .Y(n_678) );
INVx1_ASAP7_75t_L g923 ( .A(n_297), .Y(n_923) );
INVx1_ASAP7_75t_L g566 ( .A(n_298), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_299), .Y(n_1052) );
INVx1_ASAP7_75t_L g1565 ( .A(n_300), .Y(n_1565) );
CKINVDCx5p33_ASAP7_75t_R g1382 ( .A(n_301), .Y(n_1382) );
OAI211xp5_ASAP7_75t_SL g727 ( .A1(n_303), .A2(n_661), .B(n_662), .C(n_728), .Y(n_727) );
OAI211xp5_ASAP7_75t_SL g738 ( .A1(n_303), .A2(n_688), .B(n_739), .C(n_740), .Y(n_738) );
INVx1_ASAP7_75t_L g1245 ( .A(n_304), .Y(n_1245) );
INVx1_ASAP7_75t_L g1790 ( .A(n_305), .Y(n_1790) );
XOR2x2_ASAP7_75t_L g1224 ( .A(n_306), .B(n_1225), .Y(n_1224) );
OAI211xp5_ASAP7_75t_L g1152 ( .A1(n_308), .A2(n_722), .B(n_753), .C(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1164 ( .A(n_308), .Y(n_1164) );
INVxp67_ASAP7_75t_SL g1197 ( .A(n_310), .Y(n_1197) );
AOI22xp33_ASAP7_75t_SL g1332 ( .A1(n_311), .A2(n_341), .B1(n_1333), .B2(n_1336), .Y(n_1332) );
INVx1_ASAP7_75t_L g1180 ( .A(n_312), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1731 ( .A1(n_313), .A2(n_323), .B1(n_1339), .B2(n_1732), .Y(n_1731) );
OAI211xp5_ASAP7_75t_SL g749 ( .A1(n_315), .A2(n_750), .B(n_753), .C(n_754), .Y(n_749) );
INVx1_ASAP7_75t_L g772 ( .A(n_315), .Y(n_772) );
INVx1_ASAP7_75t_L g785 ( .A(n_316), .Y(n_785) );
INVx1_ASAP7_75t_L g1288 ( .A(n_317), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_318), .Y(n_641) );
INVx1_ASAP7_75t_L g1070 ( .A(n_319), .Y(n_1070) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_320), .Y(n_358) );
INVx1_ASAP7_75t_L g488 ( .A(n_322), .Y(n_488) );
INVx1_ASAP7_75t_L g827 ( .A(n_326), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_327), .Y(n_1016) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_328), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_329), .Y(n_703) );
INVx1_ASAP7_75t_L g405 ( .A(n_332), .Y(n_405) );
INVx2_ASAP7_75t_L g466 ( .A(n_332), .Y(n_466) );
INVx1_ASAP7_75t_L g529 ( .A(n_332), .Y(n_529) );
INVx1_ASAP7_75t_L g851 ( .A(n_333), .Y(n_851) );
INVx1_ASAP7_75t_L g1125 ( .A(n_334), .Y(n_1125) );
INVx1_ASAP7_75t_L g1108 ( .A(n_336), .Y(n_1108) );
INVx1_ASAP7_75t_L g491 ( .A(n_337), .Y(n_491) );
AOI21xp33_ASAP7_75t_L g1383 ( .A1(n_338), .A2(n_1214), .B(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1402 ( .A(n_338), .Y(n_1402) );
INVx1_ASAP7_75t_L g902 ( .A(n_339), .Y(n_902) );
INVx1_ASAP7_75t_L g1100 ( .A(n_340), .Y(n_1100) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_342), .Y(n_1003) );
CKINVDCx5p33_ASAP7_75t_R g1369 ( .A(n_343), .Y(n_1369) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_1411), .B(n_1424), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_1263), .B1(n_1264), .B2(n_1410), .Y(n_345) );
INVx1_ASAP7_75t_L g1410 ( .A(n_346), .Y(n_1410) );
AO22x1_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_861), .B1(n_1261), .B2(n_1262), .Y(n_346) );
INVx1_ASAP7_75t_L g1262 ( .A(n_347), .Y(n_1262) );
XNOR2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_743), .Y(n_347) );
XOR2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_620), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_532), .B1(n_618), .B2(n_619), .Y(n_349) );
INVx2_ASAP7_75t_L g618 ( .A(n_350), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_406), .C(n_460), .Y(n_351) );
OAI31xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_369), .A3(n_389), .B(n_398), .Y(n_352) );
INVx3_ASAP7_75t_L g567 ( .A(n_354), .Y(n_567) );
OR2x6_ASAP7_75t_L g354 ( .A(n_355), .B(n_360), .Y(n_354) );
OR2x6_ASAP7_75t_L g391 ( .A(n_355), .B(n_365), .Y(n_391) );
BUFx4f_ASAP7_75t_L g470 ( .A(n_355), .Y(n_470) );
INVx1_ASAP7_75t_L g656 ( .A(n_355), .Y(n_656) );
OR2x2_ASAP7_75t_L g733 ( .A(n_355), .B(n_365), .Y(n_733) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx4f_ASAP7_75t_L g500 ( .A(n_356), .Y(n_500) );
INVx3_ASAP7_75t_L g674 ( .A(n_356), .Y(n_674) );
INVx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AND2x2_ASAP7_75t_L g367 ( .A(n_358), .B(n_368), .Y(n_367) );
NAND2x1_ASAP7_75t_L g374 ( .A(n_358), .B(n_359), .Y(n_374) );
AND2x2_ASAP7_75t_L g379 ( .A(n_358), .B(n_359), .Y(n_379) );
INVx1_ASAP7_75t_L g387 ( .A(n_358), .Y(n_387) );
INVx2_ASAP7_75t_L g397 ( .A(n_358), .Y(n_397) );
INVx2_ASAP7_75t_L g481 ( .A(n_358), .Y(n_481) );
INVx2_ASAP7_75t_L g368 ( .A(n_359), .Y(n_368) );
BUFx2_ASAP7_75t_L g383 ( .A(n_359), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_359), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g480 ( .A(n_359), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g582 ( .A(n_359), .Y(n_582) );
AND2x2_ASAP7_75t_L g598 ( .A(n_359), .B(n_397), .Y(n_598) );
OR2x6_ASAP7_75t_L g673 ( .A(n_360), .B(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g1368 ( .A1(n_360), .A2(n_1369), .B1(n_1370), .B2(n_1371), .Y(n_1368) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g377 ( .A(n_361), .Y(n_377) );
AND2x4_ASAP7_75t_L g1385 ( .A(n_361), .B(n_401), .Y(n_1385) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g382 ( .A(n_362), .Y(n_382) );
AND2x4_ASAP7_75t_L g385 ( .A(n_362), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g494 ( .A(n_362), .B(n_401), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g363 ( .A(n_364), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_364), .A2(n_566), .B1(n_567), .B2(n_568), .Y(n_565) );
INVx4_ASAP7_75t_L g734 ( .A(n_364), .Y(n_734) );
INVx3_ASAP7_75t_SL g856 ( .A(n_364), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_364), .A2(n_567), .B1(n_923), .B2(n_924), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_364), .A2(n_1195), .B1(n_1196), .B2(n_1197), .Y(n_1194) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g968 ( .A(n_367), .Y(n_968) );
BUFx6f_ASAP7_75t_L g1215 ( .A(n_367), .Y(n_1215) );
BUFx3_ASAP7_75t_L g1320 ( .A(n_367), .Y(n_1320) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g590 ( .A1(n_372), .A2(n_545), .B1(n_552), .B2(n_591), .C(n_593), .Y(n_590) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_372), .A2(n_542), .B1(n_563), .B2(n_600), .C(n_602), .Y(n_599) );
BUFx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_SL g484 ( .A(n_373), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g790 ( .A1(n_373), .A2(n_791), .B1(n_792), .B2(n_793), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_373), .A2(n_791), .B1(n_822), .B2(n_835), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g1008 ( .A1(n_373), .A2(n_992), .B1(n_1003), .B2(n_1009), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_373), .A2(n_1007), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
OR2x2_ASAP7_75t_L g1682 ( .A(n_373), .B(n_1678), .Y(n_1682) );
BUFx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_374), .Y(n_490) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI211xp5_ASAP7_75t_L g569 ( .A1(n_376), .A2(n_570), .B(n_573), .C(n_574), .Y(n_569) );
INVx3_ASAP7_75t_L g753 ( .A(n_376), .Y(n_753) );
NOR3xp33_ASAP7_75t_L g978 ( .A(n_376), .B(n_979), .C(n_980), .Y(n_978) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x2_ASAP7_75t_L g663 ( .A(n_377), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g726 ( .A(n_377), .B(n_395), .Y(n_726) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_377), .B(n_383), .Y(n_1015) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_378), .Y(n_572) );
BUFx3_ASAP7_75t_L g1216 ( .A(n_378), .Y(n_1216) );
BUFx3_ASAP7_75t_L g1321 ( .A(n_378), .Y(n_1321) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g665 ( .A(n_379), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B1(n_385), .B2(n_388), .Y(n_380) );
INVx1_ASAP7_75t_L g575 ( .A(n_381), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_381), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_728) );
BUFx3_ASAP7_75t_L g755 ( .A(n_381), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_381), .A2(n_385), .B1(n_851), .B2(n_859), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_381), .A2(n_879), .B1(n_1098), .B2(n_1100), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_381), .A2(n_670), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_381), .A2(n_731), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
AOI222xp33_ASAP7_75t_L g1347 ( .A1(n_381), .A2(n_731), .B1(n_1321), .B2(n_1348), .C1(n_1349), .C2(n_1350), .Y(n_1347) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OR2x2_ASAP7_75t_L g394 ( .A(n_382), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g579 ( .A(n_382), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g668 ( .A(n_382), .B(n_383), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g1364 ( .A1(n_382), .A2(n_1321), .B(n_1365), .C(n_1366), .Y(n_1364) );
INVx1_ASAP7_75t_L g1370 ( .A(n_382), .Y(n_1370) );
INVx1_ASAP7_75t_L g1697 ( .A(n_383), .Y(n_1697) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_384), .A2(n_436), .B1(n_440), .B2(n_441), .Y(n_435) );
INVx2_ASAP7_75t_L g576 ( .A(n_385), .Y(n_576) );
INVx2_ASAP7_75t_L g671 ( .A(n_385), .Y(n_671) );
BUFx3_ASAP7_75t_L g731 ( .A(n_385), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_385), .A2(n_1015), .B1(n_1187), .B2(n_1189), .Y(n_1201) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_386), .B(n_1673), .Y(n_1701) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_391), .Y(n_759) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g1112 ( .A(n_393), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g1157 ( .A(n_393), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1344 ( .A1(n_393), .A2(n_579), .B1(n_1345), .B2(n_1346), .Y(n_1344) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g586 ( .A(n_394), .Y(n_586) );
BUFx2_ASAP7_75t_L g761 ( .A(n_394), .Y(n_761) );
INVx8_ASAP7_75t_L g474 ( .A(n_395), .Y(n_474) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_395), .Y(n_1088) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI31xp33_ASAP7_75t_L g854 ( .A1(n_398), .A2(n_855), .A3(n_857), .B(n_860), .Y(n_854) );
OAI31xp33_ASAP7_75t_L g1278 ( .A1(n_398), .A2(n_1279), .A3(n_1283), .B(n_1284), .Y(n_1278) );
OAI21xp5_ASAP7_75t_L g1342 ( .A1(n_398), .A2(n_1343), .B(n_1351), .Y(n_1342) );
BUFx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g587 ( .A(n_399), .Y(n_587) );
BUFx2_ASAP7_75t_L g676 ( .A(n_399), .Y(n_676) );
OAI31xp33_ASAP7_75t_L g724 ( .A1(n_399), .A2(n_725), .A3(n_727), .B(n_732), .Y(n_724) );
BUFx3_ASAP7_75t_L g885 ( .A(n_399), .Y(n_885) );
OAI31xp33_ASAP7_75t_L g1226 ( .A1(n_399), .A2(n_1227), .A3(n_1228), .B(n_1232), .Y(n_1226) );
OAI21xp5_ASAP7_75t_L g1793 ( .A1(n_399), .A2(n_1794), .B(n_1801), .Y(n_1793) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_402), .Y(n_399) );
AOI21xp5_ASAP7_75t_SL g1362 ( .A1(n_400), .A2(n_1363), .B(n_1374), .Y(n_1362) );
INVx1_ASAP7_75t_L g1423 ( .A(n_400), .Y(n_1423) );
NOR2xp33_ASAP7_75t_L g1753 ( .A(n_400), .B(n_1415), .Y(n_1753) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g1663 ( .A(n_403), .Y(n_1663) );
OR2x2_ASAP7_75t_L g1700 ( .A(n_403), .B(n_1701), .Y(n_1700) );
BUFx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g459 ( .A(n_404), .Y(n_459) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI31xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_423), .A3(n_443), .B(n_453), .Y(n_406) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g614 ( .A(n_409), .Y(n_614) );
BUFx2_ASAP7_75t_L g765 ( .A(n_409), .Y(n_765) );
BUFx2_ASAP7_75t_L g927 ( .A(n_409), .Y(n_927) );
OR2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
AND2x4_ASAP7_75t_L g448 ( .A(n_410), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g691 ( .A(n_410), .B(n_449), .Y(n_691) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x6_ASAP7_75t_L g419 ( .A(n_411), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g432 ( .A(n_411), .B(n_433), .Y(n_432) );
OR2x4_ASAP7_75t_L g446 ( .A(n_411), .B(n_413), .Y(n_446) );
NAND3x1_ASAP7_75t_L g527 ( .A(n_411), .B(n_528), .C(n_530), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g643 ( .A(n_411), .B(n_530), .Y(n_643) );
AND2x4_ASAP7_75t_L g1715 ( .A(n_411), .B(n_1716), .Y(n_1715) );
INVx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g438 ( .A(n_412), .Y(n_438) );
NAND2xp33_ASAP7_75t_SL g506 ( .A(n_412), .B(n_456), .Y(n_506) );
INVx2_ASAP7_75t_L g510 ( .A(n_413), .Y(n_510) );
BUFx4f_ASAP7_75t_L g628 ( .A(n_413), .Y(n_628) );
BUFx3_ASAP7_75t_L g804 ( .A(n_413), .Y(n_804) );
BUFx3_ASAP7_75t_L g814 ( .A(n_413), .Y(n_814) );
OR2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_414), .B(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_414), .Y(n_430) );
AND2x4_ASAP7_75t_L g433 ( .A(n_414), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
INVx1_ASAP7_75t_L g941 ( .A(n_415), .Y(n_941) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_L g451 ( .A(n_416), .Y(n_451) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g615 ( .A(n_419), .Y(n_615) );
INVx1_ASAP7_75t_L g874 ( .A(n_419), .Y(n_874) );
BUFx3_ASAP7_75t_L g1166 ( .A(n_419), .Y(n_1166) );
INVx1_ASAP7_75t_L g519 ( .A(n_420), .Y(n_519) );
BUFx3_ASAP7_75t_L g809 ( .A(n_420), .Y(n_809) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g524 ( .A(n_421), .Y(n_524) );
INVx1_ASAP7_75t_L g429 ( .A(n_422), .Y(n_429) );
INVx2_ASAP7_75t_L g434 ( .A(n_422), .Y(n_434) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_425), .A2(n_471), .B1(n_491), .B2(n_508), .Y(n_531) );
OAI22xp33_ASAP7_75t_L g1141 ( .A1(n_425), .A2(n_1125), .B1(n_1134), .B2(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g768 ( .A(n_426), .Y(n_768) );
INVx1_ASAP7_75t_L g834 ( .A(n_426), .Y(n_834) );
INVx1_ASAP7_75t_L g930 ( .A(n_426), .Y(n_930) );
INVx1_ASAP7_75t_L g1162 ( .A(n_426), .Y(n_1162) );
INVx2_ASAP7_75t_L g1394 ( .A(n_426), .Y(n_1394) );
INVx4_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_427), .Y(n_543) );
INVx3_ASAP7_75t_L g700 ( .A(n_427), .Y(n_700) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g513 ( .A(n_428), .Y(n_513) );
BUFx3_ASAP7_75t_L g562 ( .A(n_428), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
BUFx2_ASAP7_75t_L g442 ( .A(n_429), .Y(n_442) );
BUFx2_ASAP7_75t_L g439 ( .A(n_430), .Y(n_439) );
INVx2_ASAP7_75t_L g685 ( .A(n_430), .Y(n_685) );
AND2x4_ASAP7_75t_L g950 ( .A(n_430), .B(n_683), .Y(n_950) );
NAND3xp33_ASAP7_75t_SL g1185 ( .A(n_431), .B(n_1186), .C(n_1188), .Y(n_1185) );
NAND3xp33_ASAP7_75t_SL g1235 ( .A(n_431), .B(n_1236), .C(n_1238), .Y(n_1235) );
CKINVDCx8_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_432), .A2(n_606), .B(n_607), .C(n_608), .Y(n_605) );
CKINVDCx8_ASAP7_75t_R g688 ( .A(n_432), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g925 ( .A(n_432), .B(n_926), .C(n_929), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g1095 ( .A(n_432), .B(n_1096), .Y(n_1095) );
NOR3xp33_ASAP7_75t_L g1392 ( .A(n_432), .B(n_1393), .C(n_1397), .Y(n_1392) );
BUFx3_ASAP7_75t_L g607 ( .A(n_433), .Y(n_607) );
INVx2_ASAP7_75t_L g943 ( .A(n_433), .Y(n_943) );
BUFx2_ASAP7_75t_L g953 ( .A(n_433), .Y(n_953) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_433), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1237 ( .A(n_433), .Y(n_1237) );
BUFx2_ASAP7_75t_L g1788 ( .A(n_433), .Y(n_1788) );
INVx1_ASAP7_75t_L g683 ( .A(n_434), .Y(n_683) );
INVx1_ASAP7_75t_L g609 ( .A(n_436), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_436), .A2(n_441), .B1(n_1154), .B2(n_1164), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_436), .A2(n_441), .B1(n_1275), .B2(n_1276), .Y(n_1274) );
AND2x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
AND2x4_ASAP7_75t_L g441 ( .A(n_437), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g686 ( .A(n_437), .B(n_442), .Y(n_686) );
AND2x4_ASAP7_75t_L g742 ( .A(n_437), .B(n_439), .Y(n_742) );
AND2x2_ASAP7_75t_L g771 ( .A(n_437), .B(n_439), .Y(n_771) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g681 ( .A(n_438), .B(n_682), .Y(n_681) );
AND3x4_ASAP7_75t_L g933 ( .A(n_438), .B(n_456), .C(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g610 ( .A(n_441), .Y(n_610) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_441), .Y(n_773) );
AOI222xp33_ASAP7_75t_L g1097 ( .A1(n_441), .A2(n_742), .B1(n_1098), .B2(n_1099), .C1(n_1100), .C2(n_1101), .Y(n_1097) );
AOI222xp33_ASAP7_75t_L g1356 ( .A1(n_441), .A2(n_770), .B1(n_1101), .B2(n_1348), .C1(n_1349), .C2(n_1350), .Y(n_1356) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g1398 ( .A1(n_445), .A2(n_691), .B1(n_1369), .B2(n_1399), .Y(n_1398) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_SL g612 ( .A(n_446), .Y(n_612) );
INVx2_ASAP7_75t_SL g776 ( .A(n_446), .Y(n_776) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_446), .Y(n_844) );
INVx1_ASAP7_75t_L g1107 ( .A(n_446), .Y(n_1107) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_448), .A2(n_566), .B1(n_568), .B2(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g777 ( .A(n_448), .Y(n_777) );
INVx1_ASAP7_75t_L g845 ( .A(n_448), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_448), .A2(n_612), .B1(n_923), .B2(n_924), .Y(n_922) );
INVx2_ASAP7_75t_L g704 ( .A(n_449), .Y(n_704) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_449), .Y(n_808) );
INVx1_ASAP7_75t_L g830 ( .A(n_449), .Y(n_830) );
INVx2_ASAP7_75t_L g1147 ( .A(n_449), .Y(n_1147) );
BUFx6f_ASAP7_75t_L g1307 ( .A(n_449), .Y(n_1307) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_450), .Y(n_516) );
BUFx8_ASAP7_75t_L g551 ( .A(n_450), .Y(n_551) );
INVx2_ASAP7_75t_L g947 ( .A(n_450), .Y(n_947) );
AND2x4_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
AND2x4_ASAP7_75t_L g940 ( .A(n_452), .B(n_941), .Y(n_940) );
OAI31xp33_ASAP7_75t_L g842 ( .A1(n_453), .A2(n_843), .A3(n_846), .B(n_853), .Y(n_842) );
OAI31xp33_ASAP7_75t_L g1159 ( .A1(n_453), .A2(n_1160), .A3(n_1161), .B(n_1165), .Y(n_1159) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_457), .Y(n_453) );
AND2x4_ASAP7_75t_L g617 ( .A(n_454), .B(n_457), .Y(n_617) );
AND2x2_ASAP7_75t_L g692 ( .A(n_454), .B(n_457), .Y(n_692) );
AND2x2_ASAP7_75t_SL g778 ( .A(n_454), .B(n_457), .Y(n_778) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_454), .B(n_457), .Y(n_1192) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g1716 ( .A(n_456), .Y(n_1716) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g496 ( .A(n_459), .Y(n_496) );
OR2x2_ASAP7_75t_L g505 ( .A(n_459), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_SL g658 ( .A(n_459), .B(n_494), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_503), .Y(n_460) );
OAI33xp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_468), .A3(n_475), .B1(n_485), .B2(n_492), .B3(n_497), .Y(n_461) );
OAI33xp33_ASAP7_75t_L g836 ( .A1(n_462), .A2(n_794), .A3(n_837), .B1(n_839), .B2(n_840), .B3(n_841), .Y(n_836) );
INVx1_ASAP7_75t_L g959 ( .A(n_462), .Y(n_959) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI33xp33_ASAP7_75t_L g714 ( .A1(n_463), .A2(n_657), .A3(n_715), .B1(n_719), .B2(n_721), .B3(n_723), .Y(n_714) );
OAI33xp33_ASAP7_75t_L g1029 ( .A1(n_463), .A2(n_1011), .A3(n_1030), .B1(n_1034), .B2(n_1037), .B3(n_1041), .Y(n_1029) );
OAI33xp33_ASAP7_75t_L g1242 ( .A1(n_463), .A2(n_1011), .A3(n_1243), .B1(n_1246), .B2(n_1249), .B3(n_1252), .Y(n_1242) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g589 ( .A(n_464), .Y(n_589) );
INVx4_ASAP7_75t_L g781 ( .A(n_464), .Y(n_781) );
INVx2_ASAP7_75t_L g905 ( .A(n_464), .Y(n_905) );
AOI31xp33_ASAP7_75t_L g1684 ( .A1(n_464), .A2(n_1685), .A3(n_1686), .B(n_1688), .Y(n_1684) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
OR2x2_ASAP7_75t_L g642 ( .A(n_465), .B(n_643), .Y(n_642) );
OR2x6_ASAP7_75t_L g1079 ( .A(n_465), .B(n_643), .Y(n_1079) );
INVx1_ASAP7_75t_L g1389 ( .A(n_465), .Y(n_1389) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g934 ( .A(n_466), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g1692 ( .A(n_466), .B(n_1673), .Y(n_1692) );
OAI22xp33_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B1(n_471), .B2(n_472), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_469), .A2(n_488), .B1(n_508), .B2(n_511), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g1087 ( .A1(n_470), .A2(n_1070), .B1(n_1081), .B2(n_1088), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_470), .A2(n_1032), .B1(n_1074), .B2(n_1078), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1375 ( .A1(n_470), .A2(n_472), .B1(n_1376), .B2(n_1377), .Y(n_1375) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_472), .A2(n_498), .B1(n_501), .B2(n_502), .Y(n_497) );
OAI22xp33_ASAP7_75t_L g1287 ( .A1(n_472), .A2(n_1126), .B1(n_1288), .B2(n_1289), .Y(n_1287) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_472), .A2(n_1297), .B1(n_1299), .B2(n_1300), .Y(n_1296) );
INVx5_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx6_ASAP7_75t_L g786 ( .A(n_473), .Y(n_786) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g647 ( .A(n_474), .Y(n_647) );
INVx2_ASAP7_75t_L g718 ( .A(n_474), .Y(n_718) );
INVx1_ASAP7_75t_L g799 ( .A(n_474), .Y(n_799) );
INVx1_ASAP7_75t_L g838 ( .A(n_474), .Y(n_838) );
INVx2_ASAP7_75t_SL g1032 ( .A(n_474), .Y(n_1032) );
INVx2_ASAP7_75t_L g1138 ( .A(n_474), .Y(n_1138) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_482), .B2(n_483), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_476), .A2(n_501), .B1(n_515), .B2(n_517), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_477), .A2(n_720), .B1(n_825), .B2(n_829), .Y(n_839) );
INVx4_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g791 ( .A(n_478), .Y(n_791) );
INVx2_ASAP7_75t_L g1130 ( .A(n_478), .Y(n_1130) );
INVx4_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g487 ( .A(n_480), .Y(n_487) );
INVx2_ASAP7_75t_L g592 ( .A(n_480), .Y(n_592) );
INVx1_ASAP7_75t_L g650 ( .A(n_480), .Y(n_650) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_480), .Y(n_1009) );
AND2x2_ASAP7_75t_L g581 ( .A(n_481), .B(n_582), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_482), .A2(n_502), .B1(n_521), .B2(n_522), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_483), .A2(n_591), .B1(n_788), .B2(n_789), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_483), .A2(n_1133), .B1(n_1134), .B2(n_1135), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1290 ( .A1(n_483), .A2(n_1133), .B1(n_1291), .B2(n_1292), .Y(n_1290) );
INVx5_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_488), .B1(n_489), .B2(n_491), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g601 ( .A(n_487), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_487), .A2(n_701), .B1(n_713), .B2(n_722), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g1781 ( .A1(n_487), .A2(n_661), .B1(n_1770), .B2(n_1774), .Y(n_1781) );
OAI211xp5_ASAP7_75t_SL g1381 ( .A1(n_489), .A2(n_1382), .B(n_1383), .C(n_1386), .Y(n_1381) );
BUFx4f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx4_ASAP7_75t_L g652 ( .A(n_490), .Y(n_652) );
BUFx4f_ASAP7_75t_L g661 ( .A(n_490), .Y(n_661) );
BUFx4f_ASAP7_75t_L g720 ( .A(n_490), .Y(n_720) );
BUFx4f_ASAP7_75t_L g752 ( .A(n_490), .Y(n_752) );
BUFx6f_ASAP7_75t_L g1039 ( .A(n_490), .Y(n_1039) );
OR2x6_ASAP7_75t_L g1689 ( .A(n_490), .B(n_1690), .Y(n_1689) );
OAI22xp5_ASAP7_75t_SL g588 ( .A1(n_492), .A2(n_589), .B1(n_590), .B2(n_599), .Y(n_588) );
OAI33xp33_ASAP7_75t_L g904 ( .A1(n_492), .A2(n_905), .A3(n_906), .B1(n_910), .B2(n_914), .B3(n_916), .Y(n_904) );
OAI33xp33_ASAP7_75t_L g1123 ( .A1(n_492), .A2(n_781), .A3(n_1124), .B1(n_1128), .B2(n_1132), .B3(n_1136), .Y(n_1123) );
OAI33xp33_ASAP7_75t_L g1286 ( .A1(n_492), .A2(n_905), .A3(n_1287), .B1(n_1290), .B2(n_1293), .B3(n_1296), .Y(n_1286) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g794 ( .A(n_493), .Y(n_794) );
AOI33xp33_ASAP7_75t_L g958 ( .A1(n_493), .A2(n_959), .A3(n_960), .B1(n_964), .B2(n_971), .B3(n_972), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g1703 ( .A(n_493), .B(n_1704), .C(n_1707), .Y(n_1703) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g1378 ( .A1(n_494), .A2(n_911), .B1(n_1090), .B2(n_1379), .C(n_1380), .Y(n_1378) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_498), .A2(n_821), .B1(n_833), .B2(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g796 ( .A(n_499), .Y(n_796) );
INVx3_ASAP7_75t_L g1126 ( .A(n_499), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g646 ( .A(n_500), .Y(n_646) );
INVx3_ASAP7_75t_L g909 ( .A(n_500), .Y(n_909) );
OAI33xp33_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_507), .A3(n_514), .B1(n_520), .B2(n_525), .B3(n_531), .Y(n_503) );
BUFx4f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx4f_ASAP7_75t_L g536 ( .A(n_505), .Y(n_536) );
BUFx8_ASAP7_75t_L g802 ( .A(n_505), .Y(n_802) );
BUFx2_ASAP7_75t_L g888 ( .A(n_505), .Y(n_888) );
BUFx2_ASAP7_75t_L g1727 ( .A(n_506), .Y(n_1727) );
BUFx4f_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_509), .A2(n_699), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_SL g541 ( .A(n_510), .Y(n_541) );
OAI22xp33_ASAP7_75t_L g901 ( .A1(n_511), .A2(n_804), .B1(n_902), .B2(n_903), .Y(n_901) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g848 ( .A(n_513), .Y(n_848) );
INVx1_ASAP7_75t_L g1304 ( .A(n_513), .Y(n_1304) );
OR2x6_ASAP7_75t_L g1720 ( .A(n_513), .B(n_1721), .Y(n_1720) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_515), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g1047 ( .A1(n_515), .A2(n_548), .B1(n_1036), .B2(n_1043), .Y(n_1047) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
INVx5_ASAP7_75t_L g521 ( .A(n_516), .Y(n_521) );
INVx2_ASAP7_75t_SL g546 ( .A(n_516), .Y(n_546) );
INVx3_ASAP7_75t_L g636 ( .A(n_516), .Y(n_636) );
HB1xp67_ASAP7_75t_L g1330 ( .A(n_516), .Y(n_1330) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_517), .A2(n_825), .B1(n_826), .B2(n_827), .Y(n_824) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g633 ( .A(n_519), .Y(n_633) );
BUFx3_ASAP7_75t_L g826 ( .A(n_521), .Y(n_826) );
INVx8_ASAP7_75t_L g1726 ( .A(n_521), .Y(n_1726) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_522), .A2(n_829), .B1(n_830), .B2(n_831), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_522), .A2(n_826), .B1(n_894), .B2(n_895), .Y(n_893) );
OAI22xp33_ASAP7_75t_SL g1146 ( .A1(n_522), .A2(n_1131), .B1(n_1139), .B2(n_1147), .Y(n_1146) );
OAI22xp33_ASAP7_75t_L g1305 ( .A1(n_522), .A2(n_1291), .B1(n_1299), .B2(n_1306), .Y(n_1305) );
OAI221xp5_ASAP7_75t_L g1406 ( .A1(n_522), .A2(n_1377), .B1(n_1382), .B2(n_1407), .C(n_1408), .Y(n_1406) );
CKINVDCx8_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
INVx3_ASAP7_75t_L g548 ( .A(n_523), .Y(n_548) );
INVx3_ASAP7_75t_L g706 ( .A(n_523), .Y(n_706) );
INVx3_ASAP7_75t_L g710 ( .A(n_523), .Y(n_710) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g554 ( .A(n_524), .Y(n_554) );
OAI33xp33_ASAP7_75t_L g801 ( .A1(n_525), .A2(n_802), .A3(n_803), .B1(n_806), .B2(n_810), .B3(n_811), .Y(n_801) );
OAI33xp33_ASAP7_75t_L g819 ( .A1(n_525), .A2(n_802), .A3(n_820), .B1(n_824), .B2(n_828), .B3(n_832), .Y(n_819) );
OAI33xp33_ASAP7_75t_L g887 ( .A1(n_525), .A2(n_888), .A3(n_889), .B1(n_893), .B2(n_896), .B3(n_901), .Y(n_887) );
INVx1_ASAP7_75t_L g957 ( .A(n_525), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_525), .A2(n_888), .B1(n_1401), .B2(n_1406), .Y(n_1400) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g1148 ( .A(n_526), .Y(n_1148) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g558 ( .A(n_527), .Y(n_558) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g1671 ( .A(n_529), .Y(n_1671) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_529), .B(n_1665), .Y(n_1678) );
INVx1_ASAP7_75t_L g619 ( .A(n_532), .Y(n_619) );
NOR4xp25_ASAP7_75t_L g533 ( .A(n_534), .B(n_564), .C(n_588), .D(n_604), .Y(n_533) );
OAI33xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_537), .A3(n_544), .B1(n_549), .B2(n_556), .B3(n_559), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI33xp33_ASAP7_75t_L g625 ( .A1(n_536), .A2(n_626), .A3(n_630), .B1(n_635), .B2(n_639), .B3(n_642), .Y(n_625) );
OAI33xp33_ASAP7_75t_L g696 ( .A1(n_536), .A2(n_642), .A3(n_697), .B1(n_702), .B2(n_707), .B3(n_711), .Y(n_696) );
OAI33xp33_ASAP7_75t_L g989 ( .A1(n_536), .A2(n_642), .A3(n_990), .B1(n_993), .B2(n_996), .B3(n_1001), .Y(n_989) );
OAI33xp33_ASAP7_75t_L g1044 ( .A1(n_536), .A2(n_642), .A3(n_1045), .B1(n_1046), .B2(n_1047), .B3(n_1048), .Y(n_1044) );
OAI33xp33_ASAP7_75t_L g1255 ( .A1(n_536), .A2(n_642), .A3(n_1256), .B1(n_1257), .B2(n_1258), .B3(n_1259), .Y(n_1255) );
OAI22xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_542), .B2(n_543), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_541), .A2(n_560), .B1(n_561), .B2(n_563), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g1001 ( .A1(n_541), .A2(n_562), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
OAI22xp33_ASAP7_75t_L g1045 ( .A1(n_541), .A2(n_543), .B1(n_1031), .B2(n_1038), .Y(n_1045) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_541), .A2(n_562), .B1(n_1033), .B2(n_1040), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1256 ( .A1(n_541), .A2(n_562), .B1(n_1244), .B2(n_1250), .Y(n_1256) );
OAI22xp33_ASAP7_75t_L g626 ( .A1(n_543), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_543), .A2(n_804), .B1(n_1081), .B2(n_1082), .Y(n_1080) );
INVx1_ASAP7_75t_L g1273 ( .A(n_543), .Y(n_1273) );
OAI22xp33_ASAP7_75t_L g1309 ( .A1(n_543), .A2(n_1142), .B1(n_1289), .B2(n_1295), .Y(n_1309) );
OAI22xp33_ASAP7_75t_L g1776 ( .A1(n_543), .A2(n_628), .B1(n_1777), .B2(n_1778), .Y(n_1776) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_547), .B2(n_548), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g1772 ( .A1(n_548), .A2(n_1773), .B1(n_1774), .B2(n_1775), .Y(n_1772) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_552), .B1(n_553), .B2(n_555), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_SL g632 ( .A(n_551), .Y(n_632) );
INVx3_ASAP7_75t_L g1076 ( .A(n_551), .Y(n_1076) );
INVx3_ASAP7_75t_L g1773 ( .A(n_551), .Y(n_1773) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_553), .A2(n_636), .B1(n_637), .B2(n_638), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_553), .A2(n_946), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_553), .A2(n_1076), .B1(n_1077), .B2(n_1078), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1769 ( .A1(n_553), .A2(n_1407), .B1(n_1770), .B2(n_1771), .Y(n_1769) );
BUFx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_L g1340 ( .A(n_558), .Y(n_1340) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_562), .A2(n_628), .B1(n_640), .B2(n_641), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_562), .A2(n_628), .B1(n_712), .B2(n_713), .Y(n_711) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_562), .Y(n_805) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_562), .Y(n_823) );
AOI31xp33_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_569), .A3(n_577), .B(n_587), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_567), .B(n_1423), .Y(n_1422) );
AND2x4_ASAP7_75t_SL g1752 ( .A(n_567), .B(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g879 ( .A(n_576), .Y(n_879) );
INVx2_ASAP7_75t_L g1282 ( .A(n_576), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_583), .B2(n_584), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_578), .A2(n_583), .B1(n_614), .B2(n_615), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g1797 ( .A1(n_579), .A2(n_1798), .B1(n_1799), .B2(n_1800), .Y(n_1797) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_580), .Y(n_603) );
INVx3_ASAP7_75t_L g1220 ( .A(n_580), .Y(n_1220) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g595 ( .A(n_581), .Y(n_595) );
AND2x2_ASAP7_75t_L g1664 ( .A(n_581), .B(n_1665), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g1672 ( .A(n_581), .B(n_1673), .Y(n_1672) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g1372 ( .A(n_586), .B(n_1373), .Y(n_1372) );
AO21x1_ASAP7_75t_L g976 ( .A1(n_587), .A2(n_977), .B(n_978), .Y(n_976) );
AO21x1_ASAP7_75t_L g1193 ( .A1(n_587), .A2(n_1194), .B(n_1198), .Y(n_1193) );
OAI33xp33_ASAP7_75t_L g644 ( .A1(n_589), .A2(n_645), .A3(n_648), .B1(n_653), .B2(n_654), .B3(n_657), .Y(n_644) );
OAI33xp33_ASAP7_75t_L g1004 ( .A1(n_589), .A2(n_1005), .A3(n_1006), .B1(n_1008), .B2(n_1010), .B3(n_1011), .Y(n_1004) );
OAI33xp33_ASAP7_75t_L g1779 ( .A1(n_589), .A2(n_657), .A3(n_1780), .B1(n_1781), .B2(n_1782), .B3(n_1783), .Y(n_1779) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g912 ( .A(n_592), .Y(n_912) );
INVx2_ASAP7_75t_L g1007 ( .A(n_592), .Y(n_1007) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g961 ( .A(n_595), .Y(n_961) );
INVx2_ASAP7_75t_SL g973 ( .A(n_595), .Y(n_973) );
INVx2_ASAP7_75t_L g1212 ( .A(n_595), .Y(n_1212) );
INVx2_ASAP7_75t_L g1387 ( .A(n_595), .Y(n_1387) );
BUFx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g1706 ( .A(n_597), .Y(n_1706) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx3_ASAP7_75t_L g963 ( .A(n_598), .Y(n_963) );
INVx2_ASAP7_75t_L g975 ( .A(n_598), .Y(n_975) );
BUFx3_ASAP7_75t_L g1687 ( .A(n_598), .Y(n_1687) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI31xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_611), .A3(n_613), .B(n_616), .Y(n_604) );
INVx1_ASAP7_75t_L g1179 ( .A(n_607), .Y(n_1179) );
INVx2_ASAP7_75t_SL g1354 ( .A(n_612), .Y(n_1354) );
AOI22xp5_ASAP7_75t_L g1105 ( .A1(n_614), .A2(n_1106), .B1(n_1107), .B2(n_1108), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_614), .A2(n_615), .B1(n_1345), .B2(n_1346), .Y(n_1357) );
INVx1_ASAP7_75t_L g766 ( .A(n_615), .Y(n_766) );
INVx2_ASAP7_75t_L g928 ( .A(n_615), .Y(n_928) );
AO21x1_ASAP7_75t_L g921 ( .A1(n_616), .A2(n_922), .B(n_925), .Y(n_921) );
AOI31xp33_ASAP7_75t_L g1094 ( .A1(n_616), .A2(n_1095), .A3(n_1102), .B(n_1105), .Y(n_1094) );
CKINVDCx14_ASAP7_75t_R g616 ( .A(n_617), .Y(n_616) );
OAI31xp33_ASAP7_75t_L g1269 ( .A1(n_617), .A2(n_1270), .A3(n_1271), .B(n_1277), .Y(n_1269) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
XNOR2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_693), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_659), .C(n_677), .Y(n_623) );
NOR2xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_644), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_627), .A2(n_640), .B1(n_646), .B2(n_647), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_628), .A2(n_698), .B1(n_699), .B2(n_701), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_628), .A2(n_699), .B1(n_991), .B2(n_992), .Y(n_990) );
OAI22xp33_ASAP7_75t_L g1259 ( .A1(n_628), .A2(n_834), .B1(n_1245), .B2(n_1251), .Y(n_1259) );
OAI22xp33_ASAP7_75t_L g1766 ( .A1(n_628), .A2(n_1394), .B1(n_1767), .B2(n_1768), .Y(n_1766) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_629), .A2(n_641), .B1(n_649), .B2(n_651), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_631), .A2(n_637), .B1(n_649), .B2(n_651), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_633), .A2(n_997), .B1(n_998), .B2(n_1000), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_634), .A2(n_638), .B1(n_647), .B2(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g898 ( .A(n_636), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_636), .A2(n_706), .B1(n_1247), .B2(n_1253), .Y(n_1257) );
INVx3_ASAP7_75t_L g1730 ( .A(n_643), .Y(n_1730) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_646), .A2(n_717), .B1(n_991), .B2(n_1002), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_646), .A2(n_647), .B1(n_995), .B2(n_1000), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_646), .A2(n_1031), .B1(n_1032), .B2(n_1033), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_646), .A2(n_717), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1243 ( .A1(n_646), .A2(n_717), .B1(n_1244), .B2(n_1245), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_646), .A2(n_1032), .B1(n_1253), .B2(n_1254), .Y(n_1252) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_647), .A2(n_705), .B1(n_709), .B2(n_716), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g1780 ( .A1(n_647), .A2(n_716), .B1(n_1767), .B2(n_1777), .Y(n_1780) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_649), .A2(n_703), .B1(n_708), .B2(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g1133 ( .A(n_650), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_651), .A2(n_994), .B1(n_997), .B2(n_1007), .Y(n_1006) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g722 ( .A(n_652), .Y(n_722) );
INVx2_ASAP7_75t_L g913 ( .A(n_652), .Y(n_913) );
INVx1_ASAP7_75t_L g915 ( .A(n_652), .Y(n_915) );
INVx1_ASAP7_75t_L g1090 ( .A(n_652), .Y(n_1090) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g1011 ( .A(n_658), .Y(n_1011) );
AOI33xp33_ASAP7_75t_L g1210 ( .A1(n_658), .A2(n_1086), .A3(n_1211), .B1(n_1213), .B2(n_1217), .B3(n_1218), .Y(n_1210) );
NAND3xp33_ASAP7_75t_L g1325 ( .A(n_658), .B(n_1326), .C(n_1327), .Y(n_1325) );
OAI31xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_672), .A3(n_675), .B(n_676), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g1343 ( .A(n_662), .B(n_1344), .C(n_1347), .Y(n_1343) );
NAND3xp33_ASAP7_75t_SL g1794 ( .A(n_662), .B(n_1795), .C(n_1797), .Y(n_1794) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g1205 ( .A(n_663), .Y(n_1205) );
INVx1_ASAP7_75t_L g1204 ( .A(n_664), .Y(n_1204) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx2_ASAP7_75t_L g970 ( .A(n_665), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_668), .A2(n_870), .B1(n_879), .B2(n_880), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_668), .A2(n_1275), .B1(n_1281), .B2(n_1282), .Y(n_1280) );
AOI222xp33_ASAP7_75t_L g1795 ( .A1(n_668), .A2(n_731), .B1(n_1321), .B2(n_1790), .C1(n_1791), .C2(n_1796), .Y(n_1795) );
AOI32xp33_ASAP7_75t_L g680 ( .A1(n_669), .A2(n_681), .A3(n_684), .B1(n_686), .B2(n_687), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_670), .A2(n_1015), .B1(n_1016), .B2(n_1017), .Y(n_1014) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g1196 ( .A(n_673), .Y(n_1196) );
BUFx3_ASAP7_75t_L g716 ( .A(n_674), .Y(n_716) );
BUFx3_ASAP7_75t_L g784 ( .A(n_674), .Y(n_784) );
INVx2_ASAP7_75t_SL g1298 ( .A(n_674), .Y(n_1298) );
BUFx6f_ASAP7_75t_L g1784 ( .A(n_674), .Y(n_1784) );
OAI31xp33_ASAP7_75t_L g748 ( .A1(n_676), .A2(n_749), .A3(n_758), .B(n_762), .Y(n_748) );
OAI31xp33_ASAP7_75t_L g1012 ( .A1(n_676), .A2(n_1013), .A3(n_1018), .B(n_1019), .Y(n_1012) );
OAI31xp33_ASAP7_75t_L g1049 ( .A1(n_676), .A2(n_1050), .A3(n_1054), .B(n_1055), .Y(n_1049) );
INVx1_ASAP7_75t_L g1117 ( .A(n_676), .Y(n_1117) );
OAI31xp33_ASAP7_75t_L g1151 ( .A1(n_676), .A2(n_1152), .A3(n_1156), .B(n_1158), .Y(n_1151) );
OAI31xp33_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_679), .A3(n_689), .B(n_692), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_681), .A2(n_729), .B1(n_741), .B2(n_742), .Y(n_740) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_682), .B(n_1715), .Y(n_1714) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x6_ASAP7_75t_L g1718 ( .A(n_684), .B(n_1715), .Y(n_1718) );
INVx3_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_L g739 ( .A(n_686), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_686), .A2(n_742), .B1(n_1016), .B2(n_1024), .Y(n_1023) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_686), .A2(n_742), .B1(n_1052), .B2(n_1060), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_686), .A2(n_742), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_686), .A2(n_742), .B1(n_1230), .B2(n_1239), .Y(n_1238) );
INVxp67_ASAP7_75t_L g1396 ( .A(n_686), .Y(n_1396) );
AOI222xp33_ASAP7_75t_L g1787 ( .A1(n_686), .A2(n_742), .B1(n_1788), .B2(n_1789), .C1(n_1790), .C2(n_1791), .Y(n_1787) );
NAND3xp33_ASAP7_75t_L g1355 ( .A(n_688), .B(n_1356), .C(n_1357), .Y(n_1355) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_691), .A2(n_874), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
OAI31xp33_ASAP7_75t_SL g735 ( .A1(n_692), .A2(n_736), .A3(n_737), .B(n_738), .Y(n_735) );
OAI31xp33_ASAP7_75t_SL g1020 ( .A1(n_692), .A2(n_1021), .A3(n_1022), .B(n_1025), .Y(n_1020) );
OAI31xp33_ASAP7_75t_SL g1056 ( .A1(n_692), .A2(n_1057), .A3(n_1058), .B(n_1061), .Y(n_1056) );
OAI21xp5_ASAP7_75t_L g1352 ( .A1(n_692), .A2(n_1353), .B(n_1355), .Y(n_1352) );
OAI21xp5_ASAP7_75t_L g1785 ( .A1(n_692), .A2(n_1786), .B(n_1792), .Y(n_1785) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_724), .C(n_735), .Y(n_694) );
NOR2xp33_ASAP7_75t_SL g695 ( .A(n_696), .B(n_714), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_698), .A2(n_712), .B1(n_716), .B2(n_717), .Y(n_715) );
INVx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g892 ( .A(n_700), .Y(n_892) );
INVx2_ASAP7_75t_L g1150 ( .A(n_700), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_704), .A2(n_789), .B1(n_800), .B2(n_809), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_704), .A2(n_706), .B1(n_994), .B2(n_995), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_704), .A2(n_706), .B1(n_1035), .B2(n_1042), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_704), .A2(n_710), .B1(n_1248), .B2(n_1254), .Y(n_1258) );
OAI22xp5_ASAP7_75t_L g1783 ( .A1(n_717), .A2(n_1771), .B1(n_1775), .B2(n_1784), .Y(n_1783) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_720), .A2(n_1007), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
INVx1_ASAP7_75t_L g1800 ( .A(n_726), .Y(n_1800) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_731), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_731), .A2(n_1015), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
INVx1_ASAP7_75t_L g1395 ( .A(n_742), .Y(n_1395) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_815), .B2(n_816), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_763), .C(n_779), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g1128 ( .A1(n_752), .A2(n_1129), .B1(n_1130), .B2(n_1131), .Y(n_1128) );
OAI22xp5_ASAP7_75t_L g1293 ( .A1(n_752), .A2(n_1133), .B1(n_1294), .B2(n_1295), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_756), .A2(n_770), .B1(n_772), .B2(n_773), .Y(n_769) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_SL g883 ( .A(n_761), .Y(n_883) );
OAI31xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_767), .A3(n_774), .B(n_778), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g811 ( .A1(n_768), .A2(n_785), .B1(n_793), .B2(n_812), .Y(n_811) );
BUFx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
BUFx3_ASAP7_75t_L g850 ( .A(n_771), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_773), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_773), .A2(n_850), .B1(n_870), .B2(n_871), .Y(n_869) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g875 ( .A(n_778), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g1390 ( .A1(n_778), .A2(n_1391), .B(n_1400), .Y(n_1390) );
NOR2xp33_ASAP7_75t_SL g779 ( .A(n_780), .B(n_801), .Y(n_779) );
OAI33xp33_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .A3(n_787), .B1(n_790), .B2(n_794), .B3(n_795), .Y(n_780) );
INVx2_ASAP7_75t_SL g1086 ( .A(n_781), .Y(n_1086) );
INVx2_ASAP7_75t_SL g1324 ( .A(n_781), .Y(n_1324) );
OAI22xp33_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_782) );
OAI22xp33_ASAP7_75t_L g803 ( .A1(n_783), .A2(n_792), .B1(n_804), .B2(n_805), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_784), .A2(n_786), .B1(n_827), .B2(n_831), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_784), .A2(n_1137), .B1(n_1138), .B2(n_1139), .Y(n_1136) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_786), .A2(n_890), .B1(n_902), .B2(n_907), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_786), .A2(n_895), .B1(n_900), .B2(n_907), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_788), .A2(n_797), .B1(n_807), .B2(n_809), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_797), .B1(n_798), .B2(n_800), .Y(n_795) );
BUFx3_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OAI33xp33_ASAP7_75t_L g1140 ( .A1(n_802), .A2(n_1141), .A3(n_1144), .B1(n_1146), .B2(n_1148), .B3(n_1149), .Y(n_1140) );
OAI22xp33_ASAP7_75t_L g820 ( .A1(n_804), .A2(n_821), .B1(n_822), .B2(n_823), .Y(n_820) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_804), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g889 ( .A1(n_804), .A2(n_890), .B1(n_891), .B2(n_892), .Y(n_889) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_809), .A2(n_897), .B1(n_899), .B2(n_900), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_809), .A2(n_1129), .B1(n_1137), .B2(n_1145), .Y(n_1144) );
OAI22xp5_ASAP7_75t_L g1308 ( .A1(n_809), .A2(n_1145), .B1(n_1292), .B2(n_1300), .Y(n_1308) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g1143 ( .A(n_814), .Y(n_1143) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_842), .C(n_854), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_836), .Y(n_818) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g1261 ( .A(n_861), .Y(n_1261) );
XNOR2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_981), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_864), .B1(n_917), .B2(n_918), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
NAND3xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_876), .C(n_886), .Y(n_865) );
OAI31xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .A3(n_872), .B(n_875), .Y(n_866) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OAI31xp33_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_881), .A3(n_884), .B(n_885), .Y(n_876) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_904), .Y(n_886) );
OAI33xp33_ASAP7_75t_L g1068 ( .A1(n_888), .A2(n_1069), .A3(n_1072), .B1(n_1075), .B2(n_1079), .B3(n_1080), .Y(n_1068) );
OAI33xp33_ASAP7_75t_L g1301 ( .A1(n_888), .A2(n_1148), .A3(n_1302), .B1(n_1305), .B2(n_1308), .B3(n_1309), .Y(n_1301) );
OAI33xp33_ASAP7_75t_L g1765 ( .A1(n_888), .A2(n_1079), .A3(n_1766), .B1(n_1769), .B2(n_1772), .B3(n_1776), .Y(n_1765) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_891), .A2(n_903), .B1(n_911), .B2(n_915), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_894), .A2(n_899), .B1(n_911), .B2(n_913), .Y(n_910) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx2_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_911), .A2(n_1071), .B1(n_1082), .B2(n_1090), .Y(n_1091) );
INVx4_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NAND4xp25_ASAP7_75t_SL g920 ( .A(n_921), .B(n_931), .C(n_958), .D(n_976), .Y(n_920) );
AOI33xp33_ASAP7_75t_L g931 ( .A1(n_932), .A2(n_935), .A3(n_944), .B1(n_951), .B2(n_954), .B3(n_957), .Y(n_931) );
BUFx3_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_L g1176 ( .A(n_933), .Y(n_1176) );
NAND3xp33_ASAP7_75t_L g1328 ( .A(n_933), .B(n_1329), .C(n_1332), .Y(n_1328) );
AOI22xp33_ASAP7_75t_SL g1708 ( .A1(n_934), .A2(n_1709), .B1(n_1745), .B2(n_1749), .Y(n_1708) );
BUFx2_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g1178 ( .A1(n_938), .A2(n_1179), .B1(n_1180), .B2(n_1181), .C(n_1182), .Y(n_1178) );
INVx2_ASAP7_75t_SL g938 ( .A(n_939), .Y(n_938) );
BUFx3_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx8_ASAP7_75t_L g1174 ( .A(n_940), .Y(n_1174) );
BUFx3_ASAP7_75t_L g1335 ( .A(n_940), .Y(n_1335) );
NAND2x1p5_ASAP7_75t_L g1744 ( .A(n_940), .B(n_1715), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_942), .B(n_1187), .Y(n_1186) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g1336 ( .A(n_943), .Y(n_1336) );
INVx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
BUFx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g955 ( .A(n_947), .Y(n_955) );
INVx3_ASAP7_75t_L g999 ( .A(n_947), .Y(n_999) );
BUFx2_ASAP7_75t_L g1407 ( .A(n_947), .Y(n_1407) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx2_ASAP7_75t_L g956 ( .A(n_949), .Y(n_956) );
INVx5_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
BUFx3_ASAP7_75t_L g1331 ( .A(n_950), .Y(n_1331) );
BUFx12f_ASAP7_75t_L g1339 ( .A(n_950), .Y(n_1339) );
BUFx2_ASAP7_75t_L g1405 ( .A(n_950), .Y(n_1405) );
BUFx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g1739 ( .A1(n_953), .A2(n_1661), .B1(n_1702), .B2(n_1740), .Y(n_1739) );
HB1xp67_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx2_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx3_ASAP7_75t_L g1679 ( .A(n_975), .Y(n_1679) );
XOR2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_1062), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
XNOR2x1_ASAP7_75t_L g984 ( .A(n_985), .B(n_1026), .Y(n_984) );
XNOR2xp5_ASAP7_75t_L g985 ( .A(n_986), .B(n_987), .Y(n_985) );
AND3x1_ASAP7_75t_L g987 ( .A(n_988), .B(n_1012), .C(n_1020), .Y(n_987) );
NOR2xp33_ASAP7_75t_SL g988 ( .A(n_989), .B(n_1004), .Y(n_988) );
INVx2_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g1145 ( .A(n_999), .Y(n_1145) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_1007), .A2(n_1038), .B1(n_1039), .B2(n_1040), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_1007), .A2(n_1039), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
OAI22xp5_ASAP7_75t_SL g1089 ( .A1(n_1009), .A2(n_1073), .B1(n_1077), .B2(n_1090), .Y(n_1089) );
OAI33xp33_ASAP7_75t_L g1084 ( .A1(n_1011), .A2(n_1085), .A3(n_1087), .B1(n_1089), .B2(n_1091), .B3(n_1092), .Y(n_1084) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1015), .Y(n_1367) );
AND3x1_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1049), .C(n_1056), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1044), .Y(n_1028) );
OAI22xp33_ASAP7_75t_L g1124 ( .A1(n_1032), .A2(n_1125), .B1(n_1126), .B2(n_1127), .Y(n_1124) );
OAI22xp5_ASAP7_75t_L g1782 ( .A1(n_1039), .A2(n_1133), .B1(n_1768), .B2(n_1778), .Y(n_1782) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_1063), .A2(n_1064), .B1(n_1168), .B2(n_1260), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g1064 ( .A1(n_1065), .A2(n_1119), .B1(n_1120), .B2(n_1167), .Y(n_1064) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1065), .Y(n_1167) );
INVxp67_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
NOR4xp25_ASAP7_75t_L g1118 ( .A(n_1068), .B(n_1084), .C(n_1094), .D(n_1109), .Y(n_1118) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1076), .Y(n_1732) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1079), .Y(n_1182) );
INVxp67_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVxp67_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVxp67_ASAP7_75t_SL g1096 ( .A(n_1097), .Y(n_1096) );
AOI31xp67_ASAP7_75t_SL g1109 ( .A1(n_1110), .A2(n_1113), .A3(n_1115), .B(n_1117), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVxp67_ASAP7_75t_SL g1115 ( .A(n_1116), .Y(n_1115) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
NAND3xp33_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1151), .C(n_1159), .Y(n_1121) );
NOR2xp33_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1140), .Y(n_1122) );
OAI22xp33_ASAP7_75t_L g1149 ( .A1(n_1127), .A2(n_1135), .B1(n_1142), .B2(n_1150), .Y(n_1149) );
OAI22xp33_ASAP7_75t_L g1302 ( .A1(n_1142), .A2(n_1288), .B1(n_1294), .B2(n_1303), .Y(n_1302) );
INVx2_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1168), .Y(n_1260) );
XNOR2x1_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1224), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1206), .Y(n_1169) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1171), .Y(n_1208) );
AOI21xp5_ASAP7_75t_L g1171 ( .A1(n_1172), .A2(n_1175), .B(n_1177), .Y(n_1171) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx8_ASAP7_75t_L g1724 ( .A(n_1174), .Y(n_1724) );
INVx3_ASAP7_75t_L g1740 ( .A(n_1174), .Y(n_1740) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1183), .B(n_1193), .Y(n_1207) );
OAI31xp33_ASAP7_75t_SL g1183 ( .A1(n_1184), .A2(n_1185), .A3(n_1191), .B(n_1192), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1202 ( .A(n_1190), .B(n_1203), .Y(n_1202) );
OAI31xp33_ASAP7_75t_SL g1233 ( .A1(n_1192), .A2(n_1234), .A3(n_1235), .B(n_1240), .Y(n_1233) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1199), .B(n_1200), .Y(n_1198) );
NAND3xp33_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .C(n_1205), .Y(n_1200) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
OAI31xp33_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1208), .A3(n_1209), .B(n_1221), .Y(n_1206) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1210), .Y(n_1223) );
BUFx6f_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1215), .B(n_1665), .Y(n_1748) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1220), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
NAND3xp33_ASAP7_75t_SL g1225 ( .A(n_1226), .B(n_1233), .C(n_1241), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1231), .B(n_1237), .Y(n_1236) );
NOR2xp33_ASAP7_75t_L g1241 ( .A(n_1242), .B(n_1255), .Y(n_1241) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1266), .B1(n_1359), .B2(n_1409), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_1267), .A2(n_1312), .B1(n_1313), .B2(n_1358), .Y(n_1266) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1267), .Y(n_1358) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1268), .Y(n_1310) );
NAND3xp33_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1278), .C(n_1285), .Y(n_1268) );
INVx2_ASAP7_75t_SL g1272 ( .A(n_1273), .Y(n_1272) );
NOR2xp33_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1301), .Y(n_1285) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
OAI211xp5_ASAP7_75t_L g1401 ( .A1(n_1306), .A2(n_1402), .B(n_1403), .C(n_1404), .Y(n_1401) );
INVx2_ASAP7_75t_SL g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
NAND3xp33_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1342), .C(n_1352), .Y(n_1314) );
AND4x1_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1325), .C(n_1328), .D(n_1337), .Y(n_1315) );
NAND3xp33_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1322), .C(n_1324), .Y(n_1316) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
NAND3xp33_ASAP7_75t_L g1337 ( .A(n_1338), .B(n_1340), .C(n_1341), .Y(n_1337) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1359), .Y(n_1409) );
HB1xp67_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
OAI21xp5_ASAP7_75t_L g1361 ( .A1(n_1362), .A2(n_1388), .B(n_1390), .Y(n_1361) );
OAI21xp5_ASAP7_75t_L g1374 ( .A1(n_1375), .A2(n_1378), .B(n_1381), .Y(n_1374) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
BUFx2_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
NAND2xp5_ASAP7_75t_SL g1391 ( .A(n_1392), .B(n_1398), .Y(n_1391) );
BUFx2_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
BUFx4f_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
INVx3_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
OR2x2_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1421), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
NOR2xp33_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1419), .Y(n_1416) );
NOR2xp33_ASAP7_75t_L g1759 ( .A(n_1417), .B(n_1420), .Y(n_1759) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1417), .Y(n_1806) );
HB1xp67_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
NOR2xp33_ASAP7_75t_L g1808 ( .A(n_1420), .B(n_1806), .Y(n_1808) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
OAI221xp5_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1653), .B1(n_1655), .B2(n_1751), .C(n_1754), .Y(n_1424) );
AND5x1_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1567), .C(n_1614), .D(n_1636), .E(n_1649), .Y(n_1425) );
OAI31xp33_ASAP7_75t_L g1426 ( .A1(n_1427), .A2(n_1505), .A3(n_1544), .B(n_1558), .Y(n_1426) );
OAI221xp5_ASAP7_75t_L g1427 ( .A1(n_1428), .A2(n_1456), .B1(n_1467), .B2(n_1474), .C(n_1475), .Y(n_1427) );
NAND2x1_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1444), .Y(n_1428) );
NAND2xp5_ASAP7_75t_SL g1520 ( .A(n_1429), .B(n_1521), .Y(n_1520) );
CKINVDCx5p33_ASAP7_75t_R g1541 ( .A(n_1429), .Y(n_1541) );
OAI21xp33_ASAP7_75t_L g1581 ( .A1(n_1429), .A2(n_1494), .B(n_1582), .Y(n_1581) );
NOR2xp33_ASAP7_75t_L g1587 ( .A(n_1429), .B(n_1588), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1429), .B(n_1497), .Y(n_1591) );
NOR2x1_ASAP7_75t_L g1596 ( .A(n_1429), .B(n_1597), .Y(n_1596) );
OAI22xp5_ASAP7_75t_SL g1619 ( .A1(n_1429), .A2(n_1575), .B1(n_1620), .B2(n_1624), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1429), .B(n_1648), .Y(n_1647) );
INVx4_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
INVx4_ASAP7_75t_L g1468 ( .A(n_1430), .Y(n_1468) );
OR2x2_ASAP7_75t_L g1501 ( .A(n_1430), .B(n_1445), .Y(n_1501) );
NAND2xp5_ASAP7_75t_SL g1503 ( .A(n_1430), .B(n_1445), .Y(n_1503) );
NOR2xp33_ASAP7_75t_L g1534 ( .A(n_1430), .B(n_1535), .Y(n_1534) );
NOR3xp33_ASAP7_75t_L g1555 ( .A(n_1430), .B(n_1556), .C(n_1557), .Y(n_1555) );
NOR2xp33_ASAP7_75t_L g1574 ( .A(n_1430), .B(n_1478), .Y(n_1574) );
NOR2xp33_ASAP7_75t_L g1599 ( .A(n_1430), .B(n_1600), .Y(n_1599) );
AND2x4_ASAP7_75t_SL g1430 ( .A(n_1431), .B(n_1439), .Y(n_1430) );
AND2x4_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1434), .Y(n_1432) );
AND2x6_ASAP7_75t_L g1437 ( .A(n_1433), .B(n_1438), .Y(n_1437) );
AND2x6_ASAP7_75t_L g1440 ( .A(n_1433), .B(n_1441), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1433), .B(n_1443), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1433), .B(n_1443), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1433), .B(n_1443), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1433), .B(n_1434), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1436), .Y(n_1434) );
INVx2_ASAP7_75t_L g1564 ( .A(n_1437), .Y(n_1564) );
HB1xp67_ASAP7_75t_L g1805 ( .A(n_1438), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1449), .Y(n_1444) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1445), .Y(n_1471) );
OR2x2_ASAP7_75t_L g1522 ( .A(n_1445), .B(n_1523), .Y(n_1522) );
OR2x2_ASAP7_75t_L g1579 ( .A(n_1445), .B(n_1450), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1445), .B(n_1453), .Y(n_1592) );
OR2x2_ASAP7_75t_L g1600 ( .A(n_1445), .B(n_1490), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1623 ( .A(n_1445), .B(n_1490), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1447), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1446), .B(n_1447), .Y(n_1488) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1449), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1449), .B(n_1550), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1453), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1450), .B(n_1473), .Y(n_1472) );
OR2x2_ASAP7_75t_L g1478 ( .A(n_1450), .B(n_1453), .Y(n_1478) );
INVx2_ASAP7_75t_L g1490 ( .A(n_1450), .Y(n_1490) );
AOI332xp33_ASAP7_75t_L g1533 ( .A1(n_1450), .A2(n_1488), .A3(n_1526), .B1(n_1534), .B2(n_1536), .B3(n_1539), .C1(n_1542), .C2(n_1543), .Y(n_1533) );
NAND2x1p5_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1452), .Y(n_1450) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1453), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1453), .B(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1453), .Y(n_1523) );
OR2x2_ASAP7_75t_L g1588 ( .A(n_1453), .B(n_1488), .Y(n_1588) );
NAND3xp33_ASAP7_75t_L g1632 ( .A(n_1453), .B(n_1458), .C(n_1559), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1454), .B(n_1455), .Y(n_1453) );
OAI21xp33_ASAP7_75t_L g1594 ( .A1(n_1456), .A2(n_1595), .B(n_1598), .Y(n_1594) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1462), .Y(n_1457) );
INVx3_ASAP7_75t_L g1481 ( .A(n_1458), .Y(n_1481) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1458), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1458), .B(n_1463), .Y(n_1546) );
OR2x2_ASAP7_75t_L g1557 ( .A(n_1458), .B(n_1463), .Y(n_1557) );
NOR2xp33_ASAP7_75t_SL g1608 ( .A(n_1458), .B(n_1560), .Y(n_1608) );
OAI322xp33_ASAP7_75t_L g1650 ( .A1(n_1458), .A2(n_1496), .A3(n_1499), .B1(n_1545), .B2(n_1579), .C1(n_1651), .C2(n_1652), .Y(n_1650) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1459), .B(n_1460), .Y(n_1458) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx2_ASAP7_75t_L g1474 ( .A(n_1463), .Y(n_1474) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_1463), .B(n_1483), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1463), .B(n_1481), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1463), .B(n_1497), .Y(n_1526) );
OR2x2_ASAP7_75t_L g1535 ( .A(n_1463), .B(n_1484), .Y(n_1535) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
OR2x2_ASAP7_75t_L g1495 ( .A(n_1464), .B(n_1483), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_1465), .B(n_1466), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1469), .Y(n_1467) );
CKINVDCx5p33_ASAP7_75t_R g1493 ( .A(n_1468), .Y(n_1493) );
NOR2xp33_ASAP7_75t_L g1507 ( .A(n_1468), .B(n_1508), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1468), .B(n_1513), .Y(n_1604) );
OR2x2_ASAP7_75t_L g1618 ( .A(n_1468), .B(n_1583), .Y(n_1618) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
OAI211xp5_ASAP7_75t_L g1615 ( .A1(n_1470), .A2(n_1552), .B(n_1573), .C(n_1616), .Y(n_1615) );
OR2x2_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1472), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1471), .B(n_1477), .Y(n_1476) );
NOR2xp33_ASAP7_75t_L g1510 ( .A(n_1471), .B(n_1490), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1471), .B(n_1489), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1471), .B(n_1596), .Y(n_1611) );
OR2x2_ASAP7_75t_L g1643 ( .A(n_1471), .B(n_1478), .Y(n_1643) );
OR2x2_ASAP7_75t_L g1502 ( .A(n_1472), .B(n_1503), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g1537 ( .A(n_1472), .B(n_1538), .Y(n_1537) );
OR2x2_ASAP7_75t_L g1583 ( .A(n_1472), .B(n_1488), .Y(n_1583) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1472), .Y(n_1648) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1474), .Y(n_1575) );
NAND2xp5_ASAP7_75t_L g1622 ( .A(n_1474), .B(n_1559), .Y(n_1622) );
AOI221xp5_ASAP7_75t_L g1475 ( .A1(n_1476), .A2(n_1479), .B1(n_1487), .B2(n_1491), .C(n_1498), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1476), .B(n_1493), .Y(n_1553) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1477), .B(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
OR2x2_ASAP7_75t_L g1528 ( .A(n_1478), .B(n_1501), .Y(n_1528) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
OR2x2_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1482), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1496 ( .A(n_1481), .B(n_1497), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1504 ( .A(n_1481), .B(n_1497), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1481), .B(n_1513), .Y(n_1512) );
OR2x2_ASAP7_75t_L g1532 ( .A(n_1481), .B(n_1495), .Y(n_1532) );
CKINVDCx14_ASAP7_75t_R g1593 ( .A(n_1481), .Y(n_1593) );
OR2x2_ASAP7_75t_L g1635 ( .A(n_1481), .B(n_1517), .Y(n_1635) );
CKINVDCx5p33_ASAP7_75t_R g1513 ( .A(n_1482), .Y(n_1513) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1483), .Y(n_1517) );
NOR2xp33_ASAP7_75t_L g1625 ( .A(n_1483), .B(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1484), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .Y(n_1484) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1487), .Y(n_1556) );
AOI22xp5_ASAP7_75t_L g1620 ( .A1(n_1487), .A2(n_1543), .B1(n_1621), .B2(n_1623), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1488), .B(n_1489), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_1488), .B(n_1574), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1489), .B(n_1500), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1489), .B(n_1531), .Y(n_1530) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1489), .Y(n_1538) );
OAI311xp33_ASAP7_75t_L g1569 ( .A1(n_1490), .A2(n_1493), .A3(n_1570), .B1(n_1571), .C1(n_1585), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1496), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1494), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1631 ( .A(n_1493), .B(n_1513), .Y(n_1631) );
O2A1O1Ixp33_ASAP7_75t_L g1649 ( .A1(n_1494), .A2(n_1572), .B(n_1637), .C(n_1650), .Y(n_1649) );
CKINVDCx5p33_ASAP7_75t_R g1494 ( .A(n_1495), .Y(n_1494) );
INVx2_ASAP7_75t_L g1552 ( .A(n_1497), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1497), .B(n_1541), .Y(n_1580) );
AOI21xp33_ASAP7_75t_L g1498 ( .A1(n_1499), .A2(n_1502), .B(n_1504), .Y(n_1498) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
NOR2xp33_ASAP7_75t_L g1606 ( .A(n_1502), .B(n_1552), .Y(n_1606) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1503), .Y(n_1550) );
O2A1O1Ixp33_ASAP7_75t_L g1609 ( .A1(n_1504), .A2(n_1543), .B(n_1610), .C(n_1612), .Y(n_1609) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1504), .Y(n_1641) );
OAI211xp5_ASAP7_75t_SL g1505 ( .A1(n_1506), .A2(n_1511), .B(n_1514), .C(n_1533), .Y(n_1505) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
HB1xp67_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
AOI211xp5_ASAP7_75t_L g1514 ( .A1(n_1515), .A2(n_1519), .B(n_1524), .C(n_1529), .Y(n_1514) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1518), .Y(n_1516) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1517), .Y(n_1548) );
O2A1O1Ixp33_ASAP7_75t_L g1605 ( .A1(n_1517), .A2(n_1574), .B(n_1582), .C(n_1606), .Y(n_1605) );
AOI211xp5_ASAP7_75t_L g1614 ( .A1(n_1518), .A2(n_1615), .B(n_1619), .C(n_1627), .Y(n_1614) );
INVxp67_ASAP7_75t_SL g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
INVxp67_ASAP7_75t_SL g1524 ( .A(n_1525), .Y(n_1524) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1527), .Y(n_1525) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1526), .B(n_1542), .Y(n_1584) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
AOI21xp33_ASAP7_75t_L g1644 ( .A1(n_1532), .A2(n_1645), .B(n_1646), .Y(n_1644) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1534), .Y(n_1651) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1535), .Y(n_1543) );
OR2x2_ASAP7_75t_L g1570 ( .A(n_1535), .B(n_1540), .Y(n_1570) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1541), .Y(n_1539) );
OAI21xp33_ASAP7_75t_SL g1638 ( .A1(n_1540), .A2(n_1639), .B(n_1640), .Y(n_1638) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1542), .Y(n_1628) );
OAI21xp33_ASAP7_75t_L g1633 ( .A1(n_1543), .A2(n_1617), .B(n_1634), .Y(n_1633) );
OAI211xp5_ASAP7_75t_L g1544 ( .A1(n_1545), .A2(n_1547), .B(n_1551), .C(n_1554), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
NAND2xp5_ASAP7_75t_L g1598 ( .A(n_1546), .B(n_1599), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1549), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1548), .B(n_1587), .Y(n_1586) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1548), .B(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1549), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1553), .Y(n_1551) );
NAND2xp5_ASAP7_75t_SL g1616 ( .A(n_1552), .B(n_1617), .Y(n_1616) );
OR2x2_ASAP7_75t_L g1629 ( .A(n_1552), .B(n_1557), .Y(n_1629) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1553), .Y(n_1645) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1558), .Y(n_1568) );
INVx2_ASAP7_75t_L g1558 ( .A(n_1559), .Y(n_1558) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
OAI221xp5_ASAP7_75t_L g1561 ( .A1(n_1562), .A2(n_1563), .B1(n_1564), .B2(n_1565), .C(n_1566), .Y(n_1561) );
CKINVDCx20_ASAP7_75t_R g1654 ( .A(n_1564), .Y(n_1654) );
AOI211xp5_ASAP7_75t_L g1567 ( .A1(n_1568), .A2(n_1569), .B(n_1601), .C(n_1609), .Y(n_1567) );
AOI221xp5_ASAP7_75t_L g1636 ( .A1(n_1568), .A2(n_1582), .B1(n_1637), .B2(n_1638), .C(n_1644), .Y(n_1636) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1570), .Y(n_1637) );
AOI21xp5_ASAP7_75t_SL g1571 ( .A1(n_1572), .A2(n_1575), .B(n_1576), .Y(n_1571) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
NAND3xp33_ASAP7_75t_L g1577 ( .A(n_1575), .B(n_1578), .C(n_1580), .Y(n_1577) );
NAND3xp33_ASAP7_75t_SL g1576 ( .A(n_1577), .B(n_1581), .C(n_1584), .Y(n_1576) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
O2A1O1Ixp33_ASAP7_75t_L g1585 ( .A1(n_1586), .A2(n_1589), .B(n_1593), .C(n_1594), .Y(n_1585) );
INVxp67_ASAP7_75t_SL g1652 ( .A(n_1589), .Y(n_1652) );
NOR2xp33_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1592), .Y(n_1589) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1592), .Y(n_1602) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
O2A1O1Ixp33_ASAP7_75t_SL g1601 ( .A1(n_1602), .A2(n_1603), .B(n_1605), .C(n_1607), .Y(n_1601) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1613), .Y(n_1639) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
OAI221xp5_ASAP7_75t_L g1627 ( .A1(n_1628), .A2(n_1629), .B1(n_1630), .B2(n_1632), .C(n_1633), .Y(n_1627) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1640 ( .A(n_1641), .B(n_1642), .Y(n_1640) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
CKINVDCx20_ASAP7_75t_R g1653 ( .A(n_1654), .Y(n_1653) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
OAI21x1_ASAP7_75t_SL g1656 ( .A1(n_1657), .A2(n_1658), .B(n_1750), .Y(n_1656) );
NAND4xp25_ASAP7_75t_L g1750 ( .A(n_1657), .B(n_1660), .C(n_1666), .D(n_1708), .Y(n_1750) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1659), .Y(n_1658) );
NAND3xp33_ASAP7_75t_L g1659 ( .A(n_1660), .B(n_1666), .C(n_1708), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1660 ( .A(n_1661), .B(n_1662), .Y(n_1660) );
AND2x4_ASAP7_75t_L g1662 ( .A(n_1663), .B(n_1664), .Y(n_1662) );
AND2x4_ASAP7_75t_L g1747 ( .A(n_1663), .B(n_1748), .Y(n_1747) );
NOR2xp33_ASAP7_75t_L g1666 ( .A(n_1667), .B(n_1683), .Y(n_1666) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
OR2x2_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1672), .Y(n_1670) );
AOI22xp33_ASAP7_75t_L g1674 ( .A1(n_1675), .A2(n_1676), .B1(n_1680), .B2(n_1681), .Y(n_1674) );
AOI22xp33_ASAP7_75t_L g1733 ( .A1(n_1675), .A2(n_1734), .B1(n_1738), .B2(n_1741), .Y(n_1733) );
AND2x4_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1679), .Y(n_1676) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1678), .Y(n_1677) );
INVx2_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
NAND3xp33_ASAP7_75t_SL g1683 ( .A(n_1684), .B(n_1693), .C(n_1703), .Y(n_1683) );
CKINVDCx5p33_ASAP7_75t_R g1688 ( .A(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
NAND2x2_ASAP7_75t_L g1695 ( .A(n_1691), .B(n_1696), .Y(n_1695) );
INVx2_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
AOI22xp33_ASAP7_75t_SL g1693 ( .A1(n_1694), .A2(n_1698), .B1(n_1699), .B2(n_1702), .Y(n_1693) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
INVx2_ASAP7_75t_SL g1696 ( .A(n_1697), .Y(n_1696) );
INVx2_ASAP7_75t_SL g1699 ( .A(n_1700), .Y(n_1699) );
INVx1_ASAP7_75t_L g1705 ( .A(n_1706), .Y(n_1705) );
NAND3xp33_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1722), .C(n_1733), .Y(n_1709) );
NOR2xp33_ASAP7_75t_L g1710 ( .A(n_1711), .B(n_1719), .Y(n_1710) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
HB1xp67_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1715), .Y(n_1721) );
INVx4_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
CKINVDCx5p33_ASAP7_75t_R g1719 ( .A(n_1720), .Y(n_1719) );
AOI22xp33_ASAP7_75t_L g1722 ( .A1(n_1723), .A2(n_1725), .B1(n_1728), .B2(n_1731), .Y(n_1722) );
INVx3_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
BUFx2_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
HB1xp67_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx2_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx2_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1747), .Y(n_1746) );
INVx2_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1757), .Y(n_1756) );
HB1xp67_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
BUFx3_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
INVxp33_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
HB1xp67_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
NAND3xp33_ASAP7_75t_L g1763 ( .A(n_1764), .B(n_1785), .C(n_1793), .Y(n_1763) );
NOR2xp33_ASAP7_75t_L g1764 ( .A(n_1765), .B(n_1779), .Y(n_1764) );
INVx2_ASAP7_75t_SL g1802 ( .A(n_1803), .Y(n_1802) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
OAI21xp5_ASAP7_75t_L g1804 ( .A1(n_1805), .A2(n_1806), .B(n_1807), .Y(n_1804) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
endmodule