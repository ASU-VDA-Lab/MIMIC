module fake_jpeg_21926_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_4),
.B(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.C(n_1),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_10),
.C(n_11),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_6),
.C(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_26),
.Y(n_37)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_14),
.B1(n_18),
.B2(n_17),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_17),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_14),
.Y(n_38)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2x1_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_43),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_40),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_47),
.C(n_12),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_11),
.B1(n_12),
.B2(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_56),
.Y(n_60)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_46),
.C(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_37),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_43),
.B1(n_50),
.B2(n_19),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_55),
.C(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_64),
.C(n_65),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_52),
.C(n_51),
.Y(n_64)
);

FAx1_ASAP7_75t_SL g68 ( 
.A(n_66),
.B(n_35),
.CI(n_39),
.CON(n_68),
.SN(n_68)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_59),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_59),
.B(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_69),
.B1(n_35),
.B2(n_20),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_42),
.Y(n_72)
);


endmodule