module real_aes_8147_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_1), .A2(n_150), .B(n_155), .C(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g262 ( .A(n_2), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_3), .A2(n_145), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_4), .B(n_222), .Y(n_470) );
AOI21xp33_ASAP7_75t_L g223 ( .A1(n_5), .A2(n_145), .B(n_224), .Y(n_223) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_7), .A2(n_144), .B(n_152), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_8), .B(n_41), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_8), .B(n_41), .Y(n_123) );
INVx1_ASAP7_75t_L g559 ( .A(n_9), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_10), .B(n_194), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_11), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g229 ( .A(n_12), .Y(n_229) );
INVx1_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
INVx1_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_15), .A2(n_163), .B(n_177), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_16), .B(n_222), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_17), .B(n_179), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_18), .B(n_145), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_19), .B(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_20), .A2(n_210), .B(n_236), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_21), .B(n_222), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_22), .B(n_194), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g158 ( .A1(n_23), .A2(n_159), .B(n_161), .C(n_163), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_24), .B(n_194), .Y(n_456) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_25), .Y(n_487) );
INVx1_ASAP7_75t_L g455 ( .A(n_26), .Y(n_455) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_27), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_28), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_29), .B(n_194), .Y(n_263) );
INVx1_ASAP7_75t_L g480 ( .A(n_30), .Y(n_480) );
INVx1_ASAP7_75t_L g241 ( .A(n_31), .Y(n_241) );
INVx2_ASAP7_75t_L g148 ( .A(n_32), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_33), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_34), .A2(n_102), .B1(n_113), .B2(n_722), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_35), .A2(n_210), .B(n_230), .C(n_468), .Y(n_467) );
INVxp67_ASAP7_75t_L g481 ( .A(n_36), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_37), .A2(n_150), .B(n_155), .C(n_174), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_38), .A2(n_155), .B(n_454), .C(n_459), .Y(n_453) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_39), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_40), .A2(n_68), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_40), .Y(n_127) );
INVx1_ASAP7_75t_L g239 ( .A(n_42), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_43), .A2(n_181), .B(n_227), .C(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_44), .B(n_194), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g718 ( .A1(n_45), .A2(n_84), .B1(n_719), .B2(n_720), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_45), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_46), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_47), .Y(n_477) );
INVx1_ASAP7_75t_L g525 ( .A(n_48), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_49), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_50), .B(n_145), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_51), .A2(n_155), .B1(n_236), .B2(n_238), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_52), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_53), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_54), .A2(n_227), .B(n_228), .C(n_230), .Y(n_226) );
CKINVDCx14_ASAP7_75t_R g556 ( .A(n_55), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_56), .Y(n_198) );
INVx1_ASAP7_75t_L g225 ( .A(n_57), .Y(n_225) );
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_58), .A2(n_126), .B1(n_129), .B2(n_709), .C1(n_710), .C2(n_711), .Y(n_125) );
INVx1_ASAP7_75t_L g151 ( .A(n_59), .Y(n_151) );
INVx1_ASAP7_75t_L g141 ( .A(n_60), .Y(n_141) );
INVx1_ASAP7_75t_SL g469 ( .A(n_61), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_62), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_63), .B(n_222), .Y(n_529) );
INVx1_ASAP7_75t_L g490 ( .A(n_64), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_SL g249 ( .A1(n_65), .A2(n_179), .B(n_230), .C(n_250), .Y(n_249) );
INVxp67_ASAP7_75t_L g251 ( .A(n_66), .Y(n_251) );
INVx1_ASAP7_75t_L g112 ( .A(n_67), .Y(n_112) );
INVx1_ASAP7_75t_L g128 ( .A(n_68), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_69), .A2(n_145), .B(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_70), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_71), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_72), .A2(n_145), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g189 ( .A(n_73), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_74), .A2(n_144), .B(n_476), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g452 ( .A(n_75), .Y(n_452) );
INVx1_ASAP7_75t_L g517 ( .A(n_76), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_77), .A2(n_150), .B(n_155), .C(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_78), .A2(n_145), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g520 ( .A(n_79), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_80), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
INVx1_ASAP7_75t_L g509 ( .A(n_82), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_83), .B(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_84), .Y(n_719) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_85), .A2(n_150), .B(n_155), .C(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g109 ( .A(n_86), .Y(n_109) );
OR2x2_ASAP7_75t_L g120 ( .A(n_86), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g708 ( .A(n_86), .B(n_122), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_87), .A2(n_155), .B(n_489), .C(n_493), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_88), .B(n_138), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_89), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_90), .A2(n_150), .B(n_155), .C(n_207), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_91), .Y(n_215) );
INVx1_ASAP7_75t_L g248 ( .A(n_92), .Y(n_248) );
CKINVDCx16_ASAP7_75t_R g153 ( .A(n_93), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_94), .B(n_176), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_95), .B(n_167), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_96), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_97), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_98), .A2(n_145), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g528 ( .A(n_99), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_100), .Y(n_124) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx9p33_ASAP7_75t_R g723 ( .A(n_103), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_109), .C(n_110), .Y(n_107) );
AND2x2_ASAP7_75t_L g122 ( .A(n_108), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g441 ( .A(n_109), .B(n_122), .Y(n_441) );
NOR2x2_ASAP7_75t_L g713 ( .A(n_109), .B(n_121), .Y(n_713) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_125), .B1(n_714), .B2(n_716), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g715 ( .A(n_117), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_118), .A2(n_717), .B(n_721), .Y(n_716) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_124), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_120), .Y(n_721) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g709 ( .A(n_126), .Y(n_709) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_439), .B1(n_442), .B2(n_706), .Y(n_129) );
INVx2_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g710 ( .A1(n_131), .A2(n_441), .B1(n_443), .B2(n_708), .Y(n_710) );
OR4x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_335), .C(n_394), .D(n_421), .Y(n_131) );
NAND3xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_277), .C(n_302), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_200), .B(n_220), .C(n_253), .Y(n_133) );
AOI211xp5_ASAP7_75t_SL g425 ( .A1(n_134), .A2(n_426), .B(n_428), .C(n_431), .Y(n_425) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_169), .Y(n_134) );
INVx1_ASAP7_75t_L g300 ( .A(n_135), .Y(n_300) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g275 ( .A(n_136), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g307 ( .A(n_136), .Y(n_307) );
AND2x2_ASAP7_75t_L g362 ( .A(n_136), .B(n_331), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_136), .B(n_218), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_136), .B(n_219), .Y(n_420) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g281 ( .A(n_137), .Y(n_281) );
AND2x2_ASAP7_75t_L g324 ( .A(n_137), .B(n_187), .Y(n_324) );
AND2x2_ASAP7_75t_L g342 ( .A(n_137), .B(n_219), .Y(n_342) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_143), .B(n_166), .Y(n_137) );
INVx1_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
INVx2_ASAP7_75t_L g204 ( .A(n_138), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_138), .A2(n_190), .B(n_452), .C(n_453), .Y(n_451) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_138), .A2(n_554), .B(n_560), .Y(n_553) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_L g168 ( .A(n_139), .B(n_140), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_146), .B(n_150), .Y(n_190) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g458 ( .A(n_147), .Y(n_458) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
INVx1_ASAP7_75t_L g237 ( .A(n_148), .Y(n_237) );
INVx1_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
INVx3_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
INVx4_ASAP7_75t_SL g165 ( .A(n_150), .Y(n_165) );
BUFx3_ASAP7_75t_L g459 ( .A(n_150), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_158), .C(n_165), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_154), .A2(n_165), .B(n_225), .C(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_154), .A2(n_165), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_154), .A2(n_165), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g476 ( .A1(n_154), .A2(n_165), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_154), .A2(n_165), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_SL g524 ( .A1(n_154), .A2(n_165), .B(n_525), .C(n_526), .Y(n_524) );
O2A1O1Ixp33_ASAP7_75t_SL g555 ( .A1(n_154), .A2(n_165), .B(n_556), .C(n_557), .Y(n_555) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx3_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_156), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_159), .B(n_162), .Y(n_161) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_159), .A2(n_176), .B1(n_480), .B2(n_481), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_159), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_159), .B(n_528), .Y(n_527) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g238 ( .A1(n_160), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_238) );
INVx2_ASAP7_75t_L g240 ( .A(n_160), .Y(n_240) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g234 ( .A1(n_165), .A2(n_190), .B1(n_235), .B2(n_242), .Y(n_234) );
INVx1_ASAP7_75t_L g493 ( .A(n_165), .Y(n_493) );
INVx4_ASAP7_75t_L g186 ( .A(n_167), .Y(n_186) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_167), .A2(n_246), .B(n_252), .Y(n_245) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_167), .Y(n_463) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
INVx4_ASAP7_75t_L g274 ( .A(n_169), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_169), .A2(n_330), .B(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_L g410 ( .A(n_169), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_187), .Y(n_169) );
INVx1_ASAP7_75t_L g217 ( .A(n_170), .Y(n_217) );
AND2x2_ASAP7_75t_L g279 ( .A(n_170), .B(n_219), .Y(n_279) );
OR2x2_ASAP7_75t_L g308 ( .A(n_170), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g322 ( .A(n_170), .Y(n_322) );
INVx3_ASAP7_75t_L g331 ( .A(n_170), .Y(n_331) );
AND2x2_ASAP7_75t_L g341 ( .A(n_170), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g374 ( .A(n_170), .B(n_280), .Y(n_374) );
AND2x2_ASAP7_75t_L g398 ( .A(n_170), .B(n_354), .Y(n_398) );
OR2x6_ASAP7_75t_L g170 ( .A(n_171), .B(n_184), .Y(n_170) );
AOI21xp5_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B(n_182), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_178), .B(n_180), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_176), .A2(n_262), .B(n_263), .C(n_264), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_176), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
INVx5_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_177), .B(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_177), .B(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_177), .B(n_559), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_180), .A2(n_193), .B(n_195), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_180), .A2(n_490), .B(n_491), .C(n_492), .Y(n_489) );
O2A1O1Ixp5_ASAP7_75t_L g508 ( .A1(n_180), .A2(n_491), .B(n_509), .C(n_510), .Y(n_508) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g196 ( .A(n_182), .Y(n_196) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_183), .A2(n_234), .B(n_243), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_183), .B(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_183), .A2(n_258), .B(n_265), .Y(n_257) );
NOR2xp33_ASAP7_75t_SL g184 ( .A(n_185), .B(n_186), .Y(n_184) );
INVx3_ASAP7_75t_L g222 ( .A(n_186), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_186), .B(n_461), .Y(n_460) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_186), .A2(n_486), .B(n_494), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_186), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g219 ( .A(n_187), .Y(n_219) );
AND2x2_ASAP7_75t_L g434 ( .A(n_187), .B(n_276), .Y(n_434) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_196), .B(n_197), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_190), .A2(n_259), .B(n_260), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_190), .A2(n_487), .B(n_488), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_190), .A2(n_506), .B(n_507), .Y(n_505) );
INVx4_ASAP7_75t_L g210 ( .A(n_194), .Y(n_210) );
INVx2_ASAP7_75t_L g227 ( .A(n_194), .Y(n_227) );
INVx1_ASAP7_75t_L g474 ( .A(n_196), .Y(n_474) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_196), .A2(n_499), .B(n_500), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_199), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_199), .B(n_266), .Y(n_265) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_199), .A2(n_505), .B(n_511), .Y(n_504) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_216), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_202), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g354 ( .A(n_202), .B(n_342), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_202), .B(n_331), .Y(n_416) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g276 ( .A(n_203), .Y(n_276) );
AND2x2_ASAP7_75t_L g280 ( .A(n_203), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g321 ( .A(n_203), .B(n_322), .Y(n_321) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_214), .Y(n_203) );
INVx1_ASAP7_75t_L g483 ( .A(n_204), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_204), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_213), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_211), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_210), .B(n_469), .Y(n_468) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx3_ASAP7_75t_L g230 ( .A(n_212), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_216), .B(n_317), .Y(n_339) );
INVx1_ASAP7_75t_L g378 ( .A(n_216), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_216), .B(n_305), .Y(n_422) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
AND2x2_ASAP7_75t_L g285 ( .A(n_217), .B(n_280), .Y(n_285) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_219), .B(n_276), .Y(n_309) );
INVx1_ASAP7_75t_L g388 ( .A(n_219), .Y(n_388) );
AOI322xp5_ASAP7_75t_L g412 ( .A1(n_220), .A2(n_327), .A3(n_387), .B1(n_413), .B2(n_415), .C1(n_417), .C2(n_419), .Y(n_412) );
AND2x2_ASAP7_75t_SL g220 ( .A(n_221), .B(n_232), .Y(n_220) );
AND2x2_ASAP7_75t_L g267 ( .A(n_221), .B(n_245), .Y(n_267) );
INVx1_ASAP7_75t_SL g270 ( .A(n_221), .Y(n_270) );
AND2x2_ASAP7_75t_L g272 ( .A(n_221), .B(n_233), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_221), .B(n_289), .Y(n_295) );
INVx2_ASAP7_75t_L g314 ( .A(n_221), .Y(n_314) );
AND2x2_ASAP7_75t_L g327 ( .A(n_221), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g365 ( .A(n_221), .B(n_289), .Y(n_365) );
BUFx2_ASAP7_75t_L g382 ( .A(n_221), .Y(n_382) );
AND2x2_ASAP7_75t_L g396 ( .A(n_221), .B(n_256), .Y(n_396) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_231), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_232), .B(n_284), .Y(n_311) );
AND2x2_ASAP7_75t_L g438 ( .A(n_232), .B(n_314), .Y(n_438) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_245), .Y(n_232) );
OR2x2_ASAP7_75t_L g283 ( .A(n_233), .B(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g289 ( .A(n_233), .Y(n_289) );
AND2x2_ASAP7_75t_L g334 ( .A(n_233), .B(n_257), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_233), .B(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_233), .Y(n_418) );
INVx2_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g491 ( .A(n_240), .Y(n_491) );
AND2x2_ASAP7_75t_L g269 ( .A(n_245), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g291 ( .A(n_245), .Y(n_291) );
BUFx2_ASAP7_75t_L g297 ( .A(n_245), .Y(n_297) );
AND2x2_ASAP7_75t_L g316 ( .A(n_245), .B(n_289), .Y(n_316) );
INVx3_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
OR2x2_ASAP7_75t_L g338 ( .A(n_245), .B(n_289), .Y(n_338) );
AOI31xp33_ASAP7_75t_SL g253 ( .A1(n_254), .A2(n_268), .A3(n_271), .B(n_273), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_267), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_255), .B(n_290), .Y(n_301) );
OR2x2_ASAP7_75t_L g325 ( .A(n_255), .B(n_295), .Y(n_325) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_256), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g346 ( .A(n_256), .B(n_338), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_256), .B(n_328), .Y(n_356) );
AND2x2_ASAP7_75t_L g363 ( .A(n_256), .B(n_364), .Y(n_363) );
NAND2x1_ASAP7_75t_L g391 ( .A(n_256), .B(n_327), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_256), .B(n_382), .Y(n_392) );
AND2x2_ASAP7_75t_L g404 ( .A(n_256), .B(n_289), .Y(n_404) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx3_ASAP7_75t_L g284 ( .A(n_257), .Y(n_284) );
INVx1_ASAP7_75t_L g350 ( .A(n_267), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_267), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_269), .B(n_345), .Y(n_379) );
AND2x4_ASAP7_75t_L g290 ( .A(n_270), .B(n_291), .Y(n_290) );
CKINVDCx16_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g369 ( .A(n_275), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_275), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g317 ( .A(n_276), .B(n_307), .Y(n_317) );
AND2x2_ASAP7_75t_L g411 ( .A(n_276), .B(n_281), .Y(n_411) );
INVx1_ASAP7_75t_L g436 ( .A(n_276), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_282), .B1(n_285), .B2(n_286), .C(n_292), .Y(n_277) );
CKINVDCx14_ASAP7_75t_R g298 ( .A(n_278), .Y(n_298) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_279), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_282), .B(n_333), .Y(n_352) );
INVx3_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g401 ( .A(n_283), .B(n_297), .Y(n_401) );
AND2x2_ASAP7_75t_L g315 ( .A(n_284), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g345 ( .A(n_284), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_284), .B(n_328), .Y(n_373) );
NOR3xp33_ASAP7_75t_L g415 ( .A(n_284), .B(n_385), .C(n_416), .Y(n_415) );
AOI211xp5_ASAP7_75t_SL g348 ( .A1(n_285), .A2(n_349), .B(n_351), .C(n_359), .Y(n_348) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_287), .A2(n_338), .B1(n_339), .B2(n_340), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_288), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_288), .B(n_372), .Y(n_371) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g430 ( .A(n_290), .B(n_404), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_298), .B1(n_299), .B2(n_301), .Y(n_292) );
NOR2xp33_ASAP7_75t_SL g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_296), .B(n_345), .Y(n_376) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_299), .A2(n_391), .B1(n_422), .B2(n_429), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_310), .B1(n_312), .B2(n_317), .C(n_318), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_308), .A2(n_319), .B1(n_325), .B2(n_326), .C(n_329), .Y(n_318) );
INVx1_ASAP7_75t_L g361 ( .A(n_309), .Y(n_361) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_SL g333 ( .A(n_314), .Y(n_333) );
OR2x2_ASAP7_75t_L g406 ( .A(n_314), .B(n_338), .Y(n_406) );
AND2x2_ASAP7_75t_L g408 ( .A(n_314), .B(n_316), .Y(n_408) );
INVx1_ASAP7_75t_L g347 ( .A(n_317), .Y(n_347) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
AOI21xp33_ASAP7_75t_SL g377 ( .A1(n_320), .A2(n_378), .B(n_379), .Y(n_377) );
OR2x2_ASAP7_75t_L g384 ( .A(n_320), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g358 ( .A(n_321), .B(n_342), .Y(n_358) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp33_ASAP7_75t_SL g375 ( .A(n_326), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_327), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_328), .B(n_364), .Y(n_427) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_331), .A2(n_344), .B(n_346), .C(n_347), .Y(n_343) );
NAND2x1_ASAP7_75t_SL g368 ( .A(n_331), .B(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_332), .A2(n_381), .B1(n_383), .B2(n_386), .Y(n_380) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_334), .B(n_424), .Y(n_423) );
NAND5xp2_ASAP7_75t_L g335 ( .A(n_336), .B(n_348), .C(n_366), .D(n_380), .E(n_389), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_343), .Y(n_336) );
INVx1_ASAP7_75t_L g393 ( .A(n_339), .Y(n_393) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_341), .A2(n_360), .B1(n_400), .B2(n_402), .C(n_405), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_342), .B(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_345), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_345), .B(n_411), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_355), .B2(n_357), .Y(n_351) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_L g433 ( .A(n_362), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B1(n_374), .B2(n_375), .C(n_377), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g417 ( .A(n_372), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g424 ( .A(n_382), .Y(n_424) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_392), .B(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI211xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_397), .B(n_399), .C(n_412), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
A2O1A1Ixp33_ASAP7_75t_L g421 ( .A1(n_397), .A2(n_422), .B(n_423), .C(n_425), .Y(n_421) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_401), .B(n_403), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B(n_409), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B(n_437), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
XOR2xp5_ASAP7_75t_L g717 ( .A(n_443), .B(n_718), .Y(n_717) );
OR3x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_617), .C(n_664), .Y(n_443) );
NAND3xp33_ASAP7_75t_SL g444 ( .A(n_445), .B(n_563), .C(n_588), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_503), .B1(n_530), .B2(n_533), .C(n_541), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_471), .B(n_496), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_448), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_448), .B(n_546), .Y(n_661) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_462), .Y(n_448) );
AND2x2_ASAP7_75t_L g532 ( .A(n_449), .B(n_502), .Y(n_532) );
AND2x2_ASAP7_75t_L g581 ( .A(n_449), .B(n_501), .Y(n_581) );
AND2x2_ASAP7_75t_L g602 ( .A(n_449), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g607 ( .A(n_449), .B(n_574), .Y(n_607) );
OR2x2_ASAP7_75t_L g615 ( .A(n_449), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g687 ( .A(n_449), .B(n_484), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_449), .B(n_636), .Y(n_701) );
INVx3_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g547 ( .A(n_450), .B(n_462), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_450), .B(n_484), .Y(n_548) );
AND2x4_ASAP7_75t_L g569 ( .A(n_450), .B(n_502), .Y(n_569) );
AND2x2_ASAP7_75t_L g599 ( .A(n_450), .B(n_473), .Y(n_599) );
AND2x2_ASAP7_75t_L g608 ( .A(n_450), .B(n_598), .Y(n_608) );
AND2x2_ASAP7_75t_L g624 ( .A(n_450), .B(n_485), .Y(n_624) );
OR2x2_ASAP7_75t_L g633 ( .A(n_450), .B(n_616), .Y(n_633) );
AND2x2_ASAP7_75t_L g639 ( .A(n_450), .B(n_574), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_450), .B(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g653 ( .A(n_450), .B(n_498), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_450), .B(n_543), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_450), .B(n_603), .Y(n_692) );
OR2x6_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_458), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g502 ( .A(n_462), .Y(n_502) );
AND2x2_ASAP7_75t_L g598 ( .A(n_462), .B(n_484), .Y(n_598) );
AND2x2_ASAP7_75t_L g603 ( .A(n_462), .B(n_485), .Y(n_603) );
INVx1_ASAP7_75t_L g659 ( .A(n_462), .Y(n_659) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B(n_470), .Y(n_462) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_463), .A2(n_515), .B(n_521), .Y(n_514) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_463), .A2(n_523), .B(n_529), .Y(n_522) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g568 ( .A(n_472), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_484), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_473), .B(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g546 ( .A(n_473), .Y(n_546) );
OR2x2_ASAP7_75t_L g616 ( .A(n_473), .B(n_484), .Y(n_616) );
OR2x2_ASAP7_75t_L g677 ( .A(n_473), .B(n_584), .Y(n_677) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_482), .Y(n_473) );
INVx1_ASAP7_75t_L g499 ( .A(n_475), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_482), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_484), .B(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g636 ( .A(n_484), .B(n_498), .Y(n_636) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g575 ( .A(n_485), .Y(n_575) );
INVx1_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_497), .A2(n_681), .B1(n_685), .B2(n_688), .C(n_689), .Y(n_680) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .Y(n_497) );
INVx1_ASAP7_75t_SL g544 ( .A(n_498), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_498), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g675 ( .A(n_498), .B(n_532), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_501), .B(n_546), .Y(n_667) );
AND2x2_ASAP7_75t_L g574 ( .A(n_502), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g578 ( .A(n_503), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_503), .B(n_584), .Y(n_614) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
AND2x2_ASAP7_75t_L g540 ( .A(n_504), .B(n_514), .Y(n_540) );
INVx4_ASAP7_75t_L g552 ( .A(n_504), .Y(n_552) );
BUFx3_ASAP7_75t_L g594 ( .A(n_504), .Y(n_594) );
AND3x2_ASAP7_75t_L g609 ( .A(n_504), .B(n_610), .C(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g691 ( .A(n_513), .B(n_605), .Y(n_691) );
AND2x2_ASAP7_75t_L g699 ( .A(n_513), .B(n_584), .Y(n_699) );
INVx1_ASAP7_75t_SL g704 ( .A(n_513), .Y(n_704) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_522), .Y(n_513) );
INVx1_ASAP7_75t_SL g562 ( .A(n_514), .Y(n_562) );
AND2x2_ASAP7_75t_L g585 ( .A(n_514), .B(n_552), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_514), .B(n_536), .Y(n_587) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_514), .Y(n_627) );
OR2x2_ASAP7_75t_L g632 ( .A(n_514), .B(n_552), .Y(n_632) );
INVx2_ASAP7_75t_L g538 ( .A(n_522), .Y(n_538) );
AND2x2_ASAP7_75t_L g572 ( .A(n_522), .B(n_553), .Y(n_572) );
OR2x2_ASAP7_75t_L g592 ( .A(n_522), .B(n_553), .Y(n_592) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_522), .Y(n_612) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_531), .A2(n_571), .B(n_663), .Y(n_662) );
AOI322xp5_ASAP7_75t_L g698 ( .A1(n_533), .A2(n_543), .A3(n_569), .B1(n_699), .B2(n_700), .C1(n_702), .C2(n_705), .Y(n_698) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_535), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_536), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g561 ( .A(n_537), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g629 ( .A(n_538), .B(n_552), .Y(n_629) );
AND2x2_ASAP7_75t_L g696 ( .A(n_538), .B(n_553), .Y(n_696) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g637 ( .A(n_540), .B(n_591), .Y(n_637) );
AOI31xp33_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_545), .A3(n_548), .B(n_549), .Y(n_541) );
AND2x2_ASAP7_75t_L g596 ( .A(n_543), .B(n_574), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_543), .B(n_566), .Y(n_678) );
AND2x2_ASAP7_75t_L g697 ( .A(n_543), .B(n_602), .Y(n_697) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_546), .B(n_574), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_546), .B(n_603), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_546), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_546), .B(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_547), .B(n_603), .Y(n_635) );
INVx1_ASAP7_75t_L g679 ( .A(n_547), .Y(n_679) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_561), .Y(n_550) );
INVxp67_ASAP7_75t_L g631 ( .A(n_551), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_552), .B(n_562), .Y(n_567) );
INVx1_ASAP7_75t_L g673 ( .A(n_552), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_552), .B(n_650), .Y(n_684) );
BUFx3_ASAP7_75t_L g584 ( .A(n_553), .Y(n_584) );
AND2x2_ASAP7_75t_L g610 ( .A(n_553), .B(n_562), .Y(n_610) );
INVx2_ASAP7_75t_L g650 ( .A(n_553), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_561), .B(n_683), .Y(n_682) );
AOI211xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_568), .B(n_570), .C(n_579), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI21xp33_ASAP7_75t_L g613 ( .A1(n_565), .A2(n_614), .B(n_615), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_566), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_566), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g646 ( .A(n_567), .B(n_592), .Y(n_646) );
INVx3_ASAP7_75t_L g577 ( .A(n_569), .Y(n_577) );
OAI22xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_573), .B1(n_576), .B2(n_578), .Y(n_570) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_572), .A2(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g621 ( .A(n_572), .B(n_585), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_572), .B(n_673), .Y(n_672) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g576 ( .A(n_575), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g645 ( .A(n_575), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g589 ( .A1(n_576), .A2(n_590), .B(n_595), .Y(n_589) );
OAI22xp33_ASAP7_75t_SL g579 ( .A1(n_580), .A2(n_582), .B1(n_586), .B2(n_587), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_581), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g605 ( .A(n_584), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_584), .B(n_627), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_600), .C(n_613), .Y(n_588) );
OAI22xp5_ASAP7_75t_SL g655 ( .A1(n_590), .A2(n_656), .B1(n_660), .B2(n_661), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g660 ( .A(n_592), .B(n_593), .Y(n_660) );
AND2x2_ASAP7_75t_L g668 ( .A(n_593), .B(n_649), .Y(n_668) );
CKINVDCx16_ASAP7_75t_R g593 ( .A(n_594), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_SL g676 ( .A1(n_594), .A2(n_677), .B(n_678), .C(n_679), .Y(n_676) );
OR2x2_ASAP7_75t_L g703 ( .A(n_594), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_604), .B(n_606), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_602), .A2(n_639), .B(n_640), .C(n_643), .Y(n_638) );
OAI21xp33_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_608), .B(n_609), .Y(n_606) );
AND2x2_ASAP7_75t_L g671 ( .A(n_610), .B(n_629), .Y(n_671) );
INVxp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g649 ( .A(n_612), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g654 ( .A(n_614), .Y(n_654) );
NAND3xp33_ASAP7_75t_SL g617 ( .A(n_618), .B(n_638), .C(n_651), .Y(n_617) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_621), .B(n_622), .C(n_630), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g688 ( .A(n_625), .Y(n_688) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g648 ( .A(n_627), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_627), .B(n_696), .Y(n_695) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B(n_633), .C(n_634), .Y(n_630) );
INVx2_ASAP7_75t_SL g642 ( .A(n_632), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_633), .A2(n_644), .B1(n_646), .B2(n_647), .Y(n_643) );
OAI21xp33_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_636), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_655), .C(n_662), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
INVxp33_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g705 ( .A(n_659), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_680), .C(n_693), .D(n_698), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B(n_669), .C(n_676), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B(n_674), .Y(n_669) );
AOI21xp33_ASAP7_75t_L g689 ( .A1(n_670), .A2(n_690), .B(n_692), .Y(n_689) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_677), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
endmodule