module real_aes_10347_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_571;
wire n_549;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_360;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_1102;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1584;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g561 ( .A(n_0), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_0), .A2(n_171), .B1(n_293), .B2(n_332), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_1), .A2(n_243), .B1(n_483), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_1), .A2(n_243), .B1(n_319), .B2(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g757 ( .A(n_2), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_2), .A2(n_148), .B1(n_416), .B2(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g1010 ( .A(n_3), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_4), .A2(n_14), .B1(n_568), .B2(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g786 ( .A(n_4), .Y(n_786) );
INVx1_ASAP7_75t_L g867 ( .A(n_5), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_6), .A2(n_181), .B1(n_533), .B2(n_537), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_6), .A2(n_181), .B1(n_899), .B2(n_948), .Y(n_951) );
INVxp33_ASAP7_75t_L g1003 ( .A(n_7), .Y(n_1003) );
AOI21xp5_ASAP7_75t_L g1041 ( .A1(n_7), .A2(n_1042), .B(n_1043), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g1162 ( .A(n_8), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_8), .A2(n_51), .B1(n_1178), .B2(n_1181), .Y(n_1177) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_9), .Y(n_347) );
INVx1_ASAP7_75t_L g437 ( .A(n_9), .Y(n_437) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_9), .B(n_296), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_9), .B(n_206), .Y(n_1031) );
AOI22xp5_ASAP7_75t_L g1253 ( .A1(n_10), .A2(n_11), .B1(n_1229), .B2(n_1242), .Y(n_1253) );
INVx1_ASAP7_75t_L g1007 ( .A(n_12), .Y(n_1007) );
OAI21xp33_ASAP7_75t_SL g690 ( .A1(n_13), .A2(n_548), .B(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_13), .A2(n_128), .B1(n_726), .B2(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g787 ( .A(n_14), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g1235 ( .A1(n_15), .A2(n_247), .B1(n_1236), .B2(n_1239), .Y(n_1235) );
INVx1_ASAP7_75t_L g1012 ( .A(n_16), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g1024 ( .A1(n_16), .A2(n_278), .B1(n_1025), .B2(n_1032), .C(n_1034), .Y(n_1024) );
AOI221xp5_ASAP7_75t_SL g1094 ( .A1(n_17), .A2(n_42), .B1(n_1095), .B2(n_1096), .C(n_1097), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_17), .A2(n_42), .B1(n_948), .B2(n_1116), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_18), .A2(n_215), .B1(n_416), .B2(n_667), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_18), .A2(n_215), .B1(n_945), .B2(n_946), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_19), .A2(n_271), .B1(n_463), .B2(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_19), .A2(n_271), .B1(n_533), .B2(n_537), .Y(n_532) );
INVx1_ASAP7_75t_L g695 ( .A(n_20), .Y(n_695) );
OAI222xp33_ASAP7_75t_L g703 ( .A1(n_20), .A2(n_33), .B1(n_269), .B2(n_325), .C1(n_500), .C2(n_673), .Y(n_703) );
AO22x2_ASAP7_75t_L g854 ( .A1(n_21), .A2(n_855), .B1(n_908), .B2(n_909), .Y(n_854) );
INVx1_ASAP7_75t_L g908 ( .A(n_21), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_22), .A2(n_139), .B1(n_824), .B2(n_825), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_22), .A2(n_139), .B1(n_841), .B2(n_843), .Y(n_840) );
CKINVDCx14_ASAP7_75t_R g1245 ( .A(n_23), .Y(n_1245) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_24), .Y(n_751) );
INVx1_ASAP7_75t_L g1481 ( .A(n_25), .Y(n_1481) );
INVx1_ASAP7_75t_L g1136 ( .A(n_26), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g887 ( .A1(n_27), .A2(n_270), .B1(n_413), .B2(n_888), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_27), .A2(n_270), .B1(n_380), .B2(n_742), .Y(n_895) );
INVx1_ASAP7_75t_L g755 ( .A(n_28), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_28), .A2(n_277), .B1(n_767), .B2(n_768), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_29), .A2(n_209), .B1(n_474), .B2(n_489), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1102 ( .A1(n_29), .A2(n_209), .B1(n_404), .B2(n_1103), .C(n_1106), .Y(n_1102) );
INVxp67_ASAP7_75t_SL g818 ( .A(n_30), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_30), .A2(n_212), .B1(n_774), .B2(n_849), .Y(n_848) );
INVxp33_ASAP7_75t_L g333 ( .A(n_31), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_31), .A2(n_238), .B1(n_440), .B2(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g354 ( .A(n_32), .Y(n_354) );
OR2x2_ASAP7_75t_L g1498 ( .A(n_32), .B(n_1492), .Y(n_1498) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_33), .A2(n_179), .B1(n_735), .B2(n_742), .Y(n_741) );
INVxp67_ASAP7_75t_SL g1018 ( .A(n_34), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_34), .A2(n_265), .B1(n_836), .B2(n_849), .Y(n_1070) );
AOI22xp33_ASAP7_75t_SL g1566 ( .A1(n_35), .A2(n_83), .B1(n_723), .B2(n_833), .Y(n_1566) );
AOI22xp33_ASAP7_75t_L g1577 ( .A1(n_35), .A2(n_83), .B1(n_740), .B2(n_744), .Y(n_1577) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_36), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_37), .A2(n_240), .B1(n_650), .B2(n_961), .Y(n_960) );
INVxp67_ASAP7_75t_SL g988 ( .A(n_37), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_38), .A2(n_201), .B1(n_442), .B2(n_971), .Y(n_970) );
OAI211xp5_ASAP7_75t_SL g974 ( .A1(n_38), .A2(n_339), .B(n_975), .C(n_978), .Y(n_974) );
BUFx2_ASAP7_75t_L g344 ( .A(n_39), .Y(n_344) );
BUFx2_ASAP7_75t_L g400 ( .A(n_39), .Y(n_400) );
INVx1_ASAP7_75t_L g435 ( .A(n_39), .Y(n_435) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_39), .B(n_1031), .Y(n_1454) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_40), .A2(n_53), .B1(n_566), .B2(n_569), .Y(n_565) );
OAI211xp5_ASAP7_75t_L g608 ( .A1(n_40), .A2(n_339), .B(n_609), .C(n_612), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_41), .A2(n_111), .B1(n_463), .B2(n_662), .Y(n_661) );
INVxp67_ASAP7_75t_L g676 ( .A(n_41), .Y(n_676) );
INVx1_ASAP7_75t_L g697 ( .A(n_43), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_43), .A2(n_179), .B1(n_293), .B2(n_332), .Y(n_702) );
INVxp33_ASAP7_75t_L g1005 ( .A(n_44), .Y(n_1005) );
AOI221xp5_ASAP7_75t_L g1039 ( .A1(n_44), .A2(n_99), .B1(n_726), .B2(n_937), .C(n_1040), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_45), .A2(n_184), .B1(n_416), .B2(n_652), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_45), .A2(n_184), .B1(n_483), .B2(n_660), .Y(n_964) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_46), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_46), .A2(n_127), .B1(n_325), .B2(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g1482 ( .A(n_47), .Y(n_1482) );
INVxp33_ASAP7_75t_SL g1546 ( .A(n_48), .Y(n_1546) );
AOI22xp33_ASAP7_75t_SL g1581 ( .A1(n_48), .A2(n_55), .B1(n_1582), .B2(n_1583), .Y(n_1581) );
INVx1_ASAP7_75t_L g1563 ( .A(n_49), .Y(n_1563) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_49), .A2(n_180), .B1(n_318), .B2(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g378 ( .A(n_50), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_50), .A2(n_150), .B1(n_412), .B2(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_SL g1165 ( .A(n_51), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_52), .A2(n_259), .B1(n_416), .B2(n_652), .Y(n_1166) );
AOI221xp5_ASAP7_75t_SL g1173 ( .A1(n_52), .A2(n_451), .B1(n_559), .B2(n_1174), .C(n_1175), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_53), .A2(n_109), .B1(n_533), .B2(n_537), .Y(n_615) );
OAI211xp5_ASAP7_75t_L g1132 ( .A1(n_54), .A2(n_484), .B(n_1133), .C(n_1135), .Y(n_1132) );
INVx1_ASAP7_75t_L g1156 ( .A(n_54), .Y(n_1156) );
INVxp33_ASAP7_75t_SL g1547 ( .A(n_55), .Y(n_1547) );
INVx1_ASAP7_75t_L g861 ( .A(n_56), .Y(n_861) );
XNOR2xp5_ASAP7_75t_L g912 ( .A(n_57), .B(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_58), .A2(n_152), .B1(n_412), .B2(n_416), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_58), .A2(n_152), .B1(n_440), .B2(n_442), .Y(n_439) );
INVxp33_ASAP7_75t_SL g1554 ( .A(n_59), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g1580 ( .A1(n_59), .A2(n_62), .B1(n_758), .B2(n_841), .Y(n_1580) );
INVx1_ASAP7_75t_L g1083 ( .A(n_60), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_60), .A2(n_197), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
CKINVDCx5p33_ASAP7_75t_R g1099 ( .A(n_61), .Y(n_1099) );
INVx1_ASAP7_75t_L g1549 ( .A(n_62), .Y(n_1549) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_63), .A2(n_245), .B1(n_442), .B2(n_660), .Y(n_659) );
INVxp33_ASAP7_75t_L g678 ( .A(n_63), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_64), .A2(n_232), .B1(n_416), .B2(n_667), .Y(n_962) );
INVx1_ASAP7_75t_L g985 ( .A(n_64), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_65), .A2(n_86), .B1(n_474), .B2(n_479), .Y(n_473) );
INVx1_ASAP7_75t_L g506 ( .A(n_65), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g1241 ( .A1(n_66), .A2(n_96), .B1(n_1229), .B2(n_1242), .Y(n_1241) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_67), .A2(n_257), .B1(n_489), .B2(n_490), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_67), .A2(n_257), .B1(n_404), .B2(n_426), .C(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g1445 ( .A(n_68), .Y(n_1445) );
INVxp33_ASAP7_75t_SL g1559 ( .A(n_69), .Y(n_1559) );
AOI22xp33_ASAP7_75t_L g1569 ( .A1(n_69), .A2(n_149), .B1(n_723), .B2(n_1570), .Y(n_1569) );
OAI221xp5_ASAP7_75t_L g1449 ( .A1(n_70), .A2(n_224), .B1(n_1450), .B2(n_1455), .C(n_1458), .Y(n_1449) );
OAI22xp5_ASAP7_75t_L g1499 ( .A1(n_70), .A2(n_224), .B1(n_1500), .B2(n_1503), .Y(n_1499) );
INVx1_ASAP7_75t_L g604 ( .A(n_71), .Y(n_604) );
OAI211xp5_ASAP7_75t_SL g619 ( .A1(n_71), .A2(n_390), .B(n_620), .C(n_622), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_72), .A2(n_218), .B1(n_710), .B2(n_713), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_72), .A2(n_235), .B1(n_733), .B2(n_735), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_73), .A2(n_263), .B1(n_483), .B2(n_647), .Y(n_777) );
INVx1_ASAP7_75t_L g783 ( .A(n_73), .Y(n_783) );
INVxp67_ASAP7_75t_L g1472 ( .A(n_74), .Y(n_1472) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_74), .A2(n_125), .B1(n_440), .B2(n_662), .Y(n_1517) );
AOI22xp5_ASAP7_75t_SL g1249 ( .A1(n_75), .A2(n_84), .B1(n_1223), .B2(n_1229), .Y(n_1249) );
INVx1_ASAP7_75t_L g921 ( .A(n_76), .Y(n_921) );
INVx1_ASAP7_75t_L g924 ( .A(n_77), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_77), .A2(n_133), .B1(n_726), .B2(n_767), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_78), .A2(n_249), .B1(n_404), .B2(n_407), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_78), .A2(n_249), .B1(n_445), .B2(n_448), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g1227 ( .A(n_79), .Y(n_1227) );
INVx1_ASAP7_75t_L g323 ( .A(n_80), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_81), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g1079 ( .A(n_82), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_85), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_85), .A2(n_210), .B1(n_494), .B2(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g531 ( .A(n_86), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_87), .A2(n_197), .B1(n_533), .B2(n_537), .Y(n_1076) );
INVx1_ASAP7_75t_L g1120 ( .A(n_87), .Y(n_1120) );
INVx1_ASAP7_75t_L g634 ( .A(n_88), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_88), .A2(n_95), .B1(n_672), .B2(n_673), .Y(n_671) );
INVx1_ASAP7_75t_L g991 ( .A(n_89), .Y(n_991) );
INVx1_ASAP7_75t_L g398 ( .A(n_90), .Y(n_398) );
INVx1_ASAP7_75t_L g1492 ( .A(n_90), .Y(n_1492) );
INVxp33_ASAP7_75t_SL g873 ( .A(n_91), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_91), .A2(n_202), .B1(n_555), .B2(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g864 ( .A(n_92), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_92), .A2(n_192), .B1(n_710), .B2(n_888), .Y(n_893) );
INVx1_ASAP7_75t_L g980 ( .A(n_93), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_94), .A2(n_205), .B1(n_494), .B2(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_94), .A2(n_205), .B1(n_897), .B2(n_900), .Y(n_896) );
INVx1_ASAP7_75t_L g636 ( .A(n_95), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g1567 ( .A1(n_97), .A2(n_106), .B1(n_318), .B2(n_413), .Y(n_1567) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_97), .A2(n_106), .B1(n_845), .B2(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g497 ( .A(n_98), .Y(n_497) );
INVxp67_ASAP7_75t_SL g1008 ( .A(n_99), .Y(n_1008) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_100), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_100), .A2(n_262), .B1(n_832), .B2(n_833), .Y(n_831) );
INVx1_ASAP7_75t_L g760 ( .A(n_101), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g784 ( .A1(n_101), .A2(n_191), .B1(n_325), .B2(n_673), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_102), .A2(n_154), .B1(n_563), .B2(n_568), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_102), .A2(n_154), .B1(n_533), .B2(n_537), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_103), .A2(n_118), .B1(n_303), .B2(n_584), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_103), .A2(n_118), .B1(n_836), .B2(n_1061), .Y(n_1060) );
INVxp67_ASAP7_75t_L g1464 ( .A(n_104), .Y(n_1464) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_104), .A2(n_122), .B1(n_1514), .B2(n_1515), .C(n_1516), .Y(n_1513) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_105), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_107), .A2(n_252), .B1(n_1236), .B2(n_1293), .Y(n_1292) );
CKINVDCx20_ASAP7_75t_R g1333 ( .A(n_108), .Y(n_1333) );
INVx1_ASAP7_75t_L g564 ( .A(n_109), .Y(n_564) );
INVx1_ASAP7_75t_L g1550 ( .A(n_110), .Y(n_1550) );
INVxp33_ASAP7_75t_L g675 ( .A(n_111), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_112), .A2(n_135), .B1(n_474), .B2(n_489), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g722 ( .A1(n_112), .A2(n_135), .B1(n_413), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_113), .A2(n_242), .B1(n_428), .B2(n_650), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_113), .A2(n_242), .B1(n_563), .B2(n_774), .Y(n_773) );
OAI211xp5_ASAP7_75t_L g1141 ( .A1(n_114), .A2(n_339), .B(n_1142), .C(n_1143), .Y(n_1141) );
INVx1_ASAP7_75t_L g1169 ( .A(n_114), .Y(n_1169) );
INVxp33_ASAP7_75t_L g1438 ( .A(n_115), .Y(n_1438) );
AOI221xp5_ASAP7_75t_L g1505 ( .A1(n_115), .A2(n_155), .B1(n_897), .B2(n_948), .C(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g596 ( .A(n_116), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_116), .A2(n_141), .B1(n_474), .B2(n_489), .Y(n_617) );
AO22x2_ASAP7_75t_L g624 ( .A1(n_117), .A2(n_625), .B1(n_681), .B2(n_682), .Y(n_624) );
INVx1_ASAP7_75t_L g681 ( .A(n_117), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g541 ( .A(n_119), .B(n_542), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_120), .A2(n_186), .B1(n_474), .B2(n_489), .Y(n_1138) );
INVx1_ASAP7_75t_L g1148 ( .A(n_120), .Y(n_1148) );
INVx1_ASAP7_75t_L g1192 ( .A(n_121), .Y(n_1192) );
INVxp67_ASAP7_75t_L g1469 ( .A(n_122), .Y(n_1469) );
AOI221xp5_ASAP7_75t_L g493 ( .A1(n_123), .A2(n_217), .B1(n_494), .B2(n_495), .C(n_496), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_123), .A2(n_217), .B1(n_463), .B2(n_464), .Y(n_519) );
INVx1_ASAP7_75t_L g487 ( .A(n_124), .Y(n_487) );
INVx1_ASAP7_75t_L g1463 ( .A(n_125), .Y(n_1463) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_126), .A2(n_201), .B1(n_293), .B2(n_332), .Y(n_981) );
OAI22xp33_ASAP7_75t_L g990 ( .A1(n_126), .A2(n_232), .B1(n_474), .B2(n_479), .Y(n_990) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_127), .Y(n_801) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_128), .Y(n_698) );
INVx1_ASAP7_75t_L g1442 ( .A(n_129), .Y(n_1442) );
AOI22xp5_ASAP7_75t_L g1248 ( .A1(n_130), .A2(n_234), .B1(n_1236), .B2(n_1239), .Y(n_1248) );
INVx1_ASAP7_75t_L g638 ( .A(n_131), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_132), .A2(n_172), .B1(n_553), .B2(n_555), .Y(n_552) );
INVx1_ASAP7_75t_L g577 ( .A(n_132), .Y(n_577) );
INVxp67_ASAP7_75t_SL g923 ( .A(n_133), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_134), .A2(n_164), .B1(n_716), .B2(n_828), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_134), .A2(n_164), .B1(n_836), .B2(n_838), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g1294 ( .A1(n_136), .A2(n_137), .B1(n_1223), .B2(n_1295), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_138), .A2(n_145), .B1(n_447), .B2(n_464), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_138), .A2(n_145), .B1(n_428), .B2(n_650), .Y(n_665) );
INVx1_ASAP7_75t_L g288 ( .A(n_140), .Y(n_288) );
INVx1_ASAP7_75t_L g592 ( .A(n_141), .Y(n_592) );
CKINVDCx14_ASAP7_75t_R g470 ( .A(n_142), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g1252 ( .A1(n_143), .A2(n_167), .B1(n_1236), .B2(n_1239), .Y(n_1252) );
INVx1_ASAP7_75t_L g486 ( .A(n_144), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_146), .A2(n_235), .B1(n_716), .B2(n_718), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_146), .A2(n_218), .B1(n_738), .B2(n_740), .Y(n_737) );
INVxp33_ASAP7_75t_SL g628 ( .A(n_147), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_147), .A2(n_160), .B1(n_319), .B2(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g754 ( .A(n_148), .Y(n_754) );
INVxp67_ASAP7_75t_SL g1561 ( .A(n_149), .Y(n_1561) );
INVxp33_ASAP7_75t_L g350 ( .A(n_150), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_151), .A2(n_157), .B1(n_650), .B2(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_151), .A2(n_157), .B1(n_899), .B2(n_966), .Y(n_965) );
OAI22xp33_ASAP7_75t_L g925 ( .A1(n_153), .A2(n_194), .B1(n_474), .B2(n_479), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_153), .A2(n_231), .B1(n_770), .B2(n_942), .Y(n_941) );
INVxp33_ASAP7_75t_L g1447 ( .A(n_155), .Y(n_1447) );
INVx1_ASAP7_75t_L g1551 ( .A(n_156), .Y(n_1551) );
CKINVDCx5p33_ASAP7_75t_R g1080 ( .A(n_158), .Y(n_1080) );
INVxp67_ASAP7_75t_SL g362 ( .A(n_159), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_159), .A2(n_211), .B1(n_425), .B2(n_426), .Y(n_424) );
INVxp67_ASAP7_75t_SL g631 ( .A(n_160), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g1098 ( .A(n_161), .Y(n_1098) );
INVxp33_ASAP7_75t_SL g639 ( .A(n_162), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_162), .A2(n_182), .B1(n_428), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_163), .A2(n_254), .B1(n_319), .B2(n_667), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_163), .A2(n_254), .B1(n_483), .B2(n_647), .Y(n_772) );
AO221x2_ASAP7_75t_L g1243 ( .A1(n_165), .A2(n_261), .B1(n_1229), .B2(n_1242), .C(n_1244), .Y(n_1243) );
CKINVDCx16_ASAP7_75t_R g1230 ( .A(n_166), .Y(n_1230) );
INVx1_ASAP7_75t_L g301 ( .A(n_168), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g1131 ( .A1(n_169), .A2(n_233), .B1(n_479), .B2(n_490), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g1144 ( .A1(n_169), .A2(n_204), .B1(n_293), .B2(n_332), .Y(n_1144) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_170), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_170), .B(n_1192), .Y(n_1210) );
AND3x2_ASAP7_75t_L g1226 ( .A(n_170), .B(n_1192), .C(n_1213), .Y(n_1226) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_171), .A2(n_239), .B1(n_479), .B2(n_490), .Y(n_618) );
INVx1_ASAP7_75t_L g585 ( .A(n_172), .Y(n_585) );
INVxp33_ASAP7_75t_SL g806 ( .A(n_173), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_173), .A2(n_250), .B1(n_318), .B2(n_824), .Y(n_830) );
INVx1_ASAP7_75t_L g920 ( .A(n_174), .Y(n_920) );
AOI22xp5_ASAP7_75t_SL g1261 ( .A1(n_175), .A2(n_188), .B1(n_1223), .B2(n_1229), .Y(n_1261) );
INVx2_ASAP7_75t_L g300 ( .A(n_176), .Y(n_300) );
AOI22xp5_ASAP7_75t_SL g1260 ( .A1(n_177), .A2(n_256), .B1(n_1236), .B2(n_1239), .Y(n_1260) );
INVx1_ASAP7_75t_L g1477 ( .A(n_178), .Y(n_1477) );
INVxp33_ASAP7_75t_SL g1558 ( .A(n_180), .Y(n_1558) );
INVxp33_ASAP7_75t_SL g629 ( .A(n_182), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_183), .A2(n_208), .B1(n_599), .B2(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_183), .A2(n_208), .B1(n_899), .B2(n_948), .Y(n_947) );
AOI21xp33_ASAP7_75t_L g1035 ( .A1(n_185), .A2(n_729), .B(n_1036), .Y(n_1035) );
INVxp67_ASAP7_75t_SL g1059 ( .A(n_185), .Y(n_1059) );
INVx1_ASAP7_75t_L g1154 ( .A(n_186), .Y(n_1154) );
INVx1_ASAP7_75t_L g1213 ( .A(n_187), .Y(n_1213) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_189), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_189), .A2(n_230), .B1(n_461), .B2(n_464), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g928 ( .A1(n_190), .A2(n_339), .B(n_929), .C(n_930), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_190), .A2(n_275), .B1(n_647), .B2(n_946), .Y(n_950) );
INVx1_ASAP7_75t_L g759 ( .A(n_191), .Y(n_759) );
INVxp33_ASAP7_75t_SL g858 ( .A(n_192), .Y(n_858) );
INVx1_ASAP7_75t_L g1049 ( .A(n_193), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_194), .A2(n_275), .B1(n_293), .B2(n_332), .Y(n_933) );
INVx1_ASAP7_75t_L g1555 ( .A(n_195), .Y(n_1555) );
INVxp33_ASAP7_75t_SL g706 ( .A(n_196), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_196), .A2(n_258), .B1(n_740), .B2(n_744), .Y(n_743) );
INVxp67_ASAP7_75t_SL g812 ( .A(n_198), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_198), .A2(n_244), .B1(n_632), .B2(n_845), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_199), .A2(n_268), .B1(n_533), .B2(n_537), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_199), .A2(n_268), .B1(n_1171), .B2(n_1172), .Y(n_1170) );
AO221x2_ASAP7_75t_L g1330 ( .A1(n_200), .A2(n_280), .B1(n_1295), .B2(n_1331), .C(n_1332), .Y(n_1330) );
INVxp33_ASAP7_75t_SL g874 ( .A(n_202), .Y(n_874) );
INVx1_ASAP7_75t_L g521 ( .A(n_203), .Y(n_521) );
INVx1_ASAP7_75t_L g1168 ( .A(n_204), .Y(n_1168) );
INVx2_ASAP7_75t_L g296 ( .A(n_206), .Y(n_296) );
INVx1_ASAP7_75t_L g328 ( .A(n_206), .Y(n_328) );
OAI211xp5_ASAP7_75t_L g480 ( .A1(n_207), .A2(n_481), .B(n_484), .C(n_485), .Y(n_480) );
INVx1_ASAP7_75t_L g509 ( .A(n_207), .Y(n_509) );
INVxp33_ASAP7_75t_SL g859 ( .A(n_210), .Y(n_859) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_211), .Y(n_372) );
INVxp33_ASAP7_75t_SL g819 ( .A(n_212), .Y(n_819) );
AO22x2_ASAP7_75t_L g795 ( .A1(n_213), .A2(n_796), .B1(n_851), .B2(n_852), .Y(n_795) );
CKINVDCx14_ASAP7_75t_R g851 ( .A(n_213), .Y(n_851) );
XNOR2xp5_ASAP7_75t_L g999 ( .A(n_214), .B(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1475 ( .A(n_216), .Y(n_1475) );
XNOR2xp5_ASAP7_75t_L g747 ( .A(n_219), .B(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g309 ( .A(n_220), .Y(n_309) );
INVx1_ASAP7_75t_L g499 ( .A(n_221), .Y(n_499) );
INVx1_ASAP7_75t_L g1047 ( .A(n_222), .Y(n_1047) );
OAI211xp5_ASAP7_75t_L g1087 ( .A1(n_223), .A2(n_484), .B(n_620), .C(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1109 ( .A(n_223), .Y(n_1109) );
INVx1_ASAP7_75t_L g1137 ( .A(n_225), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1128 ( .A1(n_226), .A2(n_1129), .B1(n_1183), .B2(n_1184), .Y(n_1128) );
INVxp67_ASAP7_75t_SL g1184 ( .A(n_226), .Y(n_1184) );
CKINVDCx16_ASAP7_75t_R g1220 ( .A(n_227), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_228), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_229), .Y(n_1081) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_230), .Y(n_338) );
INVx1_ASAP7_75t_L g917 ( .A(n_231), .Y(n_917) );
INVx1_ASAP7_75t_L g1151 ( .A(n_233), .Y(n_1151) );
INVx1_ASAP7_75t_L g803 ( .A(n_236), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_237), .A2(n_255), .B1(n_479), .B2(n_490), .Y(n_1090) );
INVx1_ASAP7_75t_L g1107 ( .A(n_237), .Y(n_1107) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_238), .Y(n_317) );
INVx1_ASAP7_75t_L g601 ( .A(n_239), .Y(n_601) );
INVx1_ASAP7_75t_L g989 ( .A(n_240), .Y(n_989) );
INVx1_ASAP7_75t_L g1214 ( .A(n_241), .Y(n_1214) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_241), .B(n_1212), .Y(n_1219) );
INVxp33_ASAP7_75t_SL g810 ( .A(n_244), .Y(n_810) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_245), .Y(n_670) );
INVx1_ASAP7_75t_L g868 ( .A(n_246), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g1493 ( .A(n_248), .Y(n_1493) );
INVx1_ASAP7_75t_L g799 ( .A(n_250), .Y(n_799) );
INVx1_ASAP7_75t_L g979 ( .A(n_251), .Y(n_979) );
AO22x2_ASAP7_75t_L g1072 ( .A1(n_252), .A2(n_1073), .B1(n_1074), .B2(n_1125), .Y(n_1072) );
INVxp67_ASAP7_75t_L g1125 ( .A(n_252), .Y(n_1125) );
CKINVDCx5p33_ASAP7_75t_R g1037 ( .A(n_253), .Y(n_1037) );
INVx1_ASAP7_75t_L g1084 ( .A(n_255), .Y(n_1084) );
INVx1_ASAP7_75t_L g1529 ( .A(n_256), .Y(n_1529) );
AOI22xp33_ASAP7_75t_L g1534 ( .A1(n_256), .A2(n_1535), .B1(n_1539), .B2(n_1584), .Y(n_1534) );
INVxp33_ASAP7_75t_L g705 ( .A(n_258), .Y(n_705) );
INVxp67_ASAP7_75t_SL g1176 ( .A(n_259), .Y(n_1176) );
INVx2_ASAP7_75t_L g299 ( .A(n_260), .Y(n_299) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_262), .Y(n_807) );
INVx1_ASAP7_75t_L g789 ( .A(n_263), .Y(n_789) );
INVxp33_ASAP7_75t_SL g881 ( .A(n_264), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_264), .A2(n_279), .B1(n_758), .B2(n_903), .Y(n_902) );
INVxp67_ASAP7_75t_SL g1015 ( .A(n_265), .Y(n_1015) );
XOR2xp5_ASAP7_75t_L g685 ( .A(n_266), .B(n_686), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g1215 ( .A(n_267), .Y(n_1215) );
INVx1_ASAP7_75t_L g692 ( .A(n_269), .Y(n_692) );
BUFx3_ASAP7_75t_L g359 ( .A(n_272), .Y(n_359) );
INVx1_ASAP7_75t_L g376 ( .A(n_272), .Y(n_376) );
BUFx3_ASAP7_75t_L g361 ( .A(n_273), .Y(n_361) );
INVx1_ASAP7_75t_L g367 ( .A(n_273), .Y(n_367) );
INVx1_ASAP7_75t_L g522 ( .A(n_274), .Y(n_522) );
XOR2xp5_ASAP7_75t_L g1540 ( .A(n_276), .B(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g752 ( .A(n_277), .Y(n_752) );
INVx1_ASAP7_75t_L g1011 ( .A(n_278), .Y(n_1011) );
INVx1_ASAP7_75t_L g876 ( .A(n_279), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_1186), .B(n_1198), .Y(n_281) );
OAI22xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_994), .B1(n_995), .B2(n_1185), .Y(n_282) );
INVx1_ASAP7_75t_L g1185 ( .A(n_283), .Y(n_1185) );
XNOR2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_793), .Y(n_283) );
XNOR2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_539), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
XNOR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_469), .Y(n_286) );
XNOR2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_342), .B1(n_348), .B2(n_394), .C(n_401), .Y(n_289) );
NAND4xp25_ASAP7_75t_L g290 ( .A(n_291), .B(n_308), .C(n_330), .D(n_339), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_301), .B1(n_302), .B2(n_307), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_292), .A2(n_331), .B1(n_521), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_292), .A2(n_331), .B1(n_751), .B2(n_789), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g1553 ( .A1(n_292), .A2(n_331), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
INVx4_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx5_ASAP7_75t_L g679 ( .A(n_293), .Y(n_679) );
OR2x6_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
AND2x4_ASAP7_75t_L g302 ( .A(n_294), .B(n_303), .Y(n_302) );
AND2x4_ASAP7_75t_L g334 ( .A(n_294), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g534 ( .A(n_294), .Y(n_534) );
AND2x4_ASAP7_75t_L g538 ( .A(n_294), .B(n_335), .Y(n_538) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g575 ( .A(n_295), .B(n_347), .Y(n_575) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
OR2x6_ASAP7_75t_L g332 ( .A(n_297), .B(n_327), .Y(n_332) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_297), .Y(n_498) );
INVx2_ASAP7_75t_SL g508 ( .A(n_297), .Y(n_508) );
INVx2_ASAP7_75t_SL g588 ( .A(n_297), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g1036 ( .A1(n_297), .A2(n_422), .B(n_1037), .Y(n_1036) );
BUFx6f_ASAP7_75t_L g1155 ( .A(n_297), .Y(n_1155) );
INVx1_ASAP7_75t_L g1480 ( .A(n_297), .Y(n_1480) );
OR2x2_ASAP7_75t_L g1486 ( .A(n_297), .B(n_1454), .Y(n_1486) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx2_ASAP7_75t_L g304 ( .A(n_299), .Y(n_304) );
INVx1_ASAP7_75t_L g313 ( .A(n_299), .Y(n_313) );
INVx1_ASAP7_75t_L g321 ( .A(n_299), .Y(n_321) );
AND2x4_ASAP7_75t_L g337 ( .A(n_299), .B(n_322), .Y(n_337) );
AND2x2_ASAP7_75t_L g415 ( .A(n_299), .B(n_300), .Y(n_415) );
INVx1_ASAP7_75t_L g306 ( .A(n_300), .Y(n_306) );
INVx2_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
INVx1_ASAP7_75t_L g329 ( .A(n_300), .Y(n_329) );
INVx1_ASAP7_75t_L g502 ( .A(n_300), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_300), .B(n_304), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_301), .A2(n_369), .B1(n_372), .B2(n_373), .Y(n_368) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_302), .A2(n_334), .B1(n_675), .B2(n_676), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_302), .A2(n_334), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_302), .A2(n_334), .B1(n_786), .B2(n_787), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_302), .A2(n_538), .B1(n_818), .B2(n_819), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_302), .A2(n_334), .B1(n_873), .B2(n_874), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g1545 ( .A1(n_302), .A2(n_538), .B1(n_1546), .B2(n_1547), .Y(n_1545) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_303), .Y(n_406) );
BUFx2_ASAP7_75t_L g425 ( .A(n_303), .Y(n_425) );
BUFx2_ASAP7_75t_L g494 ( .A(n_303), .Y(n_494) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_303), .Y(n_650) );
INVx1_ASAP7_75t_L g717 ( .A(n_303), .Y(n_717) );
INVx1_ASAP7_75t_L g724 ( .A(n_303), .Y(n_724) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_303), .Y(n_767) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_303), .B(n_1017), .Y(n_1016) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g1033 ( .A(n_304), .Y(n_1033) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AOI222xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B1(n_317), .B2(n_318), .C1(n_323), .C2(n_324), .Y(n_308) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_309), .A2(n_323), .B1(n_378), .B2(n_379), .C1(n_383), .C2(n_388), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g527 ( .A1(n_310), .A2(n_326), .B1(n_486), .B2(n_487), .C1(n_522), .C2(n_528), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_310), .A2(n_326), .B1(n_613), .B2(n_614), .Y(n_612) );
AOI222xp33_ASAP7_75t_L g875 ( .A1(n_310), .A2(n_324), .B1(n_867), .B2(n_868), .C1(n_876), .C2(n_877), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_310), .A2(n_920), .B1(n_921), .B2(n_931), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_310), .A2(n_326), .B1(n_979), .B2(n_980), .Y(n_978) );
AOI222xp33_ASAP7_75t_L g1078 ( .A1(n_310), .A2(n_319), .B1(n_326), .B2(n_1079), .C1(n_1080), .C2(n_1081), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_310), .A2(n_324), .B1(n_1136), .B2(n_1137), .Y(n_1143) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
AND2x4_ASAP7_75t_L g1552 ( .A(n_311), .B(n_314), .Y(n_1552) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g673 ( .A(n_312), .B(n_328), .Y(n_673) );
OR2x2_ASAP7_75t_L g816 ( .A(n_312), .B(n_328), .Y(n_816) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g501 ( .A(n_313), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_313), .B(n_502), .Y(n_611) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_316), .B(n_437), .Y(n_436) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_318), .A2(n_340), .B(n_670), .C(n_671), .Y(n_669) );
AOI211xp5_ASAP7_75t_L g782 ( .A1(n_318), .A2(n_340), .B(n_783), .C(n_784), .Y(n_782) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_SL g431 ( .A(n_319), .Y(n_431) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g340 ( .A(n_320), .B(n_341), .Y(n_340) );
BUFx3_ASAP7_75t_L g417 ( .A(n_320), .Y(n_417) );
BUFx3_ASAP7_75t_L g529 ( .A(n_320), .Y(n_529) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_320), .Y(n_729) );
INVx1_ASAP7_75t_L g814 ( .A(n_320), .Y(n_814) );
BUFx2_ASAP7_75t_L g879 ( .A(n_320), .Y(n_879) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g672 ( .A(n_326), .Y(n_672) );
INVx2_ASAP7_75t_L g932 ( .A(n_326), .Y(n_932) );
AOI222xp33_ASAP7_75t_L g1548 ( .A1(n_326), .A2(n_729), .B1(n_1549), .B2(n_1550), .C1(n_1551), .C2(n_1552), .Y(n_1548) );
AND2x4_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g422 ( .A(n_328), .B(n_346), .Y(n_422) );
INVx1_ASAP7_75t_L g1027 ( .A(n_329), .Y(n_1027) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_333), .B1(n_334), .B2(n_338), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_331), .A2(n_638), .B1(n_678), .B2(n_679), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_331), .A2(n_679), .B1(n_803), .B2(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_331), .A2(n_679), .B1(n_861), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_331), .A2(n_679), .B1(n_1083), .B2(n_1084), .Y(n_1082) );
INVx8_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g1196 ( .A(n_332), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g410 ( .A(n_337), .Y(n_410) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_337), .Y(n_428) );
INVx1_ASAP7_75t_L g721 ( .A(n_337), .Y(n_721) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_339), .B(n_527), .C(n_530), .Y(n_526) );
NAND4xp25_ASAP7_75t_SL g871 ( .A(n_339), .B(n_872), .C(n_875), .D(n_880), .Y(n_871) );
NAND3xp33_ASAP7_75t_L g1077 ( .A(n_339), .B(n_1078), .C(n_1082), .Y(n_1077) );
NAND4xp25_ASAP7_75t_L g1544 ( .A(n_339), .B(n_1545), .C(n_1548), .D(n_1553), .Y(n_1544) );
CKINVDCx11_ASAP7_75t_R g339 ( .A(n_340), .Y(n_339) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_340), .B(n_702), .C(n_703), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g811 ( .A1(n_340), .A2(n_812), .B(n_813), .C(n_815), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_342), .A2(n_526), .B(n_532), .Y(n_525) );
OAI31xp33_ASAP7_75t_SL g606 ( .A1(n_342), .A2(n_607), .A3(n_608), .B(n_615), .Y(n_606) );
AOI221x1_ASAP7_75t_L g855 ( .A1(n_342), .A2(n_856), .B1(n_870), .B2(n_871), .C(n_882), .Y(n_855) );
OAI31xp33_ASAP7_75t_L g926 ( .A1(n_342), .A2(n_927), .A3(n_928), .B(n_933), .Y(n_926) );
OAI31xp33_ASAP7_75t_SL g972 ( .A1(n_342), .A2(n_973), .A3(n_974), .B(n_981), .Y(n_972) );
O2A1O1Ixp33_ASAP7_75t_L g1075 ( .A1(n_342), .A2(n_1076), .B(n_1077), .C(n_1085), .Y(n_1075) );
OAI31xp33_ASAP7_75t_L g1139 ( .A1(n_342), .A2(n_1140), .A3(n_1141), .B(n_1144), .Y(n_1139) );
AOI221xp5_ASAP7_75t_L g1543 ( .A1(n_342), .A2(n_396), .B1(n_1544), .B2(n_1556), .C(n_1564), .Y(n_1543) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_343), .Y(n_342) );
AOI31xp33_ASAP7_75t_L g781 ( .A1(n_343), .A2(n_782), .A3(n_785), .B(n_788), .Y(n_781) );
OR2x6_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x4_ASAP7_75t_L g457 ( .A(n_344), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g658 ( .A(n_344), .B(n_458), .Y(n_658) );
OR2x2_ASAP7_75t_L g680 ( .A(n_344), .B(n_345), .Y(n_680) );
AND2x4_ASAP7_75t_L g1488 ( .A(n_344), .B(n_1489), .Y(n_1488) );
INVxp67_ASAP7_75t_L g1197 ( .A(n_345), .Y(n_1197) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND4xp25_ASAP7_75t_L g348 ( .A(n_349), .B(n_368), .C(n_377), .D(n_390), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_362), .B2(n_363), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_351), .A2(n_363), .B1(n_628), .B2(n_629), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_351), .A2(n_363), .B1(n_754), .B2(n_755), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_351), .A2(n_363), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_351), .A2(n_363), .B1(n_858), .B2(n_859), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g1557 ( .A1(n_351), .A2(n_363), .B1(n_1558), .B2(n_1559), .Y(n_1557) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_355), .Y(n_351) );
AND2x6_ASAP7_75t_L g373 ( .A(n_352), .B(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g1004 ( .A(n_352), .B(n_355), .Y(n_1004) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g693 ( .A(n_353), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g365 ( .A(n_354), .Y(n_365) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_354), .Y(n_371) );
AND2x2_ASAP7_75t_L g453 ( .A(n_354), .B(n_398), .Y(n_453) );
INVx2_ASAP7_75t_L g459 ( .A(n_354), .Y(n_459) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g441 ( .A(n_356), .Y(n_441) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_356), .Y(n_739) );
INVx2_ASAP7_75t_L g842 ( .A(n_356), .Y(n_842) );
INVx2_ASAP7_75t_SL g847 ( .A(n_356), .Y(n_847) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_356), .Y(n_904) );
INVx1_ASAP7_75t_L g971 ( .A(n_356), .Y(n_971) );
INVx6_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g369 ( .A(n_357), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g648 ( .A(n_357), .Y(n_648) );
BUFx2_ASAP7_75t_L g945 ( .A(n_357), .Y(n_945) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_357), .B(n_1490), .Y(n_1489) );
AND2x4_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g366 ( .A(n_359), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_359), .B(n_361), .Y(n_382) );
INVx1_ASAP7_75t_L g387 ( .A(n_360), .Y(n_387) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g375 ( .A(n_361), .B(n_376), .Y(n_375) );
CKINVDCx6p67_ASAP7_75t_R g489 ( .A(n_363), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_363), .A2(n_373), .B1(n_923), .B2(n_924), .Y(n_922) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_363), .A2(n_373), .B1(n_988), .B2(n_989), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_363), .A2(n_1003), .B1(n_1004), .B2(n_1005), .Y(n_1002) );
AND2x6_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
INVx1_ASAP7_75t_L g475 ( .A(n_364), .Y(n_475) );
AND2x2_ASAP7_75t_L g482 ( .A(n_364), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x6_ASAP7_75t_L g388 ( .A(n_365), .B(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_366), .Y(n_447) );
BUFx3_ASAP7_75t_L g463 ( .A(n_366), .Y(n_463) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_366), .Y(n_568) );
BUFx2_ASAP7_75t_L g744 ( .A(n_366), .Y(n_744) );
INVx2_ASAP7_75t_SL g775 ( .A(n_366), .Y(n_775) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_366), .Y(n_837) );
BUFx6f_ASAP7_75t_L g899 ( .A(n_366), .Y(n_899) );
HB1xp67_ASAP7_75t_L g906 ( .A(n_366), .Y(n_906) );
BUFx2_ASAP7_75t_L g1171 ( .A(n_366), .Y(n_1171) );
INVx1_ASAP7_75t_L g478 ( .A(n_367), .Y(n_478) );
INVx4_ASAP7_75t_L g479 ( .A(n_369), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_369), .A2(n_373), .B1(n_638), .B2(n_639), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_369), .A2(n_373), .B1(n_697), .B2(n_698), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_369), .A2(n_373), .B1(n_751), .B2(n_752), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_369), .A2(n_373), .B1(n_803), .B2(n_804), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_369), .A2(n_373), .B1(n_861), .B2(n_862), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_369), .A2(n_373), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1560 ( .A1(n_369), .A2(n_373), .B1(n_1555), .B2(n_1561), .Y(n_1560) );
AND2x4_ASAP7_75t_L g384 ( .A(n_370), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_SL g635 ( .A(n_370), .B(n_385), .Y(n_635) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx4_ASAP7_75t_L g490 ( .A(n_373), .Y(n_490) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_374), .Y(n_464) );
INVx2_ASAP7_75t_L g556 ( .A(n_374), .Y(n_556) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_374), .Y(n_563) );
INVx1_ASAP7_75t_L g780 ( .A(n_374), .Y(n_780) );
INVx1_ASAP7_75t_L g839 ( .A(n_374), .Y(n_839) );
INVx1_ASAP7_75t_L g850 ( .A(n_374), .Y(n_850) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g449 ( .A(n_375), .Y(n_449) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_375), .Y(n_524) );
INVx2_ASAP7_75t_L g664 ( .A(n_375), .Y(n_664) );
INVx1_ASAP7_75t_L g967 ( .A(n_375), .Y(n_967) );
INVx1_ASAP7_75t_L g477 ( .A(n_376), .Y(n_477) );
BUFx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx4f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_381), .Y(n_468) );
INVx1_ASAP7_75t_L g633 ( .A(n_381), .Y(n_633) );
INVx2_ASAP7_75t_SL g736 ( .A(n_381), .Y(n_736) );
BUFx3_ASAP7_75t_L g758 ( .A(n_381), .Y(n_758) );
INVx1_ASAP7_75t_L g919 ( .A(n_381), .Y(n_919) );
AND2x4_ASAP7_75t_L g1512 ( .A(n_381), .B(n_1497), .Y(n_1512) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_382), .Y(n_393) );
AOI222xp33_ASAP7_75t_L g863 ( .A1(n_383), .A2(n_388), .B1(n_864), .B2(n_865), .C1(n_867), .C2(n_868), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_383), .A2(n_388), .B1(n_1079), .B2(n_1081), .Y(n_1088) );
BUFx4f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_384), .A2(n_388), .B1(n_486), .B2(n_487), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_384), .A2(n_388), .B1(n_613), .B2(n_614), .Y(n_622) );
AOI222xp33_ASAP7_75t_L g798 ( .A1(n_384), .A2(n_388), .B1(n_569), .B2(n_799), .C1(n_800), .C2(n_801), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_384), .A2(n_388), .B1(n_1136), .B2(n_1137), .Y(n_1135) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g694 ( .A(n_386), .Y(n_694) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g1180 ( .A(n_387), .Y(n_1180) );
AOI222xp33_ASAP7_75t_L g630 ( .A1(n_388), .A2(n_631), .B1(n_632), .B2(n_634), .C1(n_635), .C2(n_636), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_388), .A2(n_692), .B1(n_693), .B2(n_695), .Y(n_691) );
AOI222xp33_ASAP7_75t_L g756 ( .A1(n_388), .A2(n_635), .B1(n_757), .B2(n_758), .C1(n_759), .C2(n_760), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g916 ( .A1(n_388), .A2(n_635), .B1(n_917), .B2(n_918), .C1(n_920), .C2(n_921), .Y(n_916) );
AOI222xp33_ASAP7_75t_L g984 ( .A1(n_388), .A2(n_693), .B1(n_979), .B2(n_980), .C1(n_985), .C2(n_986), .Y(n_984) );
AOI222xp33_ASAP7_75t_L g1009 ( .A1(n_388), .A2(n_635), .B1(n_758), .B2(n_1010), .C1(n_1011), .C2(n_1012), .Y(n_1009) );
AOI222xp33_ASAP7_75t_L g1562 ( .A1(n_388), .A2(n_442), .B1(n_635), .B2(n_1550), .C1(n_1551), .C2(n_1563), .Y(n_1562) );
BUFx3_ASAP7_75t_L g1182 ( .A(n_389), .Y(n_1182) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_390), .B(n_750), .C(n_753), .D(n_756), .Y(n_749) );
BUFx2_ASAP7_75t_L g869 ( .A(n_390), .Y(n_869) );
NAND4xp25_ASAP7_75t_L g1001 ( .A(n_390), .B(n_1002), .C(n_1006), .D(n_1009), .Y(n_1001) );
INVx5_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
CKINVDCx8_ASAP7_75t_R g484 ( .A(n_391), .Y(n_484) );
NOR2xp33_ASAP7_75t_SL g689 ( .A(n_391), .B(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx2_ASAP7_75t_L g443 ( .A(n_393), .Y(n_443) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_393), .Y(n_483) );
INVx1_ASAP7_75t_L g570 ( .A(n_393), .Y(n_570) );
BUFx6f_ASAP7_75t_L g1521 ( .A(n_393), .Y(n_1521) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI31xp33_ASAP7_75t_SL g616 ( .A1(n_396), .A2(n_617), .A3(n_618), .B(n_619), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g687 ( .A1(n_396), .A2(n_688), .B(n_699), .Y(n_687) );
AOI211x1_ASAP7_75t_SL g796 ( .A1(n_396), .A2(n_797), .B(n_808), .C(n_820), .Y(n_796) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_396), .Y(n_870) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
AND2x4_ASAP7_75t_L g491 ( .A(n_397), .B(n_399), .Y(n_491) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g458 ( .A(n_398), .B(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_L g1528 ( .A(n_399), .Y(n_1528) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g421 ( .A(n_400), .Y(n_421) );
OR2x6_ASAP7_75t_L g574 ( .A(n_400), .B(n_575), .Y(n_574) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_402), .B(n_423), .C(n_438), .D(n_454), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_411), .C(n_418), .Y(n_402) );
INVx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_406), .B(n_1441), .Y(n_1448) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx3_ASAP7_75t_L g1095 ( .A(n_409), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1440 ( .A(n_409), .B(n_1441), .Y(n_1440) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g584 ( .A(n_410), .Y(n_584) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_410), .Y(n_727) );
BUFx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_SL g712 ( .A(n_414), .Y(n_712) );
INVx2_ASAP7_75t_SL g1042 ( .A(n_414), .Y(n_1042) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_415), .Y(n_654) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g714 ( .A(n_417), .Y(n_714) );
AND2x4_ASAP7_75t_L g1048 ( .A(n_417), .B(n_1020), .Y(n_1048) );
NAND3xp33_ASAP7_75t_L g883 ( .A(n_418), .B(n_884), .C(n_887), .Y(n_883) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_418), .A2(n_1094), .B1(n_1102), .B2(n_1111), .C(n_1112), .Y(n_1093) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx3_ASAP7_75t_L g503 ( .A(n_420), .Y(n_503) );
AOI33xp33_ASAP7_75t_L g657 ( .A1(n_420), .A2(n_658), .A3(n_659), .B1(n_661), .B2(n_665), .B3(n_666), .Y(n_657) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_420), .B(n_763), .C(n_764), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g935 ( .A(n_420), .B(n_936), .C(n_938), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_420), .B(n_956), .C(n_958), .Y(n_955) );
NAND3xp33_ASAP7_75t_L g1565 ( .A(n_420), .B(n_1566), .C(n_1567), .Y(n_1565) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
OR2x6_ASAP7_75t_L g451 ( .A(n_421), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g512 ( .A(n_421), .B(n_452), .Y(n_512) );
OR2x2_ASAP7_75t_L g643 ( .A(n_421), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g655 ( .A(n_421), .B(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g708 ( .A(n_421), .B(n_422), .Y(n_708) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_421), .Y(n_1056) );
NAND3xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_429), .C(n_432), .Y(n_423) );
HB1xp67_ASAP7_75t_L g1096 ( .A(n_425), .Y(n_1096) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g495 ( .A(n_428), .Y(n_495) );
INVx2_ASAP7_75t_SL g886 ( .A(n_428), .Y(n_886) );
INVx4_ASAP7_75t_L g892 ( .A(n_428), .Y(n_892) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
CKINVDCx8_ASAP7_75t_R g605 ( .A(n_432), .Y(n_605) );
AOI33xp33_ASAP7_75t_L g821 ( .A1(n_432), .A2(n_822), .A3(n_823), .B1(n_827), .B2(n_830), .B3(n_831), .Y(n_821) );
NAND3xp33_ASAP7_75t_L g889 ( .A(n_432), .B(n_890), .C(n_893), .Y(n_889) );
NAND3xp33_ASAP7_75t_L g939 ( .A(n_432), .B(n_940), .C(n_941), .Y(n_939) );
NAND3xp33_ASAP7_75t_L g1568 ( .A(n_432), .B(n_1569), .C(n_1572), .Y(n_1568) );
INVx5_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx6_ASAP7_75t_L g510 ( .A(n_433), .Y(n_510) );
OR2x6_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g1441 ( .A(n_435), .B(n_1017), .Y(n_1441) );
INVx2_ASAP7_75t_L g656 ( .A(n_436), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_444), .C(n_450), .Y(n_438) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_441), .Y(n_1122) );
INVx1_ASAP7_75t_L g866 ( .A(n_442), .Y(n_866) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx3_ASAP7_75t_L g843 ( .A(n_443), .Y(n_843) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g554 ( .A(n_447), .Y(n_554) );
BUFx3_ASAP7_75t_L g1116 ( .A(n_447), .Y(n_1116) );
AND2x4_ASAP7_75t_L g1496 ( .A(n_447), .B(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g740 ( .A(n_449), .Y(n_740) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_450), .B(n_895), .C(n_896), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_451), .A2(n_456), .B1(n_545), .B2(n_557), .Y(n_544) );
INVx2_ASAP7_75t_L g731 ( .A(n_451), .Y(n_731) );
OAI22xp5_ASAP7_75t_SL g1112 ( .A1(n_451), .A2(n_456), .B1(n_1113), .B2(n_1117), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g1578 ( .A(n_451), .Y(n_1578) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g644 ( .A(n_453), .Y(n_644) );
INVx2_ASAP7_75t_SL g1516 ( .A(n_453), .Y(n_1516) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_460), .C(n_465), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_SL g511 ( .A1(n_456), .A2(n_512), .B1(n_513), .B2(n_520), .Y(n_511) );
INVx4_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx4f_ASAP7_75t_L g745 ( .A(n_457), .Y(n_745) );
BUFx4f_ASAP7_75t_L g907 ( .A(n_457), .Y(n_907) );
HB1xp67_ASAP7_75t_L g1509 ( .A(n_458), .Y(n_1509) );
AND2x4_ASAP7_75t_L g1490 ( .A(n_459), .B(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g1244 ( .A1(n_470), .A2(n_1209), .B1(n_1218), .B2(n_1245), .Y(n_1244) );
NAND3x1_ASAP7_75t_SL g471 ( .A(n_472), .B(n_492), .C(n_525), .Y(n_471) );
OAI31xp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_480), .A3(n_488), .B(n_491), .Y(n_472) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx2_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
BUFx2_ASAP7_75t_L g547 ( .A(n_476), .Y(n_547) );
INVx1_ASAP7_75t_L g560 ( .A(n_476), .Y(n_560) );
OR2x2_ASAP7_75t_L g1524 ( .A(n_476), .B(n_1498), .Y(n_1524) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x2_ASAP7_75t_L g518 ( .A(n_477), .B(n_478), .Y(n_518) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g1515 ( .A(n_483), .Y(n_1515) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_484), .B(n_627), .C(n_630), .D(n_637), .Y(n_626) );
NAND4xp25_ASAP7_75t_SL g797 ( .A(n_484), .B(n_798), .C(n_802), .D(n_805), .Y(n_797) );
NAND3xp33_ASAP7_75t_SL g915 ( .A(n_484), .B(n_916), .C(n_922), .Y(n_915) );
NAND3xp33_ASAP7_75t_SL g983 ( .A(n_484), .B(n_984), .C(n_987), .Y(n_983) );
NAND4xp25_ASAP7_75t_SL g1556 ( .A(n_484), .B(n_1557), .C(n_1560), .D(n_1562), .Y(n_1556) );
AOI211x1_ASAP7_75t_L g625 ( .A1(n_491), .A2(n_626), .B(n_640), .C(n_668), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g748 ( .A1(n_491), .A2(n_749), .B(n_761), .C(n_781), .Y(n_748) );
OAI21xp5_ASAP7_75t_L g914 ( .A1(n_491), .A2(n_915), .B(n_925), .Y(n_914) );
OAI21xp5_ASAP7_75t_SL g982 ( .A1(n_491), .A2(n_983), .B(n_990), .Y(n_982) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_503), .B1(n_504), .B2(n_510), .C(n_511), .Y(n_492) );
INVx1_ASAP7_75t_L g1108 ( .A(n_495), .Y(n_1108) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_496) );
OAI221xp5_ASAP7_75t_L g513 ( .A1(n_497), .A2(n_499), .B1(n_514), .B2(n_516), .C(n_519), .Y(n_513) );
OAI22xp33_ASAP7_75t_SL g505 ( .A1(n_500), .A2(n_506), .B1(n_507), .B2(n_509), .Y(n_505) );
INVx1_ASAP7_75t_L g590 ( .A(n_500), .Y(n_590) );
OAI21xp5_ASAP7_75t_SL g1040 ( .A1(n_500), .A2(n_1010), .B(n_1041), .Y(n_1040) );
BUFx2_ASAP7_75t_L g1476 ( .A(n_500), .Y(n_1476) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g603 ( .A(n_501), .Y(n_603) );
INVx2_ASAP7_75t_L g977 ( .A(n_501), .Y(n_977) );
OAI22xp5_ASAP7_75t_SL g1097 ( .A1(n_507), .A2(n_1098), .B1(n_1099), .B2(n_1100), .Y(n_1097) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI33xp33_ASAP7_75t_L g707 ( .A1(n_510), .A2(n_708), .A3(n_709), .B1(n_715), .B2(n_722), .B3(n_725), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_510), .B(n_960), .C(n_962), .Y(n_959) );
INVx2_ASAP7_75t_L g1157 ( .A(n_510), .Y(n_1157) );
OAI221xp5_ASAP7_75t_L g520 ( .A1(n_514), .A2(n_516), .B1(n_521), .B2(n_522), .C(n_523), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g1167 ( .A1(n_514), .A2(n_620), .B1(n_1168), .B2(n_1169), .C(n_1170), .Y(n_1167) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_515), .Y(n_1066) );
INVx2_ASAP7_75t_L g1114 ( .A(n_515), .Y(n_1114) );
INVx2_ASAP7_75t_L g1508 ( .A(n_515), .Y(n_1508) );
OAI221xp5_ASAP7_75t_L g1113 ( .A1(n_516), .A2(n_1098), .B1(n_1099), .B2(n_1114), .C(n_1115), .Y(n_1113) );
OAI221xp5_ASAP7_75t_L g1117 ( .A1(n_516), .A2(n_1080), .B1(n_1118), .B2(n_1120), .C(n_1121), .Y(n_1117) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g621 ( .A(n_517), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g1058 ( .A1(n_517), .A2(n_559), .B1(n_1037), .B2(n_1059), .C(n_1060), .Y(n_1058) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g550 ( .A(n_518), .Y(n_550) );
BUFx2_ASAP7_75t_L g1069 ( .A(n_518), .Y(n_1069) );
INVx1_ASAP7_75t_L g1134 ( .A(n_518), .Y(n_1134) );
INVx1_ASAP7_75t_L g1507 ( .A(n_518), .Y(n_1507) );
BUFx6f_ASAP7_75t_L g948 ( .A(n_524), .Y(n_948) );
INVx1_ASAP7_75t_L g1124 ( .A(n_524), .Y(n_1124) );
BUFx3_ASAP7_75t_L g1583 ( .A(n_524), .Y(n_1583) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x6_ASAP7_75t_L g1443 ( .A(n_529), .B(n_1441), .Y(n_1443) );
NAND2x1p5_ASAP7_75t_L g1459 ( .A(n_529), .B(n_1453), .Y(n_1459) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g1161 ( .A(n_535), .Y(n_1161) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g580 ( .A(n_536), .Y(n_580) );
INVx1_ASAP7_75t_L g595 ( .A(n_536), .Y(n_595) );
INVx5_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_684), .B1(n_791), .B2(n_792), .Y(n_539) );
INVx1_ASAP7_75t_L g791 ( .A(n_540), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_623), .B1(n_624), .B2(n_683), .Y(n_540) );
INVx1_ASAP7_75t_L g683 ( .A(n_541), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_606), .C(n_616), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_571), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_548), .B2(n_551), .C(n_552), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_546), .A2(n_551), .B1(n_587), .B2(n_589), .Y(n_586) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g1514 ( .A(n_554), .Y(n_1514) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g900 ( .A(n_556), .Y(n_900) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B1(n_562), .B2(n_564), .C(n_565), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g734 ( .A(n_568), .Y(n_734) );
BUFx3_ASAP7_75t_L g1119 ( .A(n_568), .Y(n_1119) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI33xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .A3(n_586), .B1(n_591), .B2(n_597), .B3(n_605), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g1158 ( .A1(n_574), .A2(n_1071), .B1(n_1159), .B2(n_1167), .Y(n_1158) );
OAI33xp33_ASAP7_75t_L g1460 ( .A1(n_574), .A2(n_605), .A3(n_1461), .B1(n_1465), .B2(n_1473), .B3(n_1478), .Y(n_1460) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_581), .B2(n_585), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g1468 ( .A(n_580), .Y(n_1468) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g600 ( .A(n_584), .Y(n_600) );
INVx2_ASAP7_75t_L g829 ( .A(n_584), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g591 ( .A1(n_587), .A2(n_592), .B1(n_593), .B2(n_596), .Y(n_591) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g1461 ( .A1(n_589), .A2(n_1462), .B1(n_1463), .B2(n_1464), .Y(n_1461) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g1142 ( .A(n_590), .Y(n_1142) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g1150 ( .A(n_595), .Y(n_1150) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_601), .B1(n_602), .B2(n_604), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI22xp33_ASAP7_75t_SL g1153 ( .A1(n_602), .A2(n_1154), .B1(n_1155), .B2(n_1156), .Y(n_1153) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g929 ( .A(n_603), .Y(n_929) );
INVx1_ASAP7_75t_L g1111 ( .A(n_605), .Y(n_1111) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_609), .Y(n_1110) );
BUFx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g1101 ( .A(n_610), .Y(n_1101) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI21xp33_ASAP7_75t_SL g1175 ( .A1(n_620), .A2(n_1176), .B(n_1177), .Y(n_1175) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g682 ( .A(n_625), .Y(n_682) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_657), .Y(n_640) );
AOI33xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_645), .A3(n_646), .B1(n_649), .B2(n_651), .B3(n_655), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_642), .B(n_772), .C(n_773), .Y(n_771) );
NAND3xp33_ASAP7_75t_L g943 ( .A(n_642), .B(n_944), .C(n_947), .Y(n_943) );
NAND3xp33_ASAP7_75t_L g963 ( .A(n_642), .B(n_964), .C(n_965), .Y(n_963) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_SL g660 ( .A(n_648), .Y(n_660) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_SL g667 ( .A(n_653), .Y(n_667) );
INVx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g770 ( .A(n_654), .Y(n_770) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_654), .B(n_1017), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g1105 ( .A(n_654), .Y(n_1105) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_655), .B(n_766), .C(n_769), .Y(n_765) );
INVx1_ASAP7_75t_L g1043 ( .A(n_656), .Y(n_1043) );
NAND3xp33_ASAP7_75t_L g776 ( .A(n_658), .B(n_777), .C(n_778), .Y(n_776) );
AOI33xp33_ASAP7_75t_L g834 ( .A1(n_658), .A2(n_731), .A3(n_835), .B1(n_840), .B2(n_844), .B3(n_848), .Y(n_834) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_658), .B(n_950), .C(n_951), .Y(n_949) );
NAND3xp33_ASAP7_75t_L g968 ( .A(n_658), .B(n_969), .C(n_970), .Y(n_968) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g1062 ( .A(n_663), .Y(n_1062) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g1526 ( .A(n_664), .B(n_1498), .Y(n_1526) );
AOI31xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_674), .A3(n_677), .B(n_680), .Y(n_668) );
AO21x1_ASAP7_75t_SL g700 ( .A1(n_680), .A2(n_701), .B(n_704), .Y(n_700) );
AOI31xp33_ASAP7_75t_L g808 ( .A1(n_680), .A2(n_809), .A3(n_811), .B(n_817), .Y(n_808) );
INVx1_ASAP7_75t_L g792 ( .A(n_684), .Y(n_792) );
AO22x2_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_746), .B1(n_747), .B2(n_790), .Y(n_684) );
INVx1_ASAP7_75t_L g790 ( .A(n_685), .Y(n_790) );
NAND4xp25_ASAP7_75t_L g686 ( .A(n_687), .B(n_700), .C(n_707), .D(n_730), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_696), .Y(n_688) );
BUFx2_ASAP7_75t_L g822 ( .A(n_708), .Y(n_822) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_L g824 ( .A(n_712), .Y(n_824) );
AND2x4_ASAP7_75t_L g1446 ( .A(n_712), .B(n_1441), .Y(n_1446) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g1571 ( .A(n_720), .Y(n_1571) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g1022 ( .A(n_721), .Y(n_1022) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g832 ( .A(n_724), .Y(n_832) );
INVx1_ASAP7_75t_L g937 ( .A(n_724), .Y(n_937) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g768 ( .A(n_727), .Y(n_768) );
INVx2_ASAP7_75t_L g957 ( .A(n_727), .Y(n_957) );
INVx2_ASAP7_75t_L g961 ( .A(n_727), .Y(n_961) );
INVx2_ASAP7_75t_L g1164 ( .A(n_727), .Y(n_1164) );
BUFx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_SL g826 ( .A(n_729), .Y(n_826) );
AOI33xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .A3(n_737), .B1(n_741), .B2(n_743), .B3(n_745), .Y(n_730) );
INVx1_ASAP7_75t_L g1063 ( .A(n_731), .Y(n_1063) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g946 ( .A(n_736), .Y(n_946) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx4_ASAP7_75t_L g742 ( .A(n_739), .Y(n_742) );
CKINVDCx5p33_ASAP7_75t_R g1071 ( .A(n_745), .Y(n_1071) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND4xp25_ASAP7_75t_L g761 ( .A(n_762), .B(n_765), .C(n_771), .D(n_776), .Y(n_761) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AO22x1_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_911), .B1(n_992), .B2(n_993), .Y(n_793) );
INVx1_ASAP7_75t_L g992 ( .A(n_794), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_853), .B1(n_854), .B2(n_910), .Y(n_794) );
INVx1_ASAP7_75t_L g910 ( .A(n_795), .Y(n_910) );
INVx1_ASAP7_75t_L g852 ( .A(n_796), .Y(n_852) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_834), .Y(n_820) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g942 ( .A(n_826), .Y(n_942) );
INVx2_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g833 ( .A(n_829), .Y(n_833) );
BUFx4f_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
BUFx6f_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g1172 ( .A(n_850), .Y(n_1172) );
OAI22xp33_ASAP7_75t_L g1332 ( .A1(n_851), .A2(n_1333), .B1(n_1334), .B2(n_1335), .Y(n_1332) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g909 ( .A(n_855), .Y(n_909) );
NAND4xp25_ASAP7_75t_L g856 ( .A(n_857), .B(n_860), .C(n_863), .D(n_869), .Y(n_856) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AOI221x1_ASAP7_75t_L g1000 ( .A1(n_870), .A2(n_1001), .B1(n_1013), .B2(n_1054), .C(n_1057), .Y(n_1000) );
INVx1_ASAP7_75t_L g1092 ( .A(n_870), .Y(n_1092) );
OAI31xp33_ASAP7_75t_L g1130 ( .A1(n_870), .A2(n_1131), .A3(n_1132), .B(n_1138), .Y(n_1130) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g888 ( .A(n_878), .Y(n_888) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND4xp25_ASAP7_75t_L g882 ( .A(n_883), .B(n_889), .C(n_894), .D(n_901), .Y(n_882) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g1478 ( .A1(n_892), .A2(n_1479), .B1(n_1481), .B2(n_1482), .Y(n_1478) );
INVx2_ASAP7_75t_SL g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
BUFx3_ASAP7_75t_L g1582 ( .A(n_899), .Y(n_1582) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_905), .C(n_907), .Y(n_901) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
NAND3xp33_ASAP7_75t_L g1579 ( .A(n_907), .B(n_1580), .C(n_1581), .Y(n_1579) );
INVx2_ASAP7_75t_L g993 ( .A(n_911), .Y(n_993) );
XOR2x2_ASAP7_75t_L g911 ( .A(n_912), .B(n_952), .Y(n_911) );
NAND3x1_ASAP7_75t_L g913 ( .A(n_914), .B(n_926), .C(n_934), .Y(n_913) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g986 ( .A(n_919), .Y(n_986) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
AND4x1_ASAP7_75t_L g934 ( .A(n_935), .B(n_939), .C(n_943), .D(n_949), .Y(n_934) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_945), .Y(n_1174) );
XOR2xp5_ASAP7_75t_L g952 ( .A(n_953), .B(n_991), .Y(n_952) );
NAND3xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_972), .C(n_982), .Y(n_953) );
AND4x1_ASAP7_75t_L g954 ( .A(n_955), .B(n_959), .C(n_963), .D(n_968), .Y(n_954) );
INVx1_ASAP7_75t_L g1152 ( .A(n_957), .Y(n_1152) );
HB1xp67_ASAP7_75t_L g1471 ( .A(n_961), .Y(n_1471) );
INVx2_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
OR2x6_ASAP7_75t_L g1045 ( .A(n_977), .B(n_1029), .Y(n_1045) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
XOR2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_1127), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_998), .B1(n_1072), .B2(n_1126), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
AOI222xp33_ASAP7_75t_L g1046 ( .A1(n_1007), .A2(n_1047), .B1(n_1048), .B2(n_1049), .C1(n_1050), .C2(n_1051), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1023), .C(n_1046), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_1015), .A2(n_1016), .B1(n_1018), .B2(n_1019), .Y(n_1014) );
INVx2_ASAP7_75t_L g1021 ( .A(n_1017), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1022), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
NOR3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1039), .C(n_1044), .Y(n_1023) );
NAND2x1p5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1028), .Y(n_1025) );
NAND2x1_ASAP7_75t_SL g1452 ( .A(n_1026), .B(n_1453), .Y(n_1452) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
OR2x6_ASAP7_75t_L g1032 ( .A(n_1029), .B(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1029), .Y(n_1053) );
INVx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1033), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1038), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_1042), .B(n_1053), .Y(n_1052) );
BUFx2_ASAP7_75t_L g1573 ( .A(n_1042), .Y(n_1573) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
OAI221xp5_ASAP7_75t_SL g1064 ( .A1(n_1047), .A2(n_1049), .B1(n_1065), .B2(n_1067), .C(n_1070), .Y(n_1064) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
CKINVDCx8_ASAP7_75t_R g1055 ( .A(n_1056), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_1058), .A2(n_1063), .B1(n_1064), .B2(n_1071), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1061 ( .A(n_1062), .Y(n_1061) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx2_ASAP7_75t_SL g1068 ( .A(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1072), .Y(n_1126) );
INVx2_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1093), .Y(n_1074) );
AOI21xp5_ASAP7_75t_L g1085 ( .A1(n_1086), .A2(n_1089), .B(n_1092), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1091), .Y(n_1089) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
OAI22xp33_ASAP7_75t_SL g1106 ( .A1(n_1107), .A2(n_1108), .B1(n_1109), .B2(n_1110), .Y(n_1106) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1129), .Y(n_1183) );
NAND3xp33_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1139), .C(n_1145), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
NOR3xp33_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1158), .C(n_1173), .Y(n_1145) );
NOR3xp33_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1153), .C(n_1157), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_1148), .A2(n_1149), .B1(n_1151), .B2(n_1152), .Y(n_1147) );
BUFx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
BUFx2_ASAP7_75t_L g1462 ( .A(n_1155), .Y(n_1462) );
OAI221xp5_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1162), .B1(n_1163), .B2(n_1165), .C(n_1166), .Y(n_1159) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1180), .Y(n_1502) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1182), .B(n_1490), .Y(n_1504) );
BUFx2_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
INVx3_ASAP7_75t_SL g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_SL g1188 ( .A(n_1189), .Y(n_1188) );
AND2x4_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1195), .Y(n_1189) );
AND2x4_ASAP7_75t_L g1533 ( .A(n_1190), .B(n_1196), .Y(n_1533) );
NOR2xp33_ASAP7_75t_SL g1190 ( .A(n_1191), .B(n_1193), .Y(n_1190) );
INVx1_ASAP7_75t_SL g1538 ( .A(n_1191), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1585 ( .A(n_1191), .B(n_1193), .Y(n_1585) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1193), .B(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI221xp5_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1430), .B1(n_1432), .B2(n_1530), .C(n_1534), .Y(n_1198) );
AND3x1_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1388), .C(n_1418), .Y(n_1199) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_1201), .A2(n_1288), .B1(n_1296), .B2(n_1339), .C(n_1366), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1273), .Y(n_1201) );
O2A1O1Ixp33_ASAP7_75t_L g1202 ( .A1(n_1203), .A2(n_1254), .B(n_1257), .C(n_1262), .Y(n_1202) );
AOI21xp5_ASAP7_75t_L g1400 ( .A1(n_1203), .A2(n_1401), .B(n_1403), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1231), .Y(n_1203) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1204), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1204), .B(n_1286), .Y(n_1387) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1204), .Y(n_1403) );
INVx2_ASAP7_75t_SL g1204 ( .A(n_1205), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1205), .B(n_1276), .Y(n_1279) );
AND2x4_ASAP7_75t_L g1287 ( .A(n_1205), .B(n_1258), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1205), .B(n_1259), .Y(n_1301) );
HB1xp67_ASAP7_75t_L g1317 ( .A(n_1205), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1205), .B(n_1289), .Y(n_1323) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_1206), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1206), .B(n_1258), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1206), .B(n_1259), .Y(n_1306) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1221), .Y(n_1206) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_1208), .A2(n_1215), .B1(n_1216), .B2(n_1220), .Y(n_1207) );
BUFx3_ASAP7_75t_L g1334 ( .A(n_1208), .Y(n_1334) );
BUFx6f_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1211), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1210), .B(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1210), .Y(n_1238) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1211), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1214), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1214), .Y(n_1225) );
HB1xp67_ASAP7_75t_L g1335 ( .A(n_1216), .Y(n_1335) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1219), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_1222), .A2(n_1227), .B1(n_1228), .B2(n_1230), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
BUFx3_ASAP7_75t_L g1331 ( .A(n_1223), .Y(n_1331) );
AND2x4_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1226), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1224), .B(n_1226), .Y(n_1242) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
AND2x4_ASAP7_75t_L g1229 ( .A(n_1225), .B(n_1226), .Y(n_1229) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1228), .Y(n_1295) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1246), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1232), .B(n_1286), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1232), .B(n_1251), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1232), .B(n_1265), .Y(n_1384) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
NOR2xp33_ASAP7_75t_L g1352 ( .A(n_1233), .B(n_1286), .Y(n_1352) );
NOR2xp33_ASAP7_75t_L g1389 ( .A(n_1233), .B(n_1390), .Y(n_1389) );
OR2x2_ASAP7_75t_L g1429 ( .A(n_1233), .B(n_1329), .Y(n_1429) );
OR2x2_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1243), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1234), .B(n_1243), .Y(n_1256) );
INVx2_ASAP7_75t_L g1270 ( .A(n_1234), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1234), .B(n_1284), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1234), .B(n_1283), .Y(n_1349) );
NOR2xp33_ASAP7_75t_L g1381 ( .A(n_1234), .B(n_1284), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1241), .Y(n_1234) );
AND2x4_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1238), .Y(n_1236) );
OAI21xp33_ASAP7_75t_SL g1584 ( .A1(n_1237), .A2(n_1538), .B(n_1585), .Y(n_1584) );
AND2x4_ASAP7_75t_L g1239 ( .A(n_1238), .B(n_1240), .Y(n_1239) );
BUFx2_ASAP7_75t_L g1293 ( .A(n_1239), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1243), .B(n_1270), .Y(n_1269) );
INVx2_ASAP7_75t_SL g1283 ( .A(n_1243), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1243), .B(n_1251), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1243), .B(n_1284), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1246), .B(n_1256), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1246), .B(n_1269), .Y(n_1300) );
INVxp67_ASAP7_75t_SL g1350 ( .A(n_1246), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1250), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1247), .B(n_1256), .Y(n_1266) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1247), .Y(n_1276) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1247), .Y(n_1286) );
BUFx2_ASAP7_75t_L g1305 ( .A(n_1247), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1247), .B(n_1284), .Y(n_1329) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1247), .B(n_1311), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1249), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1250), .B(n_1269), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1250), .B(n_1256), .Y(n_1313) );
NOR2x1_ASAP7_75t_L g1360 ( .A(n_1250), .B(n_1283), .Y(n_1360) );
NOR2xp33_ASAP7_75t_L g1413 ( .A(n_1250), .B(n_1270), .Y(n_1413) );
BUFx2_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVxp67_ASAP7_75t_L g1265 ( .A(n_1251), .Y(n_1265) );
BUFx3_ASAP7_75t_L g1284 ( .A(n_1251), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1253), .Y(n_1251) );
AOI21xp5_ASAP7_75t_L g1423 ( .A1(n_1254), .A2(n_1403), .B(n_1424), .Y(n_1423) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1256), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1256), .B(n_1328), .Y(n_1327) );
OAI221xp5_ASAP7_75t_L g1346 ( .A1(n_1256), .A2(n_1347), .B1(n_1348), .B2(n_1350), .C(n_1351), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1256), .B(n_1286), .Y(n_1409) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1257), .Y(n_1416) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1257), .B(n_1305), .Y(n_1421) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1258), .B(n_1291), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1258), .B(n_1373), .Y(n_1372) );
A2O1A1Ixp33_ASAP7_75t_SL g1418 ( .A1(n_1258), .A2(n_1336), .B(n_1419), .C(n_1420), .Y(n_1418) );
INVx3_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1259), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1345 ( .A(n_1259), .B(n_1291), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1259), .B(n_1290), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1261), .Y(n_1259) );
AOI21xp5_ASAP7_75t_L g1262 ( .A1(n_1263), .A2(n_1267), .B(n_1271), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
AOI22xp5_ASAP7_75t_L g1405 ( .A1(n_1264), .A2(n_1320), .B1(n_1406), .B2(n_1408), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1266), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1265), .B(n_1269), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1265), .B(n_1349), .Y(n_1399) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1269), .B(n_1286), .Y(n_1395) );
A2O1A1Ixp33_ASAP7_75t_L g1354 ( .A1(n_1270), .A2(n_1355), .B(n_1358), .C(n_1361), .Y(n_1354) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
O2A1O1Ixp33_ASAP7_75t_L g1326 ( .A1(n_1272), .A2(n_1327), .B(n_1330), .C(n_1336), .Y(n_1326) );
OAI21xp5_ASAP7_75t_L g1367 ( .A1(n_1272), .A2(n_1275), .B(n_1368), .Y(n_1367) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1272), .B(n_1276), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1272), .B(n_1426), .Y(n_1425) );
AOI211xp5_ASAP7_75t_SL g1273 ( .A1(n_1274), .A2(n_1275), .B(n_1278), .C(n_1280), .Y(n_1273) );
A2O1A1Ixp33_ASAP7_75t_SL g1397 ( .A1(n_1274), .A2(n_1396), .B(n_1398), .C(n_1400), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1277), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1276), .B(n_1413), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1277), .B(n_1279), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1422 ( .A(n_1277), .B(n_1315), .Y(n_1422) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1279), .Y(n_1347) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1285), .Y(n_1280) );
OAI221xp5_ASAP7_75t_L g1296 ( .A1(n_1281), .A2(n_1297), .B1(n_1318), .B2(n_1319), .C(n_1321), .Y(n_1296) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1284), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1284), .B(n_1299), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1284), .B(n_1409), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1287), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1286), .B(n_1311), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1286), .B(n_1315), .Y(n_1314) );
OAI21xp33_ASAP7_75t_L g1382 ( .A1(n_1286), .A2(n_1309), .B(n_1383), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1287), .B(n_1289), .Y(n_1320) );
AOI221xp5_ASAP7_75t_L g1378 ( .A1(n_1287), .A2(n_1322), .B1(n_1379), .B2(n_1382), .C(n_1385), .Y(n_1378) );
AOI21xp5_ASAP7_75t_L g1394 ( .A1(n_1287), .A2(n_1395), .B(n_1396), .Y(n_1394) );
INVx2_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1289), .B(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1290), .Y(n_1338) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1291), .Y(n_1318) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1291), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1294), .Y(n_1291) );
AOI22xp5_ASAP7_75t_L g1339 ( .A1(n_1297), .A2(n_1340), .B1(n_1343), .B2(n_1354), .Y(n_1339) );
AND3x1_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1302), .C(n_1312), .Y(n_1297) );
OAI21xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1300), .B(n_1301), .Y(n_1298) );
AOI221xp5_ASAP7_75t_L g1321 ( .A1(n_1300), .A2(n_1322), .B1(n_1324), .B2(n_1325), .C(n_1326), .Y(n_1321) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1301), .B(n_1357), .Y(n_1356) );
A2O1A1Ixp33_ASAP7_75t_L g1410 ( .A1(n_1301), .A2(n_1330), .B(n_1411), .C(n_1414), .Y(n_1410) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_1303), .A2(n_1306), .B1(n_1307), .B2(n_1310), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
AOI21xp5_ASAP7_75t_L g1414 ( .A1(n_1304), .A2(n_1308), .B(n_1383), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1306), .Y(n_1304) );
INVx2_ASAP7_75t_L g1357 ( .A(n_1305), .Y(n_1357) );
NAND2xp5_ASAP7_75t_SL g1380 ( .A(n_1305), .B(n_1381), .Y(n_1380) );
CKINVDCx5p33_ASAP7_75t_R g1377 ( .A(n_1306), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1309), .Y(n_1307) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1310), .Y(n_1393) );
OAI21xp33_ASAP7_75t_L g1312 ( .A1(n_1313), .A2(n_1314), .B(n_1316), .Y(n_1312) );
AOI221xp5_ASAP7_75t_L g1370 ( .A1(n_1313), .A2(n_1314), .B1(n_1325), .B2(n_1371), .C(n_1374), .Y(n_1370) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1314), .Y(n_1392) );
INVxp67_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
NOR2xp33_ASAP7_75t_L g1428 ( .A(n_1317), .B(n_1429), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1318), .B(n_1365), .Y(n_1364) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1320), .B(n_1324), .Y(n_1417) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1325), .Y(n_1407) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1330), .B(n_1337), .Y(n_1336) );
INVx3_ASAP7_75t_L g1342 ( .A(n_1330), .Y(n_1342) );
AOI31xp33_ASAP7_75t_L g1366 ( .A1(n_1330), .A2(n_1367), .A3(n_1370), .B(n_1378), .Y(n_1366) );
INVx3_ASAP7_75t_L g1396 ( .A(n_1330), .Y(n_1396) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1334), .Y(n_1431) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
AOI211xp5_ASAP7_75t_L g1343 ( .A1(n_1338), .A2(n_1344), .B(n_1346), .C(n_1353), .Y(n_1343) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1338), .Y(n_1376) );
NAND3xp33_ASAP7_75t_SL g1386 ( .A(n_1338), .B(n_1349), .C(n_1387), .Y(n_1386) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
NOR2xp33_ASAP7_75t_L g1374 ( .A(n_1348), .B(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
AOI21xp33_ASAP7_75t_L g1415 ( .A1(n_1353), .A2(n_1416), .B(n_1417), .Y(n_1415) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1357), .B(n_1360), .Y(n_1359) );
OR2x2_ASAP7_75t_L g1398 ( .A(n_1357), .B(n_1399), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1357), .B(n_1381), .Y(n_1402) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1364), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1365), .B(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1377), .Y(n_1375) );
A2O1A1Ixp33_ASAP7_75t_L g1391 ( .A1(n_1377), .A2(n_1392), .B(n_1393), .C(n_1394), .Y(n_1391) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
O2A1O1Ixp33_ASAP7_75t_L g1388 ( .A1(n_1389), .A2(n_1391), .B(n_1397), .C(n_1404), .Y(n_1388) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1398), .Y(n_1419) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1399), .Y(n_1426) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
NAND3xp33_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1410), .C(n_1415), .Y(n_1404) );
INVxp67_ASAP7_75t_SL g1411 ( .A(n_1412), .Y(n_1411) );
OAI211xp5_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1422), .B(n_1423), .C(n_1427), .Y(n_1420) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx2_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
XNOR2x1_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1529), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1483), .Y(n_1434) );
NOR3xp33_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1449), .C(n_1460), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1444), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1437 ( .A1(n_1438), .A2(n_1439), .B1(n_1442), .B2(n_1443), .Y(n_1437) );
BUFx2_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
OAI221xp5_ASAP7_75t_L g1506 ( .A1(n_1442), .A2(n_1445), .B1(n_1507), .B2(n_1508), .C(n_1509), .Y(n_1506) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_1445), .A2(n_1446), .B1(n_1447), .B2(n_1448), .Y(n_1444) );
INVx2_ASAP7_75t_SL g1450 ( .A(n_1451), .Y(n_1450) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
NAND2x1p5_ASAP7_75t_L g1456 ( .A(n_1453), .B(n_1457), .Y(n_1456) );
INVx3_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
BUFx4f_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
BUFx2_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
OAI22xp5_ASAP7_75t_L g1465 ( .A1(n_1466), .A2(n_1469), .B1(n_1470), .B2(n_1472), .Y(n_1465) );
INVx2_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
INVx2_ASAP7_75t_L g1474 ( .A(n_1467), .Y(n_1474) );
INVx2_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
OAI22xp5_ASAP7_75t_L g1473 ( .A1(n_1474), .A2(n_1475), .B1(n_1476), .B2(n_1477), .Y(n_1473) );
AOI211xp5_ASAP7_75t_L g1495 ( .A1(n_1475), .A2(n_1496), .B(n_1499), .C(n_1505), .Y(n_1495) );
AOI221xp5_ASAP7_75t_L g1510 ( .A1(n_1477), .A2(n_1511), .B1(n_1513), .B2(n_1517), .C(n_1518), .Y(n_1510) );
INVx2_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
AOI22xp33_ASAP7_75t_L g1522 ( .A1(n_1481), .A2(n_1482), .B1(n_1523), .B2(n_1525), .Y(n_1522) );
AOI21xp33_ASAP7_75t_SL g1483 ( .A1(n_1484), .A2(n_1493), .B(n_1494), .Y(n_1483) );
INVx5_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
AND2x4_ASAP7_75t_L g1485 ( .A(n_1486), .B(n_1487), .Y(n_1485) );
INVx2_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
AND2x4_ASAP7_75t_L g1501 ( .A(n_1490), .B(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1490), .Y(n_1520) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
AOI31xp33_ASAP7_75t_L g1494 ( .A1(n_1495), .A2(n_1510), .A3(n_1522), .B(n_1527), .Y(n_1494) );
INVx2_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
INVx3_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
BUFx6f_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
AND2x4_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1521), .Y(n_1518) );
INVx1_ASAP7_75t_SL g1519 ( .A(n_1520), .Y(n_1519) );
BUFx6f_ASAP7_75t_L g1576 ( .A(n_1521), .Y(n_1576) );
INVx6_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
INVx4_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
INVx2_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx4_ASAP7_75t_SL g1530 ( .A(n_1531), .Y(n_1530) );
BUFx3_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
BUFx2_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
CKINVDCx5p33_ASAP7_75t_R g1536 ( .A(n_1537), .Y(n_1536) );
INVxp33_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
HB1xp67_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
NAND4xp25_ASAP7_75t_SL g1564 ( .A(n_1565), .B(n_1568), .C(n_1574), .D(n_1579), .Y(n_1564) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
NAND3xp33_ASAP7_75t_L g1574 ( .A(n_1575), .B(n_1577), .C(n_1578), .Y(n_1574) );
endmodule