module real_jpeg_12250_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_298, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;
input n_298;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_221;
wire n_292;
wire n_166;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_2),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_2),
.A2(n_22),
.B1(n_27),
.B2(n_40),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_2),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_287)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_22),
.B1(n_27),
.B2(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_4),
.A2(n_33),
.B1(n_37),
.B2(n_100),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_100),
.Y(n_176)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_33),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_43),
.B1(n_57),
.B2(n_58),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_43),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_7),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_10),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_28),
.B1(n_51),
.B2(n_52),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_10),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_10),
.A2(n_28),
.B1(n_57),
.B2(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_10),
.B(n_69),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_10),
.B(n_22),
.C(n_36),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_10),
.B(n_85),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_10),
.B(n_38),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_10),
.A2(n_58),
.B(n_71),
.C(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_10),
.B(n_56),
.Y(n_196)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_276),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_121),
.B(n_274),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_101),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_16),
.B(n_101),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_61),
.C(n_78),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_17),
.A2(n_18),
.B1(n_61),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_19),
.A2(n_20),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_20),
.A2(n_45),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_20),
.B(n_179),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_20),
.A2(n_29),
.B1(n_45),
.B2(n_265),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_26),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_21),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_21),
.B(n_26),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_21),
.A2(n_210),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_22),
.B(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_25),
.B(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_25),
.B(n_82),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_25),
.A2(n_81),
.B(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_28),
.A2(n_37),
.B(n_72),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_28),
.B(n_54),
.C(n_58),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_29),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_39),
.B(n_41),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_30),
.A2(n_66),
.B(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_31),
.B(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_31),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_31),
.B(n_65),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_33),
.A2(n_37),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_33),
.B(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_38),
.B(n_138),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_39),
.A2(n_63),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_41),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_41),
.B(n_149),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_59),
.B(n_60),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_48),
.B(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_49),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_49),
.B(n_109),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_52),
.B(n_208),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_56),
.B(n_99),
.Y(n_216)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_59),
.A2(n_238),
.B(n_287),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_61),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B(n_77),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_67),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_63),
.B(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_64),
.B(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_73),
.Y(n_67)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_69),
.B(n_176),
.Y(n_175)
);

NAND2x1_ASAP7_75t_SL g227 ( 
.A(n_69),
.B(n_93),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_69),
.A2(n_92),
.B(n_93),
.Y(n_239)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_76),
.Y(n_89)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_73),
.B(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_73),
.B(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_74),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_104),
.B1(n_105),
.B2(n_120),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_77),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_77),
.B(n_102),
.C(n_104),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_78),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_88),
.C(n_94),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_79),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_80),
.B(n_86),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_81),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_88),
.A2(n_94),
.B1(n_95),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_88),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_89),
.B(n_192),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_91),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_98),
.B(n_108),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_106),
.B(n_115),
.C(n_116),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_106),
.A2(n_107),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_111),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_114),
.A2(n_115),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_114),
.B(n_214),
.C(n_219),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_114),
.A2(n_115),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_116),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_268),
.B(n_273),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_255),
.B(n_267),
.Y(n_122)
);

AOI321xp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_222),
.A3(n_248),
.B1(n_253),
.B2(n_254),
.C(n_298),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_199),
.B(n_221),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_183),
.B(n_198),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_170),
.B(n_182),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_150),
.B(n_169),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_143),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_143),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_142),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_130),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_140),
.C(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_163),
.B(n_168),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_158),
.B(n_162),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_161),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_166),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_172),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_177),
.C(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_197),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_197),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_188),
.C(n_190),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_195),
.C(n_196),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_201),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_212),
.B2(n_213),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_205),
.C(n_212),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_211),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_211),
.Y(n_229)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_243),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_243),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_231),
.C(n_242),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.C(n_229),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_226),
.CI(n_229),
.CON(n_245),
.SN(n_245)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_227),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_242),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_239),
.C(n_240),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_245),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_245),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_252),
.Y(n_253)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_264),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_294),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_288),
.B1(n_289),
.B2(n_293),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_286),
.Y(n_293)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);


endmodule