module fake_jpeg_21578_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_46),
.C(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_71),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_48),
.B1(n_59),
.B2(n_37),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_69),
.B1(n_50),
.B2(n_1),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_47),
.B1(n_48),
.B2(n_38),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_61),
.B1(n_64),
.B2(n_70),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_44),
.B(n_40),
.C(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_0),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_73),
.B1(n_10),
.B2(n_14),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_2),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_3),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_4),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_84),
.B1(n_6),
.B2(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_5),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_6),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_23),
.C(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_15),
.Y(n_98)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_9),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_26),
.B(n_27),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_72),
.B1(n_83),
.B2(n_18),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_98),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_107),
.B1(n_101),
.B2(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_105),
.B(n_101),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_108),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_86),
.Y(n_111)
);

OAI321xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_86),
.A3(n_102),
.B1(n_90),
.B2(n_91),
.C(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_29),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_30),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_114),
.B(n_31),
.Y(n_115)
);


endmodule