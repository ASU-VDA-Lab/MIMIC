module fake_jpeg_29289_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_9),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_2),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_0),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_1),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_44),
.C(n_29),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_2),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_20),
.Y(n_57)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_66),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_19),
.B1(n_18),
.B2(n_15),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_80),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_34),
.B1(n_35),
.B2(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_29),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_16),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_12),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_22),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_26),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_37),
.B(n_61),
.Y(n_108)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_50),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_54),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_53),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_54),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_50),
.A3(n_14),
.B1(n_22),
.B2(n_37),
.Y(n_103)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_53),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_63),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_90),
.B(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_24),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_109),
.Y(n_121)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_104),
.B(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_115),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_93),
.B1(n_103),
.B2(n_78),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_97),
.B1(n_48),
.B2(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_85),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_100),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_79),
.B(n_77),
.Y(n_132)
);

OAI22x1_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_71),
.B1(n_26),
.B2(n_67),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_108),
.B(n_76),
.C(n_22),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_133),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_134),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_91),
.C(n_83),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_110),
.A3(n_121),
.B1(n_120),
.B2(n_113),
.C1(n_116),
.C2(n_119),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_111),
.A3(n_110),
.B1(n_124),
.B2(n_114),
.C1(n_131),
.C2(n_117),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_115),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_136),
.C(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_144),
.A2(n_124),
.B1(n_112),
.B2(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_118),
.B(n_131),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_141),
.B(n_11),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_8),
.B(n_7),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_155),
.B(n_92),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_154),
.A2(n_8),
.B(n_131),
.C(n_4),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_139),
.B(n_136),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_153),
.A2(n_139),
.B(n_145),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_157),
.A3(n_158),
.B1(n_159),
.B2(n_76),
.C1(n_24),
.C2(n_58),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_142),
.B1(n_58),
.B2(n_81),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_161),
.C(n_61),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_152),
.A3(n_76),
.B1(n_52),
.B2(n_24),
.C1(n_81),
.C2(n_6),
.Y(n_161)
);

OAI21x1_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_22),
.B(n_24),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_22),
.Y(n_164)
);


endmodule