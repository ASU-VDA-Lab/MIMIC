module fake_jpeg_10776_n_583 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_583);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_583;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_59),
.B(n_60),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_63),
.B(n_66),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_67),
.B(n_87),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_68),
.B(n_70),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_71),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_72),
.Y(n_171)
);

NAND2x1_ASAP7_75t_L g73 ( 
.A(n_27),
.B(n_38),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_73),
.A2(n_7),
.B(n_9),
.Y(n_215)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_75),
.Y(n_192)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_76),
.Y(n_191)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_78),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_80),
.Y(n_178)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_81),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_103),
.Y(n_132)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_58),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g197 ( 
.A(n_85),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_21),
.B(n_0),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_86),
.B(n_90),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_0),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_89),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_1),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_28),
.B(n_1),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_99),
.B(n_117),
.Y(n_181)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_101),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_28),
.B(n_2),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_44),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_106),
.A2(n_56),
.B1(n_55),
.B2(n_42),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_110),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_111),
.Y(n_198)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_30),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_118),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_119),
.B(n_121),
.Y(n_203)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

BUFx16f_ASAP7_75t_L g121 ( 
.A(n_33),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_30),
.B(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_125),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_124),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_31),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_31),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_126),
.B(n_127),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_32),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_34),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_50),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_85),
.A2(n_35),
.B1(n_46),
.B2(n_40),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_133),
.A2(n_153),
.B1(n_157),
.B2(n_159),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_76),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_134),
.B(n_138),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_141),
.B(n_143),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_50),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_74),
.A2(n_33),
.B1(n_35),
.B2(n_40),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_145),
.A2(n_167),
.B1(n_187),
.B2(n_188),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_35),
.B1(n_46),
.B2(n_40),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g283 ( 
.A1(n_146),
.A2(n_177),
.B(n_179),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_65),
.A2(n_35),
.B1(n_46),
.B2(n_40),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_88),
.B(n_34),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_154),
.B(n_155),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_73),
.B(n_37),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_77),
.A2(n_46),
.B1(n_57),
.B2(n_47),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_84),
.A2(n_57),
.B1(n_47),
.B2(n_52),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_94),
.A2(n_57),
.B1(n_47),
.B2(n_52),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_163),
.A2(n_193),
.B1(n_15),
.B2(n_17),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_164),
.A2(n_165),
.B1(n_104),
.B2(n_15),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_106),
.A2(n_116),
.B1(n_123),
.B2(n_72),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_112),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_61),
.B(n_56),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_168),
.B(n_174),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_81),
.B(n_89),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_53),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_176),
.B(n_186),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_118),
.A2(n_54),
.B1(n_53),
.B2(n_48),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_110),
.A2(n_96),
.B1(n_54),
.B2(n_48),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_43),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_62),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_64),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_94),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_80),
.B(n_6),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_199),
.B(n_191),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_121),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_121),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_91),
.Y(n_208)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_69),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_212)
);

AO22x1_ASAP7_75t_SL g226 ( 
.A1(n_212),
.A2(n_217),
.B1(n_188),
.B2(n_215),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_71),
.A2(n_82),
.B1(n_111),
.B2(n_107),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_217),
.B1(n_93),
.B2(n_102),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_215),
.B(n_174),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_75),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_132),
.B(n_98),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_218),
.B(n_224),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_219),
.Y(n_292)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_140),
.Y(n_220)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_220),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_221),
.A2(n_240),
.B1(n_194),
.B2(n_166),
.Y(n_313)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_160),
.Y(n_225)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_225),
.Y(n_327)
);

OA22x2_ASAP7_75t_L g319 ( 
.A1(n_226),
.A2(n_228),
.B1(n_149),
.B2(n_169),
.Y(n_319)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_227),
.Y(n_300)
);

AO22x2_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_79),
.B1(n_101),
.B2(n_97),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g229 ( 
.A(n_197),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_229),
.B(n_264),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_137),
.Y(n_231)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_231),
.Y(n_295)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_232),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_168),
.B(n_95),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_235),
.A2(n_239),
.B(n_264),
.Y(n_340)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_236),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_148),
.B(n_119),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_177),
.A2(n_104),
.B1(n_119),
.B2(n_14),
.Y(n_240)
);

NAND2x1_ASAP7_75t_SL g242 ( 
.A(n_174),
.B(n_11),
.Y(n_242)
);

NAND2x1_ASAP7_75t_SL g318 ( 
.A(n_242),
.B(n_277),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_162),
.B(n_12),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_243),
.B(n_245),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_244),
.A2(n_195),
.B1(n_196),
.B2(n_171),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_135),
.B(n_14),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_246),
.Y(n_339)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_161),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_248),
.B(n_252),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_SL g249 ( 
.A1(n_212),
.A2(n_15),
.B(n_17),
.C(n_18),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_249),
.A2(n_192),
.B(n_200),
.C(n_239),
.Y(n_329)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_250),
.Y(n_334)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_136),
.Y(n_251)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_170),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_203),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_253),
.B(n_262),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_140),
.Y(n_256)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_139),
.A2(n_183),
.B1(n_206),
.B2(n_173),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_147),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_129),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_158),
.Y(n_263)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_211),
.B(n_181),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_265),
.B(n_266),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_174),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_129),
.Y(n_267)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_152),
.Y(n_269)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_130),
.Y(n_270)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_270),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_182),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_271),
.A2(n_273),
.B1(n_275),
.B2(n_278),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_187),
.B(n_175),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_274),
.Y(n_307)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_150),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_139),
.A2(n_156),
.B1(n_210),
.B2(n_180),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_209),
.B(n_144),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_276),
.Y(n_335)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_147),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_151),
.B(n_178),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_193),
.C(n_159),
.Y(n_303)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_190),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_280),
.Y(n_338)
);

INVx4_ASAP7_75t_SL g281 ( 
.A(n_151),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_281),
.A2(n_282),
.B1(n_285),
.B2(n_288),
.Y(n_316)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_178),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_167),
.B(n_180),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_284),
.A2(n_163),
.B1(n_133),
.B2(n_157),
.Y(n_294)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_172),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_198),
.B(n_145),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_289),
.Y(n_315)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_184),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_179),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_184),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_290),
.A2(n_189),
.B1(n_196),
.B2(n_195),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_182),
.B(n_131),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_291),
.B(n_171),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_294),
.A2(n_299),
.B1(n_319),
.B2(n_323),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_244),
.A2(n_214),
.B1(n_146),
.B2(n_153),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_303),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_131),
.B1(n_194),
.B2(n_166),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_304),
.A2(n_313),
.B1(n_346),
.B2(n_246),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_264),
.A2(n_189),
.B(n_184),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_320),
.A2(n_231),
.B(n_281),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_322),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_238),
.B(n_149),
.C(n_169),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_279),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_329),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_239),
.B(n_192),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_336),
.A2(n_271),
.B(n_290),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_255),
.B(n_200),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_245),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_341),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_235),
.A2(n_272),
.B(n_284),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_286),
.A2(n_283),
.B1(n_221),
.B2(n_228),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_309),
.Y(n_348)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_346),
.A2(n_230),
.B1(n_226),
.B2(n_228),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_349),
.A2(n_354),
.B1(n_366),
.B2(n_375),
.Y(n_405)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_309),
.Y(n_350)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_352),
.B(n_359),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_344),
.B(n_234),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_359),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_315),
.A2(n_319),
.B1(n_313),
.B2(n_307),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_241),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_357),
.Y(n_392)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_301),
.B(n_243),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_299),
.A2(n_228),
.B1(n_283),
.B2(n_279),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_382),
.B1(n_384),
.B2(n_314),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_300),
.Y(n_365)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_315),
.A2(n_226),
.B1(n_249),
.B2(n_242),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_334),
.Y(n_367)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_296),
.B(n_251),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_L g407 ( 
.A1(n_368),
.A2(n_377),
.B(n_385),
.Y(n_407)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_302),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_372),
.Y(n_402)
);

BUFx24_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_371),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_222),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_373),
.A2(n_378),
.B(n_381),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_312),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_379),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_319),
.A2(n_269),
.B1(n_227),
.B2(n_247),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_319),
.A2(n_232),
.B1(n_270),
.B2(n_257),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_376),
.A2(n_386),
.B1(n_389),
.B2(n_351),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_296),
.B(n_250),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_307),
.A2(n_229),
.B(n_263),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_333),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_302),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_380),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_336),
.A2(n_220),
.B1(n_268),
.B2(n_256),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_336),
.A2(n_236),
.B1(n_273),
.B2(n_278),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_233),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_318),
.Y(n_416)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_388),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_329),
.A2(n_261),
.B1(n_267),
.B2(n_303),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_390),
.A2(n_345),
.B1(n_342),
.B2(n_300),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_362),
.A2(n_310),
.B1(n_321),
.B2(n_328),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_394),
.A2(n_406),
.B1(n_409),
.B2(n_410),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_395),
.A2(n_371),
.B(n_342),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_330),
.C(n_340),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_399),
.B(n_412),
.C(n_421),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_362),
.A2(n_358),
.B1(n_349),
.B2(n_369),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_358),
.A2(n_310),
.B1(n_321),
.B2(n_320),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_387),
.A2(n_325),
.B1(n_305),
.B2(n_336),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_411),
.A2(n_418),
.B1(n_419),
.B2(n_422),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_369),
.B(n_330),
.C(n_305),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_416),
.B(n_371),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_368),
.A2(n_341),
.B1(n_292),
.B2(n_318),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_369),
.A2(n_330),
.B1(n_316),
.B2(n_345),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_420),
.A2(n_382),
.B1(n_384),
.B2(n_381),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_352),
.B(n_324),
.C(n_327),
.Y(n_421)
);

OAI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_354),
.A2(n_347),
.B1(n_297),
.B2(n_308),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_377),
.A2(n_338),
.B1(n_347),
.B2(n_311),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_361),
.B1(n_388),
.B2(n_385),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_351),
.A2(n_389),
.B(n_373),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_424),
.A2(n_298),
.B(n_326),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_425),
.B(n_367),
.C(n_363),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_405),
.A2(n_386),
.B1(n_375),
.B2(n_376),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_426),
.A2(n_427),
.B1(n_418),
.B2(n_411),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_404),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_431),
.Y(n_484)
);

OAI21xp33_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_374),
.B(n_378),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_438),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_357),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_443),
.C(n_447),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_424),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_403),
.A2(n_366),
.B(n_355),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_432),
.A2(n_440),
.B(n_449),
.Y(n_473)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_400),
.Y(n_433)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_400),
.Y(n_434)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_434),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_392),
.B(n_353),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_435),
.B(n_398),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_403),
.A2(n_356),
.B(n_360),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g441 ( 
.A1(n_394),
.A2(n_372),
.B1(n_348),
.B2(n_350),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_441),
.Y(n_482)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_311),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_416),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_406),
.A2(n_410),
.B1(n_422),
.B2(n_409),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_445),
.A2(n_405),
.B1(n_393),
.B2(n_407),
.Y(n_466)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_401),
.Y(n_446)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_419),
.A2(n_379),
.B(n_371),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_414),
.Y(n_450)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_404),
.B(n_326),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_451),
.B(n_454),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_452),
.A2(n_420),
.B(n_396),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_399),
.B(n_317),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_402),
.C(n_413),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_421),
.B(n_298),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_391),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_455),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_393),
.B(n_402),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_380),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_423),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_457),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_461),
.A2(n_471),
.B1(n_445),
.B2(n_436),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_463),
.A2(n_449),
.B(n_438),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_459),
.Y(n_499)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_431),
.A2(n_396),
.B1(n_414),
.B2(n_417),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_467),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_472),
.C(n_478),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_428),
.A2(n_417),
.B1(n_413),
.B2(n_391),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_439),
.B(n_397),
.C(n_408),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_474),
.B(n_479),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_408),
.C(n_397),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_452),
.A2(n_395),
.B(n_398),
.Y(n_479)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_481),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_297),
.Y(n_483)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_483),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_436),
.A2(n_415),
.B1(n_365),
.B2(n_308),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_426),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_447),
.Y(n_486)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_486),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_489),
.A2(n_473),
.B(n_469),
.Y(n_517)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_492),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_453),
.C(n_443),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_501),
.C(n_504),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_494),
.A2(n_507),
.B1(n_508),
.B2(n_475),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_430),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_503),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_432),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_499),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_457),
.Y(n_498)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_498),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_465),
.B(n_444),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_470),
.B(n_442),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_437),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_440),
.C(n_461),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_509),
.C(n_510),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_R g506 ( 
.A(n_469),
.B(n_437),
.C(n_433),
.Y(n_506)
);

OAI322xp33_ASAP7_75t_L g528 ( 
.A1(n_506),
.A2(n_390),
.A3(n_331),
.B1(n_293),
.B2(n_343),
.C1(n_267),
.C2(n_261),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_464),
.A2(n_455),
.B1(n_448),
.B2(n_446),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_464),
.A2(n_434),
.B1(n_450),
.B2(n_415),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_331),
.C(n_370),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_466),
.B(n_339),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_500),
.A2(n_470),
.B1(n_482),
.B2(n_473),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_511),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_516),
.A2(n_523),
.B1(n_527),
.B2(n_492),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_517),
.A2(n_528),
.B(n_508),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_469),
.C(n_463),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_521),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_487),
.B(n_462),
.C(n_479),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_490),
.B(n_475),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_524),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_494),
.A2(n_482),
.B1(n_485),
.B2(n_481),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_503),
.B(n_480),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_488),
.A2(n_477),
.B1(n_476),
.B2(n_460),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_525),
.B(n_498),
.Y(n_530)
);

AO221x1_ASAP7_75t_L g526 ( 
.A1(n_489),
.A2(n_476),
.B1(n_477),
.B2(n_460),
.C(n_458),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_526),
.A2(n_509),
.B(n_505),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_500),
.A2(n_458),
.B1(n_480),
.B2(n_365),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_529),
.A2(n_534),
.B1(n_512),
.B2(n_513),
.Y(n_544)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_530),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_521),
.A2(n_502),
.B(n_495),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_533),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_491),
.Y(n_533)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_535),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_520),
.B(n_504),
.C(n_499),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_537),
.B(n_538),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_497),
.C(n_493),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_539),
.B(n_518),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_488),
.C(n_501),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_540),
.B(n_541),
.C(n_542),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_510),
.C(n_507),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_514),
.B(n_506),
.C(n_293),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_517),
.A2(n_513),
.B(n_511),
.Y(n_543)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_543),
.Y(n_553)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_544),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_541),
.B(n_515),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_545),
.B(n_540),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_547),
.B(n_548),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_519),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_532),
.B(n_522),
.Y(n_550)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_550),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_542),
.B(n_515),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_554),
.B(n_534),
.Y(n_561)
);

NOR3xp33_ASAP7_75t_L g556 ( 
.A(n_546),
.B(n_539),
.C(n_538),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_556),
.B(n_557),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_555),
.B(n_537),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_560),
.B(n_565),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_561),
.B(n_563),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_532),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_550),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_564),
.B(n_558),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_552),
.B(n_543),
.Y(n_565)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_568),
.Y(n_576)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_564),
.A2(n_524),
.B(n_553),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_569),
.A2(n_571),
.B(n_551),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_559),
.B(n_545),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_562),
.B(n_551),
.C(n_547),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_572),
.B(n_544),
.C(n_529),
.Y(n_574)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_573),
.Y(n_578)
);

AOI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_574),
.A2(n_575),
.B(n_570),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_567),
.Y(n_575)
);

OAI321xp33_ASAP7_75t_L g580 ( 
.A1(n_577),
.A2(n_512),
.A3(n_569),
.B1(n_526),
.B2(n_528),
.C(n_527),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_566),
.C(n_576),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_579),
.B(n_580),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_516),
.B(n_523),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_582),
.B(n_525),
.Y(n_583)
);


endmodule