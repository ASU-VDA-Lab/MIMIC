module real_jpeg_29451_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_0),
.A2(n_24),
.B1(n_26),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_4),
.A2(n_9),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_4),
.A2(n_30),
.B1(n_67),
.B2(n_68),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_4),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_52)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_9),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_8),
.A2(n_24),
.B1(n_26),
.B2(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_33),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_8),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_9),
.B(n_72),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_70),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_10),
.B(n_24),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_8),
.A2(n_38),
.B(n_42),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_8),
.B(n_23),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_9),
.A2(n_10),
.B1(n_25),
.B2(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_9),
.A2(n_28),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_33),
.B(n_157),
.C(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_10),
.Y(n_157)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_11),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_117),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_116),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_90),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_90),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_76),
.B2(n_89),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_49),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_35),
.B(n_48),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_20),
.A2(n_83),
.B1(n_94),
.B2(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_20),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_20),
.B(n_147),
.C(n_148),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_20),
.A2(n_123),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_22),
.B(n_23),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_24),
.A2(n_33),
.B(n_39),
.C(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_29),
.A2(n_34),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_31),
.B(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_33),
.A2(n_67),
.B(n_71),
.C(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_33),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_33),
.B(n_40),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_36),
.A2(n_40),
.B1(n_61),
.B2(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_36),
.B(n_40),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_44),
.B(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_41),
.B(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_62),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_63),
.B1(n_64),
.B2(n_75),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_58),
.B1(n_75),
.B2(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_55),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_54),
.B(n_103),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_55),
.A2(n_80),
.B1(n_104),
.B2(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_58),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_60),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_70),
.B1(n_73),
.B2(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_73),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_67),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.C(n_86),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_78),
.A2(n_81),
.B1(n_172),
.B2(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_78),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_80),
.A2(n_101),
.B(n_129),
.Y(n_147)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_81),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_81),
.A2(n_172),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_81),
.B(n_128),
.C(n_182),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_81),
.B(n_163),
.C(n_171),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_83),
.B(n_123),
.C(n_124),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_87),
.B1(n_133),
.B2(n_134),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_86),
.B(n_106),
.C(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_86),
.A2(n_87),
.B1(n_105),
.B2(n_106),
.Y(n_202)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_113),
.C(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_97),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_95),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_97),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.C(n_112),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_98),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_105),
.B1(n_106),
.B2(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_105),
.A2(n_106),
.B1(n_177),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_106),
.B(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_113),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_223),
.B(n_228),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_150),
.B(n_211),
.C(n_222),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_140),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_120),
.B(n_140),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_130),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_121),
.B(n_131),
.C(n_138),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_128),
.A2(n_145),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_128),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_128),
.B(n_195),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_137),
.B2(n_138),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_144),
.B(n_146),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_147),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_210),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_205),
.B(n_209),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_173),
.B(n_204),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_154),
.B(n_162),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_161),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_165),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_170),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_199),
.B(n_203),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_184),
.B(n_198),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_179),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_177),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_180),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_188),
.B(n_197),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_194),
.B(n_196),
.Y(n_188)
);

INVx5_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_220),
.B2(n_221),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);


endmodule