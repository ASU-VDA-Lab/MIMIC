module fake_jpeg_21558_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_39),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_59)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_42),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_57),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

A2O1A1O1Ixp25_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_18),
.B(n_27),
.C(n_14),
.D(n_23),
.Y(n_52)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_18),
.Y(n_75)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_49),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_17),
.B1(n_15),
.B2(n_22),
.Y(n_74)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_89),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_20),
.B(n_17),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_6),
.B(n_7),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_72),
.Y(n_90)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_43),
.A3(n_31),
.B1(n_41),
.B2(n_22),
.Y(n_72)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_76),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_85),
.B1(n_56),
.B2(n_62),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_R g103 ( 
.A(n_75),
.B(n_86),
.Y(n_103)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_45),
.B1(n_55),
.B2(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_18),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_95),
.B1(n_100),
.B2(n_109),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_60),
.B1(n_38),
.B2(n_5),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_27),
.C(n_23),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_19),
.C(n_70),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_2),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_105),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_19),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_3),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_63),
.B(n_6),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_68),
.A2(n_73),
.A3(n_63),
.B1(n_83),
.B2(n_87),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_114),
.B(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_64),
.B(n_82),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_9),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_105),
.B(n_12),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_71),
.B(n_88),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_88),
.C(n_67),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_120),
.C(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_67),
.C(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_84),
.B(n_7),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_84),
.C(n_76),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_91),
.C(n_103),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_135),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_91),
.B(n_109),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_95),
.B(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_128),
.C(n_134),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_134),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_146),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_110),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_144),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_122),
.B(n_111),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_130),
.Y(n_147)
);

AO21x1_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_123),
.B(n_101),
.Y(n_151)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_148),
.B(n_125),
.CI(n_137),
.CON(n_153),
.SN(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_139),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_146),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_137),
.C(n_97),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_155),
.C(n_144),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_126),
.A3(n_131),
.B1(n_100),
.B2(n_97),
.C1(n_99),
.C2(n_93),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_160),
.C(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_161),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_156),
.B(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_145),
.Y(n_162)
);

AOI31xp67_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_151),
.A3(n_154),
.B(n_153),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_165),
.A3(n_150),
.B1(n_158),
.B2(n_100),
.C1(n_147),
.C2(n_102),
.Y(n_167)
);

NOR2xp67_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_152),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_166),
.B1(n_12),
.B2(n_13),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_13),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_169),
.Y(n_172)
);


endmodule