module fake_jpeg_7004_n_264 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_264);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_27),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_40),
.C(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_26),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_23),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_23),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_41),
.B1(n_25),
.B2(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_13),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_18),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_51),
.C(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_73),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_41),
.B1(n_25),
.B2(n_40),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_69),
.B1(n_41),
.B2(n_47),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_18),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_91),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_79),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_82),
.B1(n_68),
.B2(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_75),
.B1(n_63),
.B2(n_74),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_41),
.B1(n_25),
.B2(n_45),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_61),
.B(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_90),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_93),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_60),
.Y(n_97)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_43),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_65),
.B(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_109),
.Y(n_115)
);

AOI221xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_79),
.B1(n_17),
.B2(n_22),
.C(n_24),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_106),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_68),
.B1(n_71),
.B2(n_76),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_108),
.B1(n_78),
.B2(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_67),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_71),
.B1(n_69),
.B2(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_43),
.B1(n_13),
.B2(n_18),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_77),
.B1(n_78),
.B2(n_14),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_81),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_22),
.B(n_54),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_49),
.CI(n_19),
.CON(n_128),
.SN(n_128)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_120),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_121),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_89),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_97),
.C(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_83),
.B1(n_85),
.B2(n_79),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_100),
.B1(n_98),
.B2(n_95),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_130),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_111),
.B(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_22),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_136),
.B(n_138),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_128),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_101),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_141),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_97),
.C(n_98),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_32),
.C(n_35),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_115),
.B(n_108),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_144),
.B1(n_124),
.B2(n_128),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_100),
.B1(n_95),
.B2(n_112),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_28),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_147),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_28),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_31),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_150),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_31),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_114),
.B(n_32),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_130),
.C(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_156),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_122),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_159),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_90),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_131),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_167),
.C(n_169),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_124),
.C(n_116),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_133),
.C(n_94),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_90),
.C(n_45),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_174),
.C(n_21),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_170),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_62),
.B(n_19),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_148),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_135),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_188),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_35),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_160),
.A2(n_149),
.B1(n_145),
.B2(n_64),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_62),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_193),
.B(n_178),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_58),
.C(n_38),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_192),
.C(n_58),
.Y(n_204)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_24),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_38),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_189),
.Y(n_197)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_174),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_58),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_12),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_201),
.B(n_203),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_173),
.B(n_19),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_198),
.B(n_209),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_173),
.B(n_24),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_38),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_0),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_180),
.C(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_207),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_35),
.B1(n_38),
.B2(n_10),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_38),
.C(n_35),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_21),
.C(n_20),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_15),
.B(n_20),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_206),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_197),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_207),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_210),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_206),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_217),
.C(n_220),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_183),
.B(n_10),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_223),
.B(n_224),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_9),
.C(n_12),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_199),
.B(n_9),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_221),
.A2(n_194),
.B1(n_209),
.B2(n_202),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_229),
.B(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_15),
.C(n_21),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_36),
.A3(n_21),
.B1(n_20),
.B2(n_15),
.C1(n_17),
.C2(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_36),
.Y(n_234)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_0),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_8),
.B(n_11),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_36),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_218),
.B(n_211),
.C(n_216),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_240),
.B(n_241),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_226),
.C(n_2),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_36),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_20),
.B(n_15),
.C(n_7),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_225),
.B(n_10),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_247),
.B(n_249),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_250),
.C(n_251),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_226),
.B(n_17),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_11),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_1),
.B(n_2),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_1),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_253),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_252),
.A2(n_245),
.B1(n_2),
.B2(n_4),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_6),
.Y(n_261)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_1),
.B(n_4),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_4),
.B(n_5),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_255),
.C(n_6),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_260),
.A2(n_261),
.B(n_258),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);


endmodule