module fake_ibex_1742_n_875 (n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_120, n_93, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_126, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_875);

input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_120;
input n_93;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_126;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_875;

wire n_151;
wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_153;
wire n_862;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_317;
wire n_280;
wire n_340;
wire n_375;
wire n_698;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_723;
wire n_170;
wire n_270;
wire n_383;
wire n_346;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_798;
wire n_832;
wire n_732;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_155;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_392;
wire n_354;
wire n_206;
wire n_179;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_562;
wire n_564;
wire n_506;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_820;
wire n_805;
wire n_670;
wire n_728;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_202;
wire n_298;
wire n_159;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_1),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_102),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_0),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_77),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_61),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_78),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_17),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_41),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_L g167 ( 
.A(n_58),
.B(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_35),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_L g173 ( 
.A(n_23),
.B(n_18),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_53),
.Y(n_174)
);

NOR2xp67_ASAP7_75t_L g175 ( 
.A(n_17),
.B(n_81),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_67),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_18),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_59),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_44),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_116),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_47),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_87),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_20),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_52),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_82),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_27),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_8),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_101),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_112),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_15),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_43),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_88),
.B(n_95),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_49),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_128),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_40),
.Y(n_202)
);

INVxp33_ASAP7_75t_SL g203 ( 
.A(n_122),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_28),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_45),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_16),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_38),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_79),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_66),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_21),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_99),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_19),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_135),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_127),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_48),
.B(n_100),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_29),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_103),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_110),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_132),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_138),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_54),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_33),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_19),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_39),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_108),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_133),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_105),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_20),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_70),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_134),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_28),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_15),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_14),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_14),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_84),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_29),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_62),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_124),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_34),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_34),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_68),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_25),
.B(n_139),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_94),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_71),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_163),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_162),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_228),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_0),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

AND2x6_ASAP7_75t_L g261 ( 
.A(n_165),
.B(n_42),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_200),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_163),
.Y(n_263)
);

OAI22x1_ASAP7_75t_SL g264 ( 
.A1(n_206),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_163),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_237),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_182),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_185),
.B(n_3),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_229),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_157),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_203),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_165),
.B(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_154),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_149),
.B(n_9),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_164),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_158),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_168),
.B(n_9),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_197),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_178),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_241),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_150),
.B(n_10),
.Y(n_289)
);

CKINVDCx6p67_ASAP7_75t_R g290 ( 
.A(n_191),
.Y(n_290)
);

AOI22x1_ASAP7_75t_SL g291 ( 
.A1(n_206),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_202),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_202),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_204),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_182),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_197),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_199),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_13),
.Y(n_298)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_201),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_188),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_201),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_208),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_303)
);

BUFx8_ASAP7_75t_L g304 ( 
.A(n_219),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_184),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_305)
);

OA21x2_ASAP7_75t_L g306 ( 
.A1(n_222),
.A2(n_80),
.B(n_147),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_216),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_236),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_253),
.B(n_46),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_151),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_152),
.B(n_153),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_166),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_170),
.Y(n_317)
);

CKINVDCx6p67_ASAP7_75t_R g318 ( 
.A(n_184),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_171),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_205),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_172),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_174),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_177),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_189),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_180),
.B(n_26),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_181),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_205),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_259),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_298),
.B(n_183),
.Y(n_332)
);

OR2x6_ASAP7_75t_L g333 ( 
.A(n_283),
.B(n_173),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_297),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_266),
.B(n_158),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_L g339 ( 
.A1(n_278),
.A2(n_274),
.B1(n_318),
.B2(n_322),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_298),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_266),
.B(n_213),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_297),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_256),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_317),
.B(n_187),
.Y(n_346)
);

AO22x2_ASAP7_75t_L g347 ( 
.A1(n_291),
.A2(n_250),
.B1(n_247),
.B2(n_214),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_256),
.Y(n_349)
);

AND3x2_ASAP7_75t_L g350 ( 
.A(n_275),
.B(n_325),
.C(n_300),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_266),
.B(n_159),
.Y(n_353)
);

AOI21x1_ASAP7_75t_L g354 ( 
.A1(n_306),
.A2(n_192),
.B(n_190),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_301),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_258),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_261),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_277),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_255),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_258),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_261),
.A2(n_203),
.B1(n_212),
.B2(n_225),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_262),
.B(n_245),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_268),
.B(n_194),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_258),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_261),
.A2(n_230),
.B1(n_235),
.B2(n_234),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_279),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_159),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_270),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_210),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_254),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_317),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_317),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_265),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_270),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_257),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_304),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_302),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_296),
.B(n_227),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_304),
.Y(n_384)
);

OR2x6_ASAP7_75t_L g385 ( 
.A(n_305),
.B(n_175),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_302),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g387 ( 
.A(n_267),
.B(n_304),
.C(n_319),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_285),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_302),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_285),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_295),
.A2(n_207),
.B1(n_217),
.B2(n_218),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_267),
.B(n_249),
.C(n_196),
.Y(n_392)
);

OR2x6_ASAP7_75t_L g393 ( 
.A(n_303),
.B(n_167),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_296),
.B(n_299),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_286),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_292),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_280),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_290),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_282),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_321),
.B(n_211),
.C(n_239),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_265),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_296),
.B(n_160),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_287),
.Y(n_403)
);

BUFx6f_ASAP7_75t_SL g404 ( 
.A(n_311),
.Y(n_404)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_306),
.A2(n_186),
.B(n_176),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_265),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_324),
.B(n_160),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_290),
.A2(n_289),
.B1(n_281),
.B2(n_272),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_294),
.B(n_161),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_286),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_293),
.B(n_161),
.Y(n_411)
);

NAND3xp33_ASAP7_75t_L g412 ( 
.A(n_326),
.B(n_240),
.C(n_242),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_286),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_286),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_286),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_296),
.B(n_169),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_313),
.B(n_169),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_309),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_310),
.B(n_193),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_316),
.B(n_193),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_299),
.B(n_195),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_255),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_316),
.B(n_323),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_328),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_368),
.B(n_315),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_315),
.Y(n_427)
);

NOR3xp33_ASAP7_75t_L g428 ( 
.A(n_339),
.B(n_391),
.C(n_392),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_315),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_381),
.B(n_217),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_315),
.Y(n_433)
);

AOI221xp5_ASAP7_75t_L g434 ( 
.A1(n_339),
.A2(n_307),
.B1(n_364),
.B2(n_369),
.C(n_367),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_358),
.B(n_195),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_338),
.B(n_315),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_353),
.B(n_320),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_408),
.B(n_221),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_354),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_371),
.B(n_323),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_401),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_341),
.B(n_327),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_417),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_405),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_332),
.A2(n_306),
.B(n_284),
.Y(n_446)
);

A2O1A1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_336),
.A2(n_276),
.B(n_273),
.C(n_231),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_345),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_349),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_420),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_370),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_384),
.B(n_328),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_406),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_397),
.B(n_224),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

AOI221xp5_ASAP7_75t_SL g457 ( 
.A1(n_330),
.A2(n_331),
.B1(n_335),
.B2(n_332),
.C(n_340),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_399),
.B(n_226),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_398),
.B(n_264),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_359),
.B(n_363),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_418),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_365),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_350),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_379),
.B(n_218),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_411),
.B(n_232),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_396),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_362),
.B(n_155),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_412),
.B(n_387),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_362),
.A2(n_261),
.B1(n_311),
.B2(n_299),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_400),
.B(n_156),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_366),
.B(n_402),
.Y(n_473)
);

BUFx5_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_333),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_393),
.A2(n_233),
.B1(n_223),
.B2(n_311),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_179),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_416),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_416),
.B(n_421),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_333),
.B(n_223),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_383),
.A2(n_299),
.B(n_198),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_393),
.A2(n_233),
.B1(n_385),
.B2(n_333),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_383),
.B(n_243),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_424),
.B(n_30),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_393),
.B(n_30),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_372),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_385),
.A2(n_311),
.B1(n_299),
.B2(n_314),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_394),
.Y(n_490)
);

NOR3xp33_ASAP7_75t_L g491 ( 
.A(n_346),
.B(n_347),
.C(n_238),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_404),
.A2(n_311),
.B1(n_314),
.B2(n_308),
.Y(n_492)
);

NOR3xp33_ASAP7_75t_L g493 ( 
.A(n_347),
.B(n_246),
.C(n_308),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_394),
.B(n_311),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_347),
.B(n_288),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_372),
.B(n_374),
.Y(n_496)
);

AND2x6_ASAP7_75t_SL g497 ( 
.A(n_404),
.B(n_31),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_374),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_376),
.B(n_288),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_376),
.B(n_288),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_395),
.Y(n_501)
);

INVx8_ASAP7_75t_L g502 ( 
.A(n_360),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_410),
.B(n_32),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_476),
.A2(n_413),
.B1(n_415),
.B2(n_414),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_474),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_474),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_442),
.B(n_33),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_465),
.Y(n_508)
);

BUFx12f_ASAP7_75t_L g509 ( 
.A(n_497),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_482),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_474),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_446),
.A2(n_352),
.B(n_329),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_461),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

O2A1O1Ixp33_ASAP7_75t_L g516 ( 
.A1(n_447),
.A2(n_355),
.B(n_389),
.C(n_386),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_444),
.B(n_36),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_473),
.A2(n_344),
.B(n_389),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_468),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_428),
.A2(n_434),
.B1(n_450),
.B2(n_443),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_425),
.A2(n_348),
.B(n_334),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_452),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_436),
.A2(n_355),
.B(n_337),
.Y(n_523)
);

O2A1O1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_428),
.A2(n_356),
.B(n_386),
.C(n_382),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_427),
.A2(n_356),
.B(n_342),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_430),
.B(n_343),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_429),
.A2(n_343),
.B(n_375),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_375),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_471),
.A2(n_434),
.B1(n_460),
.B2(n_440),
.Y(n_529)
);

AND2x6_ASAP7_75t_SL g530 ( 
.A(n_459),
.B(n_37),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_433),
.A2(n_480),
.B(n_494),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_481),
.A2(n_378),
.B(n_422),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_430),
.B(n_312),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_431),
.B(n_38),
.Y(n_534)
);

A2O1A1Ixp33_ASAP7_75t_L g535 ( 
.A1(n_470),
.A2(n_312),
.B(n_255),
.C(n_269),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_445),
.A2(n_439),
.B(n_466),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_437),
.B(n_50),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_430),
.Y(n_538)
);

INVx11_ASAP7_75t_L g539 ( 
.A(n_475),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

A2O1A1Ixp33_ASAP7_75t_L g541 ( 
.A1(n_457),
.A2(n_312),
.B(n_269),
.C(n_263),
.Y(n_541)
);

BUFx8_ASAP7_75t_L g542 ( 
.A(n_464),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_491),
.B(n_269),
.Y(n_543)
);

INVx6_ASAP7_75t_L g544 ( 
.A(n_487),
.Y(n_544)
);

O2A1O1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_438),
.A2(n_55),
.B(n_57),
.C(n_60),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_455),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_439),
.A2(n_490),
.B(n_469),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_502),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_454),
.B(n_458),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_493),
.A2(n_263),
.B1(n_260),
.B2(n_360),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_467),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_449),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_493),
.B(n_63),
.C(n_64),
.Y(n_554)
);

OR2x6_ASAP7_75t_SL g555 ( 
.A(n_486),
.B(n_459),
.Y(n_555)
);

A2O1A1Ixp33_ASAP7_75t_L g556 ( 
.A1(n_456),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_556)
);

AO32x2_ASAP7_75t_L g557 ( 
.A1(n_483),
.A2(n_489),
.A3(n_495),
.B1(n_492),
.B2(n_463),
.Y(n_557)
);

BUFx8_ASAP7_75t_SL g558 ( 
.A(n_459),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_477),
.B(n_479),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_462),
.Y(n_560)
);

NAND2x1p5_ASAP7_75t_L g561 ( 
.A(n_432),
.B(n_426),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_478),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_472),
.B(n_92),
.Y(n_563)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_435),
.A2(n_93),
.B(n_96),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_502),
.Y(n_565)
);

A2O1A1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_485),
.A2(n_107),
.B(n_109),
.C(n_111),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_441),
.Y(n_567)
);

OAI21xp33_ASAP7_75t_L g568 ( 
.A1(n_492),
.A2(n_114),
.B(n_115),
.Y(n_568)
);

A2O1A1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_453),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_L g570 ( 
.A(n_499),
.B(n_500),
.Y(n_570)
);

AO21x1_ASAP7_75t_L g571 ( 
.A1(n_501),
.A2(n_496),
.B(n_488),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_502),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_544),
.B(n_498),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_542),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_513),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_558),
.B(n_542),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_536),
.A2(n_550),
.B(n_531),
.Y(n_577)
);

AO31x2_ASAP7_75t_L g578 ( 
.A1(n_541),
.A2(n_571),
.A3(n_535),
.B(n_566),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_572),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_520),
.B(n_519),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_517),
.A2(n_520),
.B(n_534),
.Y(n_581)
);

AO31x2_ASAP7_75t_L g582 ( 
.A1(n_548),
.A2(n_556),
.A3(n_512),
.B(n_569),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_524),
.A2(n_537),
.B(n_516),
.C(n_507),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_508),
.B(n_522),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_510),
.A2(n_544),
.B1(n_543),
.B2(n_540),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_553),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_521),
.A2(n_527),
.B(n_525),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_559),
.A2(n_505),
.B1(n_552),
.B2(n_563),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_560),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_509),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_547),
.B(n_528),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_539),
.Y(n_593)
);

CKINVDCx9p33_ASAP7_75t_R g594 ( 
.A(n_555),
.Y(n_594)
);

AO32x2_ASAP7_75t_L g595 ( 
.A1(n_504),
.A2(n_562),
.A3(n_543),
.B1(n_554),
.B2(n_551),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_567),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_565),
.B(n_561),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_523),
.A2(n_564),
.B(n_532),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_549),
.B(n_561),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_506),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_570),
.B(n_557),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_511),
.B(n_515),
.Y(n_603)
);

NAND3xp33_ASAP7_75t_SL g604 ( 
.A(n_554),
.B(n_545),
.C(n_568),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_538),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_518),
.Y(n_606)
);

AO31x2_ASAP7_75t_L g607 ( 
.A1(n_557),
.A2(n_533),
.A3(n_526),
.B(n_530),
.Y(n_607)
);

INVx3_ASAP7_75t_SL g608 ( 
.A(n_530),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_542),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_514),
.B(n_519),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_505),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_514),
.A2(n_520),
.B1(n_540),
.B2(n_529),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_549),
.B(n_451),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_513),
.A2(n_271),
.B1(n_328),
.B2(n_451),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_544),
.B(n_451),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_514),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_513),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_565),
.B(n_451),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_517),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_514),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_514),
.B(n_520),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_514),
.Y(n_622)
);

NOR2x1_ASAP7_75t_L g623 ( 
.A(n_565),
.B(n_451),
.Y(n_623)
);

AO31x2_ASAP7_75t_L g624 ( 
.A1(n_541),
.A2(n_571),
.A3(n_535),
.B(n_536),
.Y(n_624)
);

AO31x2_ASAP7_75t_L g625 ( 
.A1(n_541),
.A2(n_571),
.A3(n_535),
.B(n_536),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g626 ( 
.A1(n_514),
.A2(n_520),
.B1(n_540),
.B2(n_529),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_544),
.B(n_451),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_544),
.B(n_451),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_514),
.A2(n_520),
.B1(n_540),
.B2(n_529),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_513),
.A2(n_271),
.B1(n_328),
.B2(n_451),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_517),
.A2(n_391),
.B(n_451),
.Y(n_631)
);

AO22x2_ASAP7_75t_L g632 ( 
.A1(n_517),
.A2(n_484),
.B1(n_493),
.B2(n_491),
.Y(n_632)
);

CKINVDCx11_ASAP7_75t_R g633 ( 
.A(n_509),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_514),
.Y(n_634)
);

AO31x2_ASAP7_75t_L g635 ( 
.A1(n_541),
.A2(n_571),
.A3(n_535),
.B(n_536),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_514),
.B(n_520),
.Y(n_636)
);

CKINVDCx11_ASAP7_75t_R g637 ( 
.A(n_509),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_514),
.B(n_520),
.Y(n_638)
);

AO31x2_ASAP7_75t_L g639 ( 
.A1(n_541),
.A2(n_571),
.A3(n_535),
.B(n_536),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_513),
.B(n_442),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_513),
.B(n_451),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_514),
.A2(n_520),
.B1(n_540),
.B2(n_529),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_514),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_513),
.B(n_442),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_514),
.B(n_520),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_513),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_531),
.A2(n_446),
.B(n_541),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_514),
.Y(n_650)
);

NAND2x1p5_ASAP7_75t_L g651 ( 
.A(n_565),
.B(n_451),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_531),
.A2(n_446),
.B(n_541),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_544),
.B(n_451),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_544),
.B(n_451),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_649),
.A2(n_652),
.B(n_598),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_612),
.A2(n_642),
.B1(n_629),
.B2(n_626),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_634),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_640),
.B(n_646),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_616),
.Y(n_659)
);

OAI21x1_ASAP7_75t_L g660 ( 
.A1(n_606),
.A2(n_577),
.B(n_588),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_644),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_620),
.B(n_622),
.Y(n_662)
);

NAND2x1p5_ASAP7_75t_L g663 ( 
.A(n_645),
.B(n_643),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_618),
.Y(n_664)
);

OAI21x1_ASAP7_75t_SL g665 ( 
.A1(n_581),
.A2(n_589),
.B(n_580),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_651),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_645),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_641),
.B(n_648),
.Y(n_668)
);

BUFx12f_ASAP7_75t_L g669 ( 
.A(n_633),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_620),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_574),
.Y(n_671)
);

AO21x2_ASAP7_75t_L g672 ( 
.A1(n_604),
.A2(n_583),
.B(n_602),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_645),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_622),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_650),
.Y(n_675)
);

OA21x2_ASAP7_75t_L g676 ( 
.A1(n_636),
.A2(n_638),
.B(n_647),
.Y(n_676)
);

BUFx8_ASAP7_75t_L g677 ( 
.A(n_609),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_632),
.A2(n_610),
.B1(n_585),
.B2(n_608),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_590),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_584),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_610),
.B(n_617),
.Y(n_681)
);

AO31x2_ASAP7_75t_L g682 ( 
.A1(n_596),
.A2(n_587),
.A3(n_601),
.B(n_639),
.Y(n_682)
);

AO21x2_ASAP7_75t_L g683 ( 
.A1(n_595),
.A2(n_601),
.B(n_639),
.Y(n_683)
);

AO31x2_ASAP7_75t_L g684 ( 
.A1(n_624),
.A2(n_625),
.A3(n_635),
.B(n_639),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_632),
.B(n_631),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g686 ( 
.A1(n_592),
.A2(n_605),
.B(n_586),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_599),
.A2(n_603),
.B(n_600),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_575),
.B(n_627),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_615),
.B(n_628),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_597),
.B(n_611),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_653),
.B(n_654),
.Y(n_691)
);

BUFx4f_ASAP7_75t_SL g692 ( 
.A(n_579),
.Y(n_692)
);

NAND2x1p5_ASAP7_75t_L g693 ( 
.A(n_623),
.B(n_613),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_614),
.B(n_630),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_625),
.A2(n_582),
.B(n_578),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_594),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_607),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_573),
.A2(n_607),
.B(n_619),
.Y(n_698)
);

NAND2x1_ASAP7_75t_L g699 ( 
.A(n_593),
.B(n_576),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_591),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_637),
.B(n_641),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_634),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_620),
.B(n_622),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_634),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_L g705 ( 
.A(n_645),
.B(n_641),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_634),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_634),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_634),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_620),
.B(n_622),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_645),
.Y(n_710)
);

AO21x1_ASAP7_75t_L g711 ( 
.A1(n_589),
.A2(n_543),
.B(n_581),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_634),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_634),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_621),
.B(n_520),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_633),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_634),
.Y(n_716)
);

AND3x4_ASAP7_75t_L g717 ( 
.A(n_574),
.B(n_493),
.C(n_428),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_682),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_694),
.B(n_701),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_675),
.B(n_682),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_682),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_668),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_670),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_705),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_674),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_662),
.B(n_703),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_664),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_685),
.B(n_714),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_677),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_710),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_710),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_696),
.A2(n_665),
.B1(n_692),
.B2(n_709),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_679),
.B(n_658),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_717),
.A2(n_691),
.B1(n_689),
.B2(n_656),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_692),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_676),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_659),
.B(n_676),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_666),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_680),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_657),
.B(n_712),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_661),
.B(n_707),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_717),
.A2(n_678),
.B1(n_711),
.B2(n_681),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_702),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_704),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_690),
.B(n_713),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_706),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_678),
.B(n_688),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_708),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_716),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_663),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_667),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_667),
.Y(n_753)
);

OR2x6_ASAP7_75t_L g754 ( 
.A(n_698),
.B(n_687),
.Y(n_754)
);

OA21x2_ASAP7_75t_L g755 ( 
.A1(n_655),
.A2(n_695),
.B(n_660),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_663),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_720),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_738),
.B(n_683),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_754),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_738),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_720),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_754),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_718),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_729),
.B(n_684),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_737),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_727),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_737),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_719),
.A2(n_690),
.B1(n_697),
.B2(n_672),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_721),
.B(n_684),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_SL g770 ( 
.A(n_725),
.B(n_677),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_729),
.B(n_684),
.Y(n_771)
);

NOR4xp25_ASAP7_75t_SL g772 ( 
.A(n_730),
.B(n_715),
.C(n_700),
.D(n_669),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_723),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_769),
.B(n_724),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_763),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_760),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_769),
.B(n_764),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_763),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_773),
.B(n_733),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_763),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_765),
.Y(n_781)
);

AND2x4_ASAP7_75t_SL g782 ( 
.A(n_760),
.B(n_754),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_773),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_758),
.B(n_755),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_760),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_758),
.B(n_755),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_765),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_769),
.B(n_726),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_773),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_757),
.B(n_762),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_764),
.B(n_726),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_767),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_767),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_775),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_777),
.B(n_764),
.Y(n_795)
);

NAND4xp25_ASAP7_75t_L g796 ( 
.A(n_791),
.B(n_743),
.C(n_770),
.D(n_735),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_792),
.B(n_730),
.Y(n_797)
);

OAI332xp33_ASAP7_75t_L g798 ( 
.A1(n_791),
.A2(n_770),
.A3(n_748),
.B1(n_734),
.B2(n_771),
.B3(n_736),
.C1(n_788),
.C2(n_774),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_775),
.Y(n_799)
);

NAND2x1_ASAP7_75t_L g800 ( 
.A(n_776),
.B(n_759),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_774),
.B(n_771),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_778),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_784),
.B(n_757),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_784),
.B(n_757),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_780),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_784),
.B(n_761),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_788),
.B(n_771),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_789),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_776),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_777),
.B(n_761),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_796),
.B(n_669),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_798),
.B(n_722),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_803),
.B(n_786),
.Y(n_813)
);

NAND2x1_ASAP7_75t_L g814 ( 
.A(n_797),
.B(n_776),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_810),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_810),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_794),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_794),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_800),
.A2(n_779),
.B(n_787),
.Y(n_819)
);

OAI21xp33_ASAP7_75t_SL g820 ( 
.A1(n_809),
.A2(n_779),
.B(n_787),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_808),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_803),
.B(n_785),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_795),
.B(n_781),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_799),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_814),
.Y(n_825)
);

OAI32xp33_ASAP7_75t_L g826 ( 
.A1(n_820),
.A2(n_808),
.A3(n_795),
.B1(n_783),
.B2(n_789),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_821),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_815),
.B(n_804),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_816),
.B(n_804),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_812),
.A2(n_806),
.B1(n_807),
.B2(n_801),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_811),
.A2(n_806),
.B1(n_786),
.B2(n_790),
.Y(n_831)
);

AO22x1_ASAP7_75t_L g832 ( 
.A1(n_821),
.A2(n_715),
.B1(n_677),
.B2(n_785),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_819),
.A2(n_800),
.B(n_786),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_823),
.B(n_799),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_813),
.B(n_805),
.Y(n_835)
);

OAI221xp5_ASAP7_75t_L g836 ( 
.A1(n_833),
.A2(n_819),
.B1(n_768),
.B2(n_824),
.C(n_818),
.Y(n_836)
);

AOI221xp5_ASAP7_75t_L g837 ( 
.A1(n_826),
.A2(n_822),
.B1(n_817),
.B2(n_768),
.C(n_802),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_SL g838 ( 
.A1(n_825),
.A2(n_785),
.B1(n_792),
.B2(n_783),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_834),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_827),
.A2(n_782),
.B(n_783),
.C(n_789),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_SL g841 ( 
.A1(n_832),
.A2(n_699),
.B(n_793),
.C(n_781),
.Y(n_841)
);

OAI221xp5_ASAP7_75t_SL g842 ( 
.A1(n_837),
.A2(n_831),
.B1(n_830),
.B2(n_748),
.C(n_829),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_839),
.B(n_836),
.Y(n_843)
);

NAND4xp25_ASAP7_75t_L g844 ( 
.A(n_841),
.B(n_783),
.C(n_739),
.D(n_759),
.Y(n_844)
);

NOR2x1_ASAP7_75t_L g845 ( 
.A(n_844),
.B(n_840),
.Y(n_845)
);

NOR3xp33_ASAP7_75t_L g846 ( 
.A(n_843),
.B(n_838),
.C(n_671),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_L g847 ( 
.A(n_845),
.B(n_846),
.C(n_842),
.Y(n_847)
);

AND3x4_ASAP7_75t_L g848 ( 
.A(n_845),
.B(n_772),
.C(n_766),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_R g849 ( 
.A(n_848),
.B(n_772),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_847),
.Y(n_850)
);

AND4x1_ASAP7_75t_L g851 ( 
.A(n_850),
.B(n_828),
.C(n_835),
.D(n_686),
.Y(n_851)
);

NOR2x1_ASAP7_75t_L g852 ( 
.A(n_849),
.B(n_731),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_852),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_851),
.A2(n_728),
.B1(n_732),
.B2(n_746),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_852),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_853),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_855),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_854),
.B(n_731),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_855),
.A2(n_693),
.B(n_732),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_855),
.A2(n_693),
.B(n_741),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_856),
.A2(n_734),
.B1(n_753),
.B2(n_752),
.Y(n_861)
);

AOI22x1_ASAP7_75t_SL g862 ( 
.A1(n_857),
.A2(n_740),
.B1(n_750),
.B2(n_749),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_SL g863 ( 
.A1(n_859),
.A2(n_742),
.B(n_740),
.C(n_747),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_858),
.B(n_860),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_858),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_856),
.A2(n_745),
.B(n_750),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_857),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_867),
.A2(n_745),
.B(n_744),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_865),
.A2(n_756),
.B1(n_751),
.B2(n_723),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_864),
.Y(n_870)
);

AOI21xp33_ASAP7_75t_L g871 ( 
.A1(n_861),
.A2(n_747),
.B(n_744),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_870),
.B(n_866),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_868),
.B(n_862),
.C(n_863),
.Y(n_873)
);

AO21x2_ASAP7_75t_L g874 ( 
.A1(n_872),
.A2(n_869),
.B(n_871),
.Y(n_874)
);

AOI21xp33_ASAP7_75t_SL g875 ( 
.A1(n_874),
.A2(n_873),
.B(n_749),
.Y(n_875)
);


endmodule