module fake_netlist_5_2232_n_22012 (n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_22012);

input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_22012;

wire n_924;
wire n_19133;
wire n_977;
wire n_9936;
wire n_4706;
wire n_20081;
wire n_14870;
wire n_2380;
wire n_15741;
wire n_3006;
wire n_532;
wire n_10794;
wire n_5287;
wire n_12872;
wire n_15349;
wire n_11207;
wire n_19036;
wire n_8174;
wire n_5161;
wire n_15269;
wire n_20874;
wire n_5776;
wire n_6551;
wire n_10793;
wire n_10552;
wire n_12215;
wire n_4963;
wire n_20753;
wire n_19588;
wire n_19261;
wire n_5282;
wire n_11349;
wire n_8328;
wire n_8060;
wire n_14939;
wire n_21305;
wire n_3813;
wire n_15935;
wire n_10108;
wire n_7660;
wire n_671;
wire n_18799;
wire n_3445;
wire n_18722;
wire n_8617;
wire n_3785;
wire n_17921;
wire n_10117;
wire n_12139;
wire n_14762;
wire n_21716;
wire n_7205;
wire n_3019;
wire n_17714;
wire n_8319;
wire n_6694;
wire n_4517;
wire n_15406;
wire n_4425;
wire n_14287;
wire n_1860;
wire n_17679;
wire n_19837;
wire n_14471;
wire n_20126;
wire n_6913;
wire n_10756;
wire n_19801;
wire n_11653;
wire n_8961;
wire n_16240;
wire n_7772;
wire n_5402;
wire n_17017;
wire n_13889;
wire n_5509;
wire n_9773;
wire n_11089;
wire n_14045;
wire n_18391;
wire n_16498;
wire n_12709;
wire n_9173;
wire n_18413;
wire n_16910;
wire n_11296;
wire n_8681;
wire n_9796;
wire n_519;
wire n_5469;
wire n_6431;
wire n_12266;
wire n_9049;
wire n_11917;
wire n_7861;
wire n_9907;
wire n_5202;
wire n_14898;
wire n_16663;
wire n_9539;
wire n_14270;
wire n_569;
wire n_10421;
wire n_7523;
wire n_16256;
wire n_21022;
wire n_3631;
wire n_16182;
wire n_14959;
wire n_21785;
wire n_1566;
wire n_297;
wire n_9500;
wire n_16017;
wire n_16295;
wire n_6085;
wire n_7306;
wire n_8819;
wire n_223;
wire n_7493;
wire n_12027;
wire n_3868;
wire n_12111;
wire n_12075;
wire n_264;
wire n_21149;
wire n_3687;
wire n_13708;
wire n_21487;
wire n_5241;
wire n_6939;
wire n_882;
wire n_2384;
wire n_7528;
wire n_14519;
wire n_3156;
wire n_9206;
wire n_646;
wire n_14611;
wire n_12142;
wire n_2202;
wire n_16764;
wire n_11354;
wire n_19720;
wire n_13782;
wire n_8310;
wire n_19369;
wire n_11052;
wire n_15548;
wire n_17791;
wire n_6920;
wire n_18260;
wire n_17685;
wire n_21153;
wire n_1561;
wire n_16514;
wire n_3361;
wire n_1600;
wire n_9040;
wire n_19849;
wire n_14336;
wire n_15813;
wire n_10626;
wire n_4255;
wire n_1796;
wire n_901;
wire n_18414;
wire n_7152;
wire n_16452;
wire n_18812;
wire n_18998;
wire n_13571;
wire n_4237;
wire n_1672;
wire n_19848;
wire n_20234;
wire n_637;
wire n_8126;
wire n_17635;
wire n_18274;
wire n_5894;
wire n_19570;
wire n_2079;
wire n_7801;
wire n_11588;
wire n_11689;
wire n_10231;
wire n_7463;
wire n_20038;
wire n_342;
wire n_9369;
wire n_21179;
wire n_8305;
wire n_16557;
wire n_14458;
wire n_2072;
wire n_2738;
wire n_10730;
wire n_13095;
wire n_14856;
wire n_19607;
wire n_7779;
wire n_2968;
wire n_7316;
wire n_13612;
wire n_6098;
wire n_7019;
wire n_5062;
wire n_10202;
wire n_11398;
wire n_20085;
wire n_4469;
wire n_190;
wire n_7452;
wire n_8939;
wire n_16656;
wire n_3349;
wire n_12269;
wire n_7195;
wire n_6701;
wire n_7478;
wire n_20282;
wire n_16822;
wire n_19038;
wire n_2062;
wire n_12019;
wire n_14263;
wire n_14824;
wire n_2100;
wire n_3310;
wire n_18827;
wire n_748;
wire n_1058;
wire n_15995;
wire n_8440;
wire n_332;
wire n_1053;
wire n_21130;
wire n_10367;
wire n_4504;
wire n_9570;
wire n_15040;
wire n_15981;
wire n_20922;
wire n_1385;
wire n_793;
wire n_4408;
wire n_17166;
wire n_1819;
wire n_476;
wire n_2987;
wire n_16314;
wire n_11099;
wire n_4567;
wire n_4164;
wire n_4234;
wire n_11859;
wire n_18906;
wire n_5348;
wire n_7873;
wire n_16154;
wire n_2606;
wire n_18815;
wire n_3187;
wire n_20395;
wire n_8729;
wire n_16141;
wire n_19577;
wire n_6550;
wire n_17852;
wire n_19916;
wire n_5031;
wire n_17744;
wire n_3392;
wire n_4444;
wire n_5709;
wire n_10803;
wire n_16179;
wire n_3331;
wire n_2911;
wire n_10187;
wire n_2154;
wire n_14698;
wire n_18135;
wire n_5860;
wire n_6926;
wire n_9607;
wire n_4302;
wire n_21304;
wire n_8228;
wire n_10586;
wire n_6956;
wire n_10040;
wire n_21116;
wire n_5381;
wire n_3257;
wire n_2293;
wire n_11911;
wire n_17603;
wire n_9262;
wire n_2028;
wire n_15649;
wire n_558;
wire n_8387;
wire n_21377;
wire n_1412;
wire n_12782;
wire n_3981;
wire n_9761;
wire n_17612;
wire n_20718;
wire n_11039;
wire n_10164;
wire n_10269;
wire n_12567;
wire n_14228;
wire n_15264;
wire n_20581;
wire n_3224;
wire n_6342;
wire n_14854;
wire n_19375;
wire n_7308;
wire n_15828;
wire n_17822;
wire n_434;
wire n_18477;
wire n_21320;
wire n_21573;
wire n_12153;
wire n_935;
wire n_11730;
wire n_18194;
wire n_817;
wire n_1175;
wire n_10918;
wire n_18078;
wire n_20415;
wire n_13629;
wire n_14671;
wire n_17525;
wire n_14265;
wire n_13351;
wire n_17450;
wire n_8843;
wire n_11942;
wire n_4028;
wire n_19542;
wire n_13083;
wire n_3819;
wire n_7974;
wire n_16814;
wire n_18850;
wire n_17867;
wire n_431;
wire n_6503;
wire n_5888;
wire n_17319;
wire n_11835;
wire n_10598;
wire n_16031;
wire n_14797;
wire n_16555;
wire n_4731;
wire n_11444;
wire n_5592;
wire n_12430;
wire n_21459;
wire n_4618;
wire n_17406;
wire n_13971;
wire n_15798;
wire n_4099;
wire n_3484;
wire n_21156;
wire n_9646;
wire n_5303;
wire n_21725;
wire n_11205;
wire n_17489;
wire n_14093;
wire n_14150;
wire n_10436;
wire n_4603;
wire n_21681;
wire n_19676;
wire n_11048;
wire n_18781;
wire n_19529;
wire n_13172;
wire n_2607;
wire n_16766;
wire n_19556;
wire n_20481;
wire n_16935;
wire n_3317;
wire n_11782;
wire n_20100;
wire n_10538;
wire n_2582;
wire n_12258;
wire n_4283;
wire n_4681;
wire n_16500;
wire n_15743;
wire n_9918;
wire n_4638;
wire n_8159;
wire n_3455;
wire n_11397;
wire n_20955;
wire n_5346;
wire n_5517;
wire n_7797;
wire n_8216;
wire n_4707;
wire n_14979;
wire n_13887;
wire n_16238;
wire n_17323;
wire n_10924;
wire n_20912;
wire n_12871;
wire n_2342;
wire n_10942;
wire n_12295;
wire n_14171;
wire n_9956;
wire n_15134;
wire n_18864;
wire n_4848;
wire n_9715;
wire n_15679;
wire n_18618;
wire n_14141;
wire n_19037;
wire n_10292;
wire n_12077;
wire n_12166;
wire n_17962;
wire n_5624;
wire n_394;
wire n_21404;
wire n_11945;
wire n_12216;
wire n_2869;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_18459;
wire n_19947;
wire n_19920;
wire n_9931;
wire n_12098;
wire n_13749;
wire n_15064;
wire n_12102;
wire n_13009;
wire n_18284;
wire n_14325;
wire n_16682;
wire n_13535;
wire n_10624;
wire n_16254;
wire n_6568;
wire n_2857;
wire n_8295;
wire n_13668;
wire n_15124;
wire n_14836;
wire n_19865;
wire n_14292;
wire n_8995;
wire n_8146;
wire n_14583;
wire n_1596;
wire n_8082;
wire n_13046;
wire n_978;
wire n_20643;
wire n_19327;
wire n_7183;
wire n_1474;
wire n_16693;
wire n_19158;
wire n_15617;
wire n_6411;
wire n_2093;
wire n_9195;
wire n_12768;
wire n_10701;
wire n_14233;
wire n_15848;
wire n_15253;
wire n_4632;
wire n_20559;
wire n_16607;
wire n_14505;
wire n_12483;
wire n_21880;
wire n_16019;
wire n_14121;
wire n_4949;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_17011;
wire n_12682;
wire n_7223;
wire n_1758;
wire n_7890;
wire n_21882;
wire n_6179;
wire n_9281;
wire n_9475;
wire n_16850;
wire n_8865;
wire n_13056;
wire n_17575;
wire n_12313;
wire n_7165;
wire n_8110;
wire n_17290;
wire n_6223;
wire n_8475;
wire n_6435;
wire n_9143;
wire n_168;
wire n_974;
wire n_727;
wire n_957;
wire n_15785;
wire n_21389;
wire n_7795;
wire n_7404;
wire n_11147;
wire n_11700;
wire n_3597;
wire n_9087;
wire n_8119;
wire n_15227;
wire n_10135;
wire n_7885;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_11833;
wire n_19603;
wire n_5014;
wire n_1127;
wire n_9186;
wire n_15266;
wire n_1785;
wire n_2829;
wire n_6846;
wire n_9243;
wire n_14346;
wire n_3200;
wire n_14902;
wire n_11057;
wire n_6041;
wire n_7822;
wire n_12186;
wire n_2604;
wire n_17931;
wire n_4257;
wire n_3213;
wire n_20035;
wire n_15357;
wire n_13598;
wire n_17054;
wire n_11783;
wire n_21509;
wire n_16451;
wire n_11026;
wire n_14990;
wire n_14806;
wire n_2106;
wire n_17091;
wire n_12939;
wire n_4665;
wire n_1823;
wire n_20192;
wire n_14708;
wire n_7696;
wire n_17630;
wire n_11232;
wire n_5670;
wire n_9171;
wire n_1875;
wire n_18244;
wire n_1324;
wire n_19668;
wire n_17381;
wire n_21647;
wire n_19184;
wire n_860;
wire n_3229;
wire n_4463;
wire n_16863;
wire n_1805;
wire n_7958;
wire n_17770;
wire n_16368;
wire n_948;
wire n_5751;
wire n_4670;
wire n_15013;
wire n_4084;
wire n_4703;
wire n_15014;
wire n_18544;
wire n_8667;
wire n_3499;
wire n_16323;
wire n_19843;
wire n_15710;
wire n_16286;
wire n_14001;
wire n_6824;
wire n_11767;
wire n_8717;
wire n_1552;
wire n_6189;
wire n_3618;
wire n_20580;
wire n_2593;
wire n_19817;
wire n_16483;
wire n_19473;
wire n_6993;
wire n_20587;
wire n_6037;
wire n_3642;
wire n_3808;
wire n_8892;
wire n_359;
wire n_19838;
wire n_14550;
wire n_9067;
wire n_12712;
wire n_815;
wire n_16374;
wire n_14604;
wire n_20837;
wire n_9074;
wire n_20764;
wire n_1381;
wire n_6418;
wire n_6564;
wire n_2301;
wire n_21128;
wire n_3583;
wire n_18941;
wire n_15150;
wire n_3560;
wire n_4714;
wire n_8197;
wire n_13733;
wire n_10052;
wire n_18455;
wire n_12309;
wire n_18371;
wire n_21574;
wire n_17403;
wire n_9843;
wire n_19010;
wire n_3020;
wire n_17568;
wire n_16913;
wire n_5441;
wire n_6517;
wire n_2910;
wire n_11579;
wire n_7350;
wire n_20863;
wire n_1467;
wire n_10369;
wire n_20551;
wire n_2163;
wire n_16366;
wire n_5885;
wire n_2254;
wire n_925;
wire n_2647;
wire n_13003;
wire n_8452;
wire n_4443;
wire n_4507;
wire n_2624;
wire n_10671;
wire n_8140;
wire n_13213;
wire n_8981;
wire n_16803;
wire n_3569;
wire n_968;
wire n_19172;
wire n_4348;
wire n_619;
wire n_12611;
wire n_19305;
wire n_13767;
wire n_3494;
wire n_20806;
wire n_20915;
wire n_12322;
wire n_12303;
wire n_12507;
wire n_21796;
wire n_17801;
wire n_21746;
wire n_7844;
wire n_3771;
wire n_683;
wire n_3110;
wire n_11882;
wire n_13802;
wire n_1057;
wire n_16754;
wire n_9665;
wire n_802;
wire n_11146;
wire n_5609;
wire n_19785;
wire n_5416;
wire n_4026;
wire n_19138;
wire n_4512;
wire n_1305;
wire n_13443;
wire n_7471;
wire n_18068;
wire n_21516;
wire n_6745;
wire n_19406;
wire n_16659;
wire n_4521;
wire n_8481;
wire n_19151;
wire n_4488;
wire n_15867;
wire n_2783;
wire n_19713;
wire n_3750;
wire n_19903;
wire n_15491;
wire n_18594;
wire n_18913;
wire n_4588;
wire n_14146;
wire n_15870;
wire n_18677;
wire n_3299;
wire n_12121;
wire n_7594;
wire n_7766;
wire n_7340;
wire n_10837;
wire n_20834;
wire n_972;
wire n_8205;
wire n_12116;
wire n_8651;
wire n_14260;
wire n_1200;
wire n_13621;
wire n_14999;
wire n_3568;
wire n_9255;
wire n_15873;
wire n_10039;
wire n_8828;
wire n_17080;
wire n_17995;
wire n_7603;
wire n_6138;
wire n_16825;
wire n_9034;
wire n_20168;
wire n_1329;
wire n_15611;
wire n_9601;
wire n_13173;
wire n_5692;
wire n_7494;
wire n_19022;
wire n_10887;
wire n_13253;
wire n_9967;
wire n_18855;
wire n_21131;
wire n_16621;
wire n_10735;
wire n_8739;
wire n_8133;
wire n_8919;
wire n_17697;
wire n_2429;
wire n_17624;
wire n_883;
wire n_15478;
wire n_17154;
wire n_7396;
wire n_9912;
wire n_16649;
wire n_16292;
wire n_7116;
wire n_12779;
wire n_4352;
wire n_4441;
wire n_918;
wire n_8318;
wire n_16170;
wire n_8542;
wire n_17007;
wire n_11059;
wire n_2364;
wire n_13514;
wire n_18487;
wire n_15502;
wire n_19573;
wire n_17553;
wire n_21918;
wire n_15095;
wire n_10411;
wire n_11643;
wire n_13199;
wire n_2393;
wire n_18333;
wire n_15068;
wire n_6300;
wire n_9609;
wire n_10172;
wire n_19004;
wire n_16642;
wire n_7815;
wire n_13407;
wire n_9046;
wire n_17534;
wire n_192;
wire n_15554;
wire n_5032;
wire n_1549;
wire n_6537;
wire n_655;
wire n_21279;
wire n_21713;
wire n_9864;
wire n_13521;
wire n_3240;
wire n_18101;
wire n_12485;
wire n_12408;
wire n_9300;
wire n_15749;
wire n_387;
wire n_17153;
wire n_12238;
wire n_16271;
wire n_16373;
wire n_398;
wire n_5112;
wire n_5386;
wire n_18380;
wire n_6783;
wire n_9353;
wire n_7465;
wire n_13720;
wire n_2295;
wire n_3931;
wire n_8293;
wire n_5017;
wire n_10754;
wire n_4710;
wire n_13565;
wire n_17542;
wire n_13685;
wire n_13129;
wire n_21111;
wire n_20960;
wire n_6459;
wire n_19276;
wire n_16569;
wire n_2800;
wire n_16257;
wire n_5644;
wire n_3409;
wire n_8078;
wire n_10413;
wire n_12587;
wire n_4867;
wire n_17861;
wire n_15222;
wire n_19281;
wire n_21793;
wire n_21218;
wire n_17847;
wire n_15890;
wire n_6977;
wire n_7984;
wire n_14426;
wire n_4411;
wire n_11821;
wire n_8361;
wire n_6313;
wire n_16378;
wire n_16337;
wire n_15757;
wire n_149;
wire n_4777;
wire n_2653;
wire n_836;
wire n_20076;
wire n_17629;
wire n_6555;
wire n_16745;
wire n_14329;
wire n_13653;
wire n_7516;
wire n_15552;
wire n_13640;
wire n_5864;
wire n_6536;
wire n_3459;
wire n_3155;
wire n_8301;
wire n_19262;
wire n_1392;
wire n_3911;
wire n_19983;
wire n_6294;
wire n_18466;
wire n_7427;
wire n_21702;
wire n_13962;
wire n_17486;
wire n_12162;
wire n_20529;
wire n_4885;
wire n_7838;
wire n_7786;
wire n_21192;
wire n_9580;
wire n_5804;
wire n_18483;
wire n_12236;
wire n_6376;
wire n_3565;
wire n_7926;
wire n_2575;
wire n_7411;
wire n_12632;
wire n_17779;
wire n_5040;
wire n_6730;
wire n_10487;
wire n_13479;
wire n_15453;
wire n_6996;
wire n_9817;
wire n_15389;
wire n_1345;
wire n_1899;
wire n_8753;
wire n_7731;
wire n_11290;
wire n_15739;
wire n_2067;
wire n_8044;
wire n_15937;
wire n_14137;
wire n_2877;
wire n_7709;
wire n_9689;
wire n_3035;
wire n_21183;
wire n_19666;
wire n_21101;
wire n_19236;
wire n_6710;
wire n_7162;
wire n_18230;
wire n_1657;
wire n_19194;
wire n_768;
wire n_1475;
wire n_16096;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_9886;
wire n_1491;
wire n_20047;
wire n_12837;
wire n_18286;
wire n_17193;
wire n_735;
wire n_2501;
wire n_19874;
wire n_10264;
wire n_6426;
wire n_6634;
wire n_6836;
wire n_15735;
wire n_18379;
wire n_19470;
wire n_5197;
wire n_15792;
wire n_1979;
wire n_9297;
wire n_13460;
wire n_8788;
wire n_7111;
wire n_7549;
wire n_16978;
wire n_2484;
wire n_20288;
wire n_20648;
wire n_3731;
wire n_15849;
wire n_20841;
wire n_17928;
wire n_5994;
wire n_435;
wire n_766;
wire n_20707;
wire n_541;
wire n_15791;
wire n_15696;
wire n_13088;
wire n_8061;
wire n_6833;
wire n_21386;
wire n_687;
wire n_20263;
wire n_2489;
wire n_20556;
wire n_11103;
wire n_7481;
wire n_17177;
wire n_10341;
wire n_20106;
wire n_12230;
wire n_14511;
wire n_14176;
wire n_12995;
wire n_21944;
wire n_3561;
wire n_10498;
wire n_21373;
wire n_1011;
wire n_10508;
wire n_9662;
wire n_3536;
wire n_16610;
wire n_12406;
wire n_6821;
wire n_15740;
wire n_18419;
wire n_8545;
wire n_12725;
wire n_5788;
wire n_13404;
wire n_20026;
wire n_16534;
wire n_2103;
wire n_10865;
wire n_16984;
wire n_12185;
wire n_18399;
wire n_850;
wire n_8683;
wire n_17983;
wire n_15293;
wire n_10081;
wire n_2372;
wire n_7016;
wire n_6347;
wire n_19286;
wire n_15756;
wire n_15676;
wire n_9448;
wire n_17919;
wire n_353;
wire n_9799;
wire n_9313;
wire n_493;
wire n_2433;
wire n_7955;
wire n_19461;
wire n_7072;
wire n_5582;
wire n_7374;
wire n_20789;
wire n_12114;
wire n_13171;
wire n_11967;
wire n_9438;
wire n_7201;
wire n_2316;
wire n_1898;
wire n_12571;
wire n_10036;
wire n_20289;
wire n_15559;
wire n_10853;
wire n_12508;
wire n_12582;
wire n_12052;
wire n_2687;
wire n_1120;
wire n_4220;
wire n_1944;
wire n_5630;
wire n_1497;
wire n_3151;
wire n_20647;
wire n_4066;
wire n_11803;
wire n_16690;
wire n_11067;
wire n_12610;
wire n_5264;
wire n_1981;
wire n_7540;
wire n_4858;
wire n_15829;
wire n_18640;
wire n_19675;
wire n_14392;
wire n_15373;
wire n_7005;
wire n_1518;
wire n_18720;
wire n_15216;
wire n_14115;
wire n_12592;
wire n_1889;
wire n_14282;
wire n_13938;
wire n_2966;
wire n_14615;
wire n_1569;
wire n_20692;
wire n_11413;
wire n_19466;
wire n_19167;
wire n_6205;
wire n_19285;
wire n_21451;
wire n_756;
wire n_4456;
wire n_7607;
wire n_15973;
wire n_9159;
wire n_399;
wire n_16309;
wire n_15317;
wire n_4346;
wire n_21575;
wire n_13290;
wire n_3170;
wire n_7830;
wire n_8302;
wire n_17892;
wire n_21452;
wire n_11682;
wire n_17986;
wire n_12801;
wire n_11091;
wire n_15325;
wire n_11929;
wire n_17863;
wire n_760;
wire n_17954;
wire n_6668;
wire n_220;
wire n_18905;
wire n_15952;
wire n_1945;
wire n_3018;
wire n_7053;
wire n_8724;
wire n_14702;
wire n_19479;
wire n_5831;
wire n_12552;
wire n_8070;
wire n_6835;
wire n_13039;
wire n_14305;
wire n_17492;
wire n_4764;
wire n_19096;
wire n_9509;
wire n_6258;
wire n_167;
wire n_16601;
wire n_12256;
wire n_10057;
wire n_377;
wire n_4581;
wire n_12184;
wire n_11093;
wire n_19908;
wire n_21583;
wire n_8411;
wire n_12657;
wire n_19161;
wire n_2488;
wire n_13957;
wire n_7211;
wire n_20596;
wire n_6531;
wire n_8689;
wire n_19279;
wire n_771;
wire n_4782;
wire n_17271;
wire n_1520;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_10141;
wire n_20176;
wire n_1411;
wire n_8549;
wire n_3054;
wire n_18622;
wire n_21263;
wire n_19694;
wire n_2703;
wire n_10929;
wire n_16785;
wire n_8658;
wire n_9959;
wire n_5428;
wire n_10261;
wire n_12285;
wire n_16180;
wire n_3391;
wire n_6102;
wire n_21442;
wire n_9818;
wire n_5678;
wire n_4056;
wire n_21030;
wire n_1246;
wire n_2956;
wire n_19202;
wire n_19123;
wire n_19815;
wire n_8676;
wire n_15413;
wire n_19030;
wire n_871;
wire n_13496;
wire n_7929;
wire n_10028;
wire n_8399;
wire n_18710;
wire n_15363;
wire n_11069;
wire n_19716;
wire n_5116;
wire n_3464;
wire n_19259;
wire n_17746;
wire n_13818;
wire n_9304;
wire n_10777;
wire n_6632;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_18335;
wire n_9830;
wire n_21718;
wire n_9913;
wire n_11728;
wire n_3076;
wire n_16563;
wire n_3535;
wire n_17008;
wire n_20469;
wire n_11796;
wire n_8754;
wire n_7898;
wire n_10715;
wire n_12136;
wire n_16770;
wire n_6359;
wire n_20441;
wire n_17963;
wire n_2146;
wire n_13154;
wire n_19116;
wire n_3935;
wire n_7377;
wire n_11228;
wire n_542;
wire n_5379;
wire n_16458;
wire n_3948;
wire n_12517;
wire n_16173;
wire n_20293;
wire n_16875;
wire n_20645;
wire n_6301;
wire n_3232;
wire n_1673;
wire n_14850;
wire n_11261;
wire n_17623;
wire n_3125;
wire n_11023;
wire n_11382;
wire n_20576;
wire n_14278;
wire n_20349;
wire n_8602;
wire n_7381;
wire n_7948;
wire n_20554;
wire n_16449;
wire n_3951;
wire n_19284;
wire n_11305;
wire n_12680;
wire n_19702;
wire n_17202;
wire n_15511;
wire n_7430;
wire n_9700;
wire n_18356;
wire n_8871;
wire n_480;
wire n_425;
wire n_9476;
wire n_20080;
wire n_695;
wire n_21635;
wire n_20754;
wire n_8824;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_18154;
wire n_16058;
wire n_20663;
wire n_21792;
wire n_15533;
wire n_21393;
wire n_14160;
wire n_15576;
wire n_20614;
wire n_12666;
wire n_9882;
wire n_12205;
wire n_13177;
wire n_6145;
wire n_3577;
wire n_21906;
wire n_10242;
wire n_20544;
wire n_14899;
wire n_17641;
wire n_14166;
wire n_21888;
wire n_4314;
wire n_1621;
wire n_17078;
wire n_7846;
wire n_6076;
wire n_4288;
wire n_3567;
wire n_16549;
wire n_10673;
wire n_19409;
wire n_19737;
wire n_12917;
wire n_1634;
wire n_5843;
wire n_3321;
wire n_666;
wire n_14356;
wire n_3152;
wire n_20610;
wire n_12950;
wire n_7489;
wire n_18016;
wire n_18005;
wire n_15197;
wire n_6335;
wire n_18806;
wire n_16516;
wire n_2247;
wire n_7451;
wire n_17856;
wire n_19758;
wire n_15780;
wire n_16677;
wire n_12962;
wire n_3778;
wire n_17317;
wire n_1729;
wire n_19882;
wire n_2739;
wire n_15706;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_19249;
wire n_9702;
wire n_3256;
wire n_2386;
wire n_15301;
wire n_17351;
wire n_4217;
wire n_8807;
wire n_14207;
wire n_1099;
wire n_9924;
wire n_16848;
wire n_8732;
wire n_15954;
wire n_1738;
wire n_3728;
wire n_17835;
wire n_3088;
wire n_10527;
wire n_6951;
wire n_3713;
wire n_17294;
wire n_12584;
wire n_5046;
wire n_9252;
wire n_3246;
wire n_819;
wire n_12999;
wire n_14084;
wire n_21159;
wire n_13120;
wire n_5088;
wire n_16596;
wire n_19608;
wire n_15123;
wire n_7986;
wire n_6950;
wire n_417;
wire n_20799;
wire n_933;
wire n_11705;
wire n_8203;
wire n_14587;
wire n_16988;
wire n_7663;
wire n_13125;
wire n_11521;
wire n_17780;
wire n_14513;
wire n_2024;
wire n_14910;
wire n_755;
wire n_14590;
wire n_12293;
wire n_530;
wire n_17178;
wire n_13069;
wire n_18698;
wire n_21773;
wire n_15094;
wire n_3832;
wire n_22003;
wire n_17157;
wire n_16258;
wire n_5824;
wire n_11533;
wire n_17258;
wire n_5538;
wire n_6658;
wire n_10863;
wire n_15344;
wire n_17539;
wire n_10077;
wire n_18637;
wire n_9144;
wire n_7767;
wire n_13352;
wire n_21347;
wire n_20900;
wire n_15035;
wire n_13953;
wire n_18696;
wire n_21227;
wire n_20947;
wire n_7672;
wire n_4525;
wire n_12118;
wire n_3782;
wire n_9850;
wire n_14940;
wire n_6864;
wire n_13453;
wire n_11549;
wire n_7158;
wire n_2888;
wire n_19599;
wire n_6494;
wire n_8323;
wire n_1236;
wire n_12353;
wire n_8296;
wire n_13846;
wire n_17615;
wire n_10417;
wire n_9430;
wire n_17413;
wire n_10310;
wire n_335;
wire n_7504;
wire n_10333;
wire n_3489;
wire n_21422;
wire n_343;
wire n_8448;
wire n_20910;
wire n_16715;
wire n_5129;
wire n_7375;
wire n_5500;
wire n_15215;
wire n_12006;
wire n_16196;
wire n_5219;
wire n_16664;
wire n_14935;
wire n_3049;
wire n_16315;
wire n_21692;
wire n_8557;
wire n_19562;
wire n_21403;
wire n_1097;
wire n_1036;
wire n_6863;
wire n_9541;
wire n_18985;
wire n_13477;
wire n_21628;
wire n_15469;
wire n_7876;
wire n_6050;
wire n_15329;
wire n_15309;
wire n_15709;
wire n_7960;
wire n_17837;
wire n_670;
wire n_18607;
wire n_19112;
wire n_9555;
wire n_10959;
wire n_19861;
wire n_2551;
wire n_9994;
wire n_17950;
wire n_8538;
wire n_7043;
wire n_12753;
wire n_16248;
wire n_16945;
wire n_10859;
wire n_18981;
wire n_7751;
wire n_19304;
wire n_15430;
wire n_9142;
wire n_2699;
wire n_888;
wire n_3542;
wire n_20463;
wire n_5491;
wire n_3940;
wire n_8300;
wire n_2985;
wire n_5636;
wire n_7719;
wire n_9202;
wire n_2753;
wire n_8451;
wire n_18352;
wire n_2842;
wire n_4523;
wire n_10941;
wire n_11448;
wire n_5084;
wire n_8435;
wire n_3570;
wire n_5260;
wire n_18655;
wire n_9788;
wire n_19771;
wire n_13722;
wire n_2712;
wire n_14060;
wire n_14936;
wire n_19087;
wire n_6354;
wire n_5918;
wire n_18808;
wire n_19456;
wire n_4464;
wire n_17180;
wire n_17644;
wire n_15473;
wire n_3096;
wire n_989;
wire n_2544;
wire n_18254;
wire n_892;
wire n_9392;
wire n_18659;
wire n_6667;
wire n_12491;
wire n_14498;
wire n_6156;
wire n_13966;
wire n_21982;
wire n_5913;
wire n_5621;
wire n_13437;
wire n_2919;
wire n_8213;
wire n_7973;
wire n_18676;
wire n_18304;
wire n_13423;
wire n_15914;
wire n_17139;
wire n_2241;
wire n_2757;
wire n_8532;
wire n_15199;
wire n_21318;
wire n_11172;
wire n_8043;
wire n_20755;
wire n_7969;
wire n_6248;
wire n_884;
wire n_18018;
wire n_19691;
wire n_2921;
wire n_2720;
wire n_6088;
wire n_6894;
wire n_21745;
wire n_1856;
wire n_7267;
wire n_4959;
wire n_14520;
wire n_9898;
wire n_237;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_17079;
wire n_21754;
wire n_14669;
wire n_4103;
wire n_6204;
wire n_21235;
wire n_13951;
wire n_15236;
wire n_17329;
wire n_16110;
wire n_10921;
wire n_794;
wire n_7387;
wire n_10551;
wire n_16783;
wire n_2837;
wire n_21997;
wire n_5257;
wire n_4765;
wire n_18934;
wire n_702;
wire n_12364;
wire n_21949;
wire n_2108;
wire n_14785;
wire n_13697;
wire n_20969;
wire n_19868;
wire n_1538;
wire n_1779;
wire n_20977;
wire n_8359;
wire n_16345;
wire n_1369;
wire n_19546;
wire n_21087;
wire n_8211;
wire n_17795;
wire n_13943;
wire n_14814;
wire n_10871;
wire n_3207;
wire n_15434;
wire n_21989;
wire n_8943;
wire n_809;
wire n_8441;
wire n_10747;
wire n_15322;
wire n_5012;
wire n_1293;
wire n_15558;
wire n_4620;
wire n_11387;
wire n_8198;
wire n_15596;
wire n_15945;
wire n_7188;
wire n_8526;
wire n_10705;
wire n_2813;
wire n_2009;
wire n_18185;
wire n_6147;
wire n_17969;
wire n_3218;
wire n_21015;
wire n_10334;
wire n_11358;
wire n_18180;
wire n_6011;
wire n_7722;
wire n_8592;
wire n_747;
wire n_16343;
wire n_4325;
wire n_10235;
wire n_13247;
wire n_10153;
wire n_7193;
wire n_17185;
wire n_11489;
wire n_6897;
wire n_20071;
wire n_12420;
wire n_18626;
wire n_9071;
wire n_2629;
wire n_12314;
wire n_4379;
wire n_7128;
wire n_11373;
wire n_5882;
wire n_9606;
wire n_7881;
wire n_14416;
wire n_18156;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_10998;
wire n_21993;
wire n_9492;
wire n_13271;
wire n_19712;
wire n_18195;
wire n_9031;
wire n_17904;
wire n_18127;
wire n_11434;
wire n_11645;
wire n_4179;
wire n_18951;
wire n_9991;
wire n_18946;
wire n_11254;
wire n_13693;
wire n_14277;
wire n_368;
wire n_17798;
wire n_20218;
wire n_2539;
wire n_10253;
wire n_7248;
wire n_5339;
wire n_13376;
wire n_6099;
wire n_10946;
wire n_1617;
wire n_6904;
wire n_3760;
wire n_20334;
wire n_1760;
wire n_15480;
wire n_17497;
wire n_2856;
wire n_15651;
wire n_10473;
wire n_20605;
wire n_13104;
wire n_15339;
wire n_10893;
wire n_7533;
wire n_11548;
wire n_9777;
wire n_21240;
wire n_4787;
wire n_3667;
wire n_878;
wire n_16513;
wire n_18245;
wire n_10148;
wire n_9366;
wire n_11248;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_15669;
wire n_2787;
wire n_18234;
wire n_11901;
wire n_6116;
wire n_16081;
wire n_10337;
wire n_16912;
wire n_9869;
wire n_19182;
wire n_6819;
wire n_13929;
wire n_7936;
wire n_9741;
wire n_10956;
wire n_12131;
wire n_16834;
wire n_8391;
wire n_18518;
wire n_11381;
wire n_2982;
wire n_12453;
wire n_17887;
wire n_3545;
wire n_17305;
wire n_12557;
wire n_20639;
wire n_20634;
wire n_15295;
wire n_20223;
wire n_1614;
wire n_20539;
wire n_7148;
wire n_15582;
wire n_5782;
wire n_8340;
wire n_7250;
wire n_7828;
wire n_12020;
wire n_19336;
wire n_4935;
wire n_8691;
wire n_16044;
wire n_4785;
wire n_3820;
wire n_3454;
wire n_13502;
wire n_13468;
wire n_20825;
wire n_12920;
wire n_13403;
wire n_12785;
wire n_17654;
wire n_8704;
wire n_6355;
wire n_5596;
wire n_16787;
wire n_10078;
wire n_16162;
wire n_2346;
wire n_13201;
wire n_19576;
wire n_3990;
wire n_11106;
wire n_1215;
wire n_17967;
wire n_9289;
wire n_14687;
wire n_10827;
wire n_18685;
wire n_20442;
wire n_11218;
wire n_7356;
wire n_13291;
wire n_7294;
wire n_12629;
wire n_21750;
wire n_5290;
wire n_12972;
wire n_7018;
wire n_17515;
wire n_2721;
wire n_11167;
wire n_13440;
wire n_21722;
wire n_10452;
wire n_8707;
wire n_3002;
wire n_337;
wire n_19485;
wire n_5324;
wire n_18362;
wire n_7108;
wire n_21247;
wire n_9125;
wire n_8552;
wire n_7888;
wire n_17272;
wire n_14460;
wire n_13111;
wire n_11884;
wire n_12727;
wire n_1416;
wire n_1724;
wire n_18712;
wire n_3458;
wire n_21858;
wire n_6966;
wire n_9228;
wire n_14828;
wire n_15131;
wire n_21039;
wire n_12227;
wire n_1486;
wire n_12597;
wire n_7218;
wire n_3519;
wire n_7221;
wire n_10967;
wire n_8289;
wire n_14189;
wire n_16021;
wire n_3045;
wire n_15057;
wire n_22005;
wire n_13568;
wire n_13029;
wire n_19731;
wire n_2896;
wire n_13647;
wire n_19454;
wire n_17729;
wire n_4074;
wire n_15977;
wire n_12674;
wire n_5583;
wire n_11826;
wire n_1349;
wire n_4460;
wire n_11317;
wire n_19809;
wire n_3223;
wire n_21987;
wire n_10742;
wire n_14538;
wire n_19765;
wire n_12913;
wire n_2255;
wire n_1965;
wire n_9365;
wire n_1902;
wire n_14021;
wire n_20262;
wire n_3938;
wire n_11033;
wire n_18207;
wire n_19181;
wire n_6135;
wire n_14037;
wire n_11798;
wire n_3498;
wire n_2015;
wire n_19630;
wire n_17470;
wire n_21687;
wire n_993;
wire n_17461;
wire n_20072;
wire n_545;
wire n_21542;
wire n_450;
wire n_21810;
wire n_11079;
wire n_6141;
wire n_21229;
wire n_17589;
wire n_3965;
wire n_4349;
wire n_14931;
wire n_8493;
wire n_19100;
wire n_3788;
wire n_12400;
wire n_10244;
wire n_17989;
wire n_4313;
wire n_17902;
wire n_1935;
wire n_20171;
wire n_11469;
wire n_8958;
wire n_2696;
wire n_17149;
wire n_21134;
wire n_3242;
wire n_9624;
wire n_8161;
wire n_16403;
wire n_21581;
wire n_8734;
wire n_11341;
wire n_21651;
wire n_9901;
wire n_11619;
wire n_13378;
wire n_12756;
wire n_17926;
wire n_5100;
wire n_9189;
wire n_5849;
wire n_8495;
wire n_14255;
wire n_2578;
wire n_12218;
wire n_6635;
wire n_1821;
wire n_20162;
wire n_3894;
wire n_9472;
wire n_17757;
wire n_11553;
wire n_4015;
wire n_3890;
wire n_5367;
wire n_16802;
wire n_8994;
wire n_8901;
wire n_10725;
wire n_19856;
wire n_17800;
wire n_17788;
wire n_12387;
wire n_10627;
wire n_15846;
wire n_3524;
wire n_5034;
wire n_5988;
wire n_15194;
wire n_14651;
wire n_20136;
wire n_19157;
wire n_12798;
wire n_3549;
wire n_11032;
wire n_2092;
wire n_9434;
wire n_10604;
wire n_11110;
wire n_5959;
wire n_9052;
wire n_7645;
wire n_17020;
wire n_1776;
wire n_12780;
wire n_19063;
wire n_15314;
wire n_3026;
wire n_8157;
wire n_13651;
wire n_13830;
wire n_16307;
wire n_8309;
wire n_14998;
wire n_1047;
wire n_12589;
wire n_5754;
wire n_21986;
wire n_8096;
wire n_20571;
wire n_12043;
wire n_20165;
wire n_8222;
wire n_18795;
wire n_19978;
wire n_11971;
wire n_6726;
wire n_2266;
wire n_11320;
wire n_6554;
wire n_21096;
wire n_18007;
wire n_19258;
wire n_967;
wire n_14245;
wire n_12476;
wire n_8866;
wire n_19451;
wire n_5614;
wire n_21343;
wire n_19604;
wire n_17362;
wire n_3976;
wire n_1357;
wire n_7355;
wire n_8794;
wire n_14993;
wire n_17543;
wire n_16079;
wire n_14241;
wire n_21328;
wire n_4840;
wire n_17917;
wire n_15235;
wire n_19029;
wire n_983;
wire n_1826;
wire n_1283;
wire n_5696;
wire n_12549;
wire n_19325;
wire n_6499;
wire n_6837;
wire n_13442;
wire n_15073;
wire n_13390;
wire n_7393;
wire n_9686;
wire n_3282;
wire n_13334;
wire n_821;
wire n_13408;
wire n_20708;
wire n_12018;
wire n_20050;
wire n_2475;
wire n_8333;
wire n_8055;
wire n_5064;
wire n_12060;
wire n_5753;
wire n_10628;
wire n_507;
wire n_19385;
wire n_21447;
wire n_17337;
wire n_5536;
wire n_1605;
wire n_14071;
wire n_5173;
wire n_19294;
wire n_6305;
wire n_1228;
wire n_3920;
wire n_10819;
wire n_12315;
wire n_5794;
wire n_13098;
wire n_5027;
wire n_14447;
wire n_12484;
wire n_3866;
wire n_779;
wire n_9964;
wire n_10356;
wire n_20888;
wire n_11711;
wire n_16604;
wire n_18395;
wire n_15107;
wire n_7014;
wire n_13424;
wire n_5635;
wire n_11350;
wire n_984;
wire n_9019;
wire n_11310;
wire n_15023;
wire n_5975;
wire n_20713;
wire n_21587;
wire n_8494;
wire n_7066;
wire n_20552;
wire n_12449;
wire n_9468;
wire n_11939;
wire n_21138;
wire n_16968;
wire n_18914;
wire n_3094;
wire n_17281;
wire n_15799;
wire n_2310;
wire n_18735;
wire n_20362;
wire n_6789;
wire n_17617;
wire n_12845;
wire n_18136;
wire n_2502;
wire n_4762;
wire n_21835;
wire n_2793;
wire n_7690;
wire n_15360;
wire n_15110;
wire n_9419;
wire n_2285;
wire n_18336;
wire n_12793;
wire n_3147;
wire n_21930;
wire n_14488;
wire n_12367;
wire n_1149;
wire n_19205;
wire n_7390;
wire n_17789;
wire n_18634;
wire n_10474;
wire n_13316;
wire n_1824;
wire n_9820;
wire n_12954;
wire n_178;
wire n_16716;
wire n_17452;
wire n_11839;
wire n_11815;
wire n_2588;
wire n_12773;
wire n_8153;
wire n_12556;
wire n_4668;
wire n_17439;
wire n_849;
wire n_12789;
wire n_584;
wire n_15201;
wire n_5284;
wire n_21396;
wire n_16807;
wire n_4997;
wire n_10573;
wire n_2627;
wire n_13101;
wire n_6768;
wire n_4759;
wire n_13893;
wire n_13494;
wire n_1413;
wire n_801;
wire n_4467;
wire n_7506;
wire n_2340;
wire n_14210;
wire n_16507;
wire n_14717;
wire n_18051;
wire n_17893;
wire n_18046;
wire n_4735;
wire n_15368;
wire n_10428;
wire n_15908;
wire n_19272;
wire n_16572;
wire n_10989;
wire n_11145;
wire n_15812;
wire n_11017;
wire n_19075;
wire n_18597;
wire n_15623;
wire n_21195;
wire n_1019;
wire n_8906;
wire n_304;
wire n_7416;
wire n_12404;
wire n_21420;
wire n_7330;
wire n_15950;
wire n_8477;
wire n_16704;
wire n_10433;
wire n_778;
wire n_4068;
wire n_6000;
wire n_3192;
wire n_18590;
wire n_6655;
wire n_5792;
wire n_21186;
wire n_12002;
wire n_20719;
wire n_18133;
wire n_1929;
wire n_11543;
wire n_2807;
wire n_2313;
wire n_489;
wire n_8122;
wire n_2558;
wire n_10796;
wire n_8536;
wire n_7474;
wire n_7612;
wire n_6113;
wire n_16155;
wire n_7789;
wire n_15826;
wire n_917;
wire n_18074;
wire n_7902;
wire n_20979;
wire n_15027;
wire n_16369;
wire n_12598;
wire n_6842;
wire n_13575;
wire n_3390;
wire n_12033;
wire n_1573;
wire n_21217;
wire n_16738;
wire n_21006;
wire n_2745;
wire n_6801;
wire n_17719;
wire n_9996;
wire n_11348;
wire n_7680;
wire n_18484;
wire n_19040;
wire n_7398;
wire n_1133;
wire n_4537;
wire n_16015;
wire n_21485;
wire n_9906;
wire n_18355;
wire n_21719;
wire n_6968;
wire n_9504;
wire n_16632;
wire n_6615;
wire n_16206;
wire n_12181;
wire n_15145;
wire n_5205;
wire n_16107;
wire n_9138;
wire n_9384;
wire n_2602;
wire n_19452;
wire n_14197;
wire n_8903;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_5998;
wire n_18288;
wire n_4105;
wire n_19774;
wire n_232;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_17387;
wire n_427;
wire n_11019;
wire n_20384;
wire n_8585;
wire n_21398;
wire n_8982;
wire n_6415;
wire n_21194;
wire n_6857;
wire n_10489;
wire n_2401;
wire n_15114;
wire n_5476;
wire n_7842;
wire n_5446;
wire n_20004;
wire n_18383;
wire n_3148;
wire n_16714;
wire n_5944;
wire n_7618;
wire n_2264;
wire n_16267;
wire n_20904;
wire n_16468;
wire n_6361;
wire n_11677;
wire n_9357;
wire n_4098;
wire n_15394;
wire n_16897;
wire n_5861;
wire n_5976;
wire n_11827;
wire n_16896;
wire n_1184;
wire n_20489;
wire n_16150;
wire n_3404;
wire n_19407;
wire n_4055;
wire n_2926;
wire n_626;
wire n_3540;
wire n_16905;
wire n_8692;
wire n_7167;
wire n_18650;
wire n_20468;
wire n_10380;
wire n_4442;
wire n_16829;
wire n_14809;
wire n_19376;
wire n_20376;
wire n_10530;
wire n_4779;
wire n_8062;
wire n_2286;
wire n_19111;
wire n_16826;
wire n_10203;
wire n_13860;
wire n_19538;
wire n_2065;
wire n_10061;
wire n_4017;
wire n_13359;
wire n_8233;
wire n_9747;
wire n_620;
wire n_6953;
wire n_1081;
wire n_2705;
wire n_9061;
wire n_9168;
wire n_11690;
wire n_2977;
wire n_18851;
wire n_11155;
wire n_5674;
wire n_21103;
wire n_245;
wire n_19051;
wire n_20676;
wire n_15060;
wire n_16795;
wire n_7993;
wire n_21593;
wire n_672;
wire n_20322;
wire n_16094;
wire n_18069;
wire n_19938;
wire n_16496;
wire n_9073;
wire n_3365;
wire n_3476;
wire n_11312;
wire n_21569;
wire n_265;
wire n_11988;
wire n_7963;
wire n_443;
wire n_6599;
wire n_14978;
wire n_12311;
wire n_12914;
wire n_1747;
wire n_9068;
wire n_10537;
wire n_12787;
wire n_19655;
wire n_19053;
wire n_4740;
wire n_17417;
wire n_9544;
wire n_14108;
wire n_7800;
wire n_14700;
wire n_17853;
wire n_15633;
wire n_12263;
wire n_21270;
wire n_12959;
wire n_1868;
wire n_1613;
wire n_7581;
wire n_10131;
wire n_4049;
wire n_941;
wire n_13057;
wire n_13990;
wire n_18450;
wire n_8789;
wire n_17358;
wire n_21832;
wire n_16325;
wire n_13876;
wire n_14438;
wire n_14382;
wire n_13128;
wire n_19967;
wire n_7678;
wire n_10082;
wire n_15299;
wire n_17197;
wire n_15390;
wire n_18813;
wire n_17683;
wire n_5526;
wire n_10152;
wire n_15063;
wire n_2818;
wire n_1100;
wire n_6195;
wire n_8927;
wire n_17238;
wire n_11055;
wire n_18256;
wire n_17649;
wire n_15824;
wire n_12090;
wire n_5021;
wire n_19906;
wire n_7829;
wire n_14131;
wire n_4382;
wire n_20257;
wire n_2138;
wire n_14457;
wire n_5230;
wire n_2260;
wire n_14398;
wire n_5389;
wire n_11597;
wire n_13716;
wire n_1172;
wire n_428;
wire n_12165;
wire n_1341;
wire n_15970;
wire n_21407;
wire n_17518;
wire n_3289;
wire n_18970;
wire n_8832;
wire n_15614;
wire n_20679;
wire n_9340;
wire n_18591;
wire n_8461;
wire n_15128;
wire n_10977;
wire n_6825;
wire n_20674;
wire n_21999;
wire n_1770;
wire n_19534;
wire n_4228;
wire n_11369;
wire n_17205;
wire n_20507;
wire n_6547;
wire n_19690;
wire n_14231;
wire n_16824;
wire n_1873;
wire n_20209;
wire n_221;
wire n_6275;
wire n_3472;
wire n_21009;
wire n_4877;
wire n_20450;
wire n_20891;
wire n_21594;
wire n_11376;
wire n_5030;
wire n_3949;
wire n_9823;
wire n_14304;
wire n_11812;
wire n_19212;
wire n_8455;
wire n_11838;
wire n_17057;
wire n_20995;
wire n_4834;
wire n_20923;
wire n_11333;
wire n_1364;
wire n_9595;
wire n_5272;
wire n_2183;
wire n_6826;
wire n_8372;
wire n_7551;
wire n_1367;
wire n_11188;
wire n_4562;
wire n_16540;
wire n_16456;
wire n_7750;
wire n_18226;
wire n_12525;
wire n_17400;
wire n_13093;
wire n_20369;
wire n_8616;
wire n_3115;
wire n_4390;
wire n_5302;
wire n_6752;
wire n_5545;
wire n_2209;
wire n_4270;
wire n_8135;
wire n_10295;
wire n_5152;
wire n_16508;
wire n_9258;
wire n_3680;
wire n_12693;
wire n_201;
wire n_20359;
wire n_12203;
wire n_20068;
wire n_6329;
wire n_2940;
wire n_8529;
wire n_9763;
wire n_1495;
wire n_5128;
wire n_18656;
wire n_9965;
wire n_3322;
wire n_21108;
wire n_846;
wire n_18949;
wire n_6905;
wire n_7425;
wire n_1914;
wire n_2335;
wire n_12933;
wire n_8967;
wire n_21498;
wire n_21458;
wire n_8719;
wire n_2349;
wire n_16098;
wire n_19642;
wire n_10678;
wire n_6215;
wire n_14645;
wire n_15901;
wire n_5770;
wire n_5892;
wire n_8762;
wire n_16477;
wire n_6899;
wire n_19132;
wire n_5802;
wire n_3522;
wire n_20012;
wire n_9803;
wire n_21597;
wire n_8977;
wire n_10978;
wire n_9755;
wire n_14997;
wire n_20131;
wire n_17306;
wire n_4563;
wire n_2210;
wire n_14361;
wire n_4169;
wire n_18973;
wire n_13447;
wire n_12410;
wire n_17846;
wire n_9917;
wire n_3066;
wire n_2426;
wire n_18936;
wire n_15315;
wire n_12182;
wire n_14096;
wire n_14943;
wire n_20445;
wire n_4881;
wire n_14007;
wire n_9522;
wire n_19539;
wire n_16134;
wire n_16580;
wire n_5271;
wire n_160;
wire n_10571;
wire n_13276;
wire n_13338;
wire n_12547;
wire n_20087;
wire n_5637;
wire n_12370;
wire n_4584;
wire n_8279;
wire n_14054;
wire n_18919;
wire n_3319;
wire n_5240;
wire n_5813;
wire n_13543;
wire n_5495;
wire n_9488;
wire n_7312;
wire n_19732;
wire n_7155;
wire n_9231;
wire n_6865;
wire n_3016;
wire n_16635;
wire n_1693;
wire n_16595;
wire n_5393;
wire n_904;
wire n_7213;
wire n_9047;
wire n_18831;
wire n_8270;
wire n_4209;
wire n_11072;
wire n_17996;
wire n_1542;
wire n_13781;
wire n_14223;
wire n_15871;
wire n_11605;
wire n_19892;
wire n_8054;
wire n_12419;
wire n_1751;
wire n_13760;
wire n_21629;
wire n_9979;
wire n_785;
wire n_9093;
wire n_11959;
wire n_15883;
wire n_6482;
wire n_13012;
wire n_15148;
wire n_12865;
wire n_7715;
wire n_11881;
wire n_15210;
wire n_3596;
wire n_7007;
wire n_3906;
wire n_10045;
wire n_14672;
wire n_18654;
wire n_155;
wire n_20120;
wire n_1370;
wire n_2388;
wire n_13102;
wire n_4292;
wire n_20197;
wire n_21067;
wire n_8281;
wire n_4202;
wire n_18587;
wire n_9976;
wire n_2853;
wire n_5939;
wire n_16429;
wire n_11258;
wire n_800;
wire n_9568;
wire n_15956;
wire n_20600;
wire n_8459;
wire n_20283;
wire n_17634;
wire n_12580;
wire n_4412;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_7122;
wire n_7567;
wire n_21873;
wire n_21307;
wire n_3815;
wire n_13607;
wire n_21599;
wire n_11563;
wire n_15089;
wire n_13292;
wire n_5259;
wire n_1118;
wire n_20426;
wire n_17448;
wire n_19931;
wire n_9079;
wire n_11846;
wire n_1359;
wire n_10383;
wire n_13377;
wire n_10064;
wire n_15637;
wire n_375;
wire n_2165;
wire n_16790;
wire n_8975;
wire n_20344;
wire n_3532;
wire n_9170;
wire n_1818;
wire n_1257;
wire n_18252;
wire n_3531;
wire n_12960;
wire n_17122;
wire n_13519;
wire n_18040;
wire n_13984;
wire n_10238;
wire n_8759;
wire n_4548;
wire n_5923;
wire n_5790;
wire n_21964;
wire n_21655;
wire n_21637;
wire n_14924;
wire n_2959;
wire n_9670;
wire n_12711;
wire n_6552;
wire n_1845;
wire n_20412;
wire n_8325;
wire n_6328;
wire n_4816;
wire n_231;
wire n_19013;
wire n_19174;
wire n_15815;
wire n_16281;
wire n_14049;
wire n_7159;
wire n_1289;
wire n_8889;
wire n_13643;
wire n_6978;
wire n_12104;
wire n_18616;
wire n_19430;
wire n_16611;
wire n_12467;
wire n_4483;
wire n_21303;
wire n_19143;
wire n_19693;
wire n_19555;
wire n_7477;
wire n_2643;
wire n_12386;
wire n_10213;
wire n_18089;
wire n_21734;
wire n_10872;
wire n_5997;
wire n_955;
wire n_3028;
wire n_4350;
wire n_7295;
wire n_21556;
wire n_15900;
wire n_19247;
wire n_6058;
wire n_550;
wire n_8956;
wire n_20733;
wire n_1428;
wire n_7831;
wire n_19214;
wire n_1216;
wire n_5235;
wire n_15234;
wire n_17620;
wire n_3963;
wire n_14564;
wire n_21463;
wire n_12339;
wire n_6170;
wire n_20604;
wire n_10669;
wire n_10895;
wire n_8641;
wire n_15903;
wire n_11610;
wire n_11187;
wire n_7466;
wire n_16246;
wire n_15255;
wire n_11280;
wire n_10757;
wire n_7651;
wire n_5103;
wire n_680;
wire n_20140;
wire n_8973;
wire n_6935;
wire n_21349;
wire n_11426;
wire n_18178;
wire n_9038;
wire n_17394;
wire n_1556;
wire n_14337;
wire n_2118;
wire n_5985;
wire n_2944;
wire n_14439;
wire n_468;
wire n_6907;
wire n_11706;
wire n_13284;
wire n_7661;
wire n_10782;
wire n_6541;
wire n_19912;
wire n_5896;
wire n_13303;
wire n_17490;
wire n_3690;
wire n_13813;
wire n_3716;
wire n_5133;
wire n_8412;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_6226;
wire n_21526;
wire n_20245;
wire n_11211;
wire n_9668;
wire n_2275;
wire n_3273;
wire n_17613;
wire n_9877;
wire n_4310;
wire n_1950;
wire n_2370;
wire n_9395;
wire n_17163;
wire n_20937;
wire n_18096;
wire n_14734;
wire n_9209;
wire n_5097;
wire n_19595;
wire n_15010;
wire n_21929;
wire n_15308;
wire n_18615;
wire n_3071;
wire n_3739;
wire n_593;
wire n_5816;
wire n_17391;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_7241;
wire n_18116;
wire n_11011;
wire n_10009;
wire n_11776;
wire n_4850;
wire n_17741;
wire n_11165;
wire n_4813;
wire n_17508;
wire n_21548;
wire n_8274;
wire n_16699;
wire n_18417;
wire n_8550;
wire n_8264;
wire n_12817;
wire n_18907;
wire n_9009;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_10044;
wire n_13207;
wire n_16219;
wire n_1825;
wire n_12586;
wire n_21353;
wire n_5400;
wire n_8266;
wire n_10169;
wire n_4252;
wire n_15707;
wire n_6063;
wire n_10329;
wire n_20337;
wire n_21148;
wire n_19293;
wire n_10891;
wire n_15099;
wire n_8946;
wire n_9716;
wire n_14543;
wire n_18532;
wire n_3481;
wire n_6890;
wire n_9116;
wire n_21644;
wire n_13308;
wire n_9006;
wire n_13381;
wire n_17112;
wire n_10029;
wire n_3514;
wire n_4132;
wire n_13483;
wire n_9852;
wire n_7543;
wire n_2611;
wire n_9914;
wire n_6184;
wire n_16157;
wire n_20269;
wire n_21354;
wire n_2529;
wire n_15466;
wire n_21950;
wire n_15874;
wire n_17945;
wire n_4001;
wire n_3047;
wire n_14873;
wire n_6716;
wire n_16043;
wire n_12776;
wire n_17484;
wire n_21259;
wire n_7475;
wire n_759;
wire n_12578;
wire n_4824;
wire n_4120;
wire n_11864;
wire n_3745;
wire n_14232;
wire n_21288;
wire n_2990;
wire n_18756;
wire n_21807;
wire n_20650;
wire n_9669;
wire n_9958;
wire n_4082;
wire n_4085;
wire n_4073;
wire n_16457;
wire n_1649;
wire n_4163;
wire n_17981;
wire n_13345;
wire n_3500;
wire n_9588;
wire n_21481;
wire n_2621;
wire n_13756;
wire n_19800;
wire n_19923;
wire n_17137;
wire n_2671;
wire n_6646;
wire n_8936;
wire n_8414;
wire n_15529;
wire n_10137;
wire n_17141;
wire n_11861;
wire n_17388;
wire n_6903;
wire n_9050;
wire n_11724;
wire n_14775;
wire n_13970;
wire n_18846;
wire n_10196;
wire n_4334;
wire n_1674;
wire n_18887;
wire n_20189;
wire n_19469;
wire n_8831;
wire n_18184;
wire n_18086;
wire n_14100;
wire n_15704;
wire n_139;
wire n_11459;
wire n_11355;
wire n_6604;
wire n_4014;
wire n_12267;
wire n_12569;
wire n_16903;
wire n_17111;
wire n_9640;
wire n_8348;
wire n_5607;
wire n_21741;
wire n_20419;
wire n_20981;
wire n_14452;
wire n_16046;
wire n_10840;
wire n_10335;
wire n_19316;
wire n_6566;
wire n_18103;
wire n_13152;
wire n_1443;
wire n_18897;
wire n_946;
wire n_19549;
wire n_4892;
wire n_16071;
wire n_3816;
wire n_12513;
wire n_12091;
wire n_6047;
wire n_14788;
wire n_12307;
wire n_18017;
wire n_11890;
wire n_8913;
wire n_18061;
wire n_15550;
wire n_8800;
wire n_6861;
wire n_13702;
wire n_2045;
wire n_2040;
wire n_10919;
wire n_3199;
wire n_17456;
wire n_3843;
wire n_12288;
wire n_18856;
wire n_12415;
wire n_13037;
wire n_9432;
wire n_16849;
wire n_20765;
wire n_3685;
wire n_4249;
wire n_7748;
wire n_20211;
wire n_12949;
wire n_7556;
wire n_8881;
wire n_9704;
wire n_4718;
wire n_3555;
wire n_3236;
wire n_20538;
wire n_12859;
wire n_3396;
wire n_11282;
wire n_1445;
wire n_21113;
wire n_7050;
wire n_4023;
wire n_9915;
wire n_14156;
wire n_4420;
wire n_14772;
wire n_5773;
wire n_12188;
wire n_12943;
wire n_16297;
wire n_7318;
wire n_15136;
wire n_10373;
wire n_6108;
wire n_16353;
wire n_14387;
wire n_16694;
wire n_13148;
wire n_15645;
wire n_484;
wire n_12588;
wire n_12652;
wire n_8523;
wire n_20523;
wire n_11458;
wire n_4396;
wire n_16855;
wire n_16214;
wire n_18057;
wire n_6480;
wire n_13531;
wire n_20275;
wire n_2087;
wire n_7733;
wire n_11255;
wire n_6597;
wire n_10561;
wire n_15282;
wire n_18097;
wire n_12523;
wire n_7817;
wire n_21334;
wire n_14312;
wire n_6933;
wire n_16411;
wire n_8338;
wire n_4951;
wire n_12579;
wire n_17952;
wire n_11442;
wire n_19031;
wire n_13052;
wire n_7289;
wire n_17002;
wire n_5805;
wire n_9552;
wire n_11008;
wire n_11243;
wire n_2399;
wire n_14659;
wire n_473;
wire n_17650;
wire n_18511;
wire n_16960;
wire n_2133;
wire n_8027;
wire n_10096;
wire n_3830;
wire n_11425;
wire n_6817;
wire n_11992;
wire n_614;
wire n_18803;
wire n_5175;
wire n_3883;
wire n_4152;
wire n_17000;
wire n_21268;
wire n_19019;
wire n_11536;
wire n_773;
wire n_17584;
wire n_9069;
wire n_8966;
wire n_142;
wire n_8487;
wire n_14995;
wire n_16570;
wire n_15817;
wire n_13471;
wire n_296;
wire n_11327;
wire n_8533;
wire n_4281;
wire n_21003;
wire n_19441;
wire n_4962;
wire n_14956;
wire n_15684;
wire n_20092;
wire n_1237;
wire n_6327;
wire n_11140;
wire n_761;
wire n_6607;
wire n_9188;
wire n_18334;
wire n_11078;
wire n_4958;
wire n_9743;
wire n_16422;
wire n_10749;
wire n_4921;
wire n_1980;
wire n_8911;
wire n_11352;
wire n_20125;
wire n_18932;
wire n_7725;
wire n_3065;
wire n_1093;
wire n_15039;
wire n_1265;
wire n_19695;
wire n_9113;
wire n_4945;
wire n_4732;
wire n_19671;
wire n_11986;
wire n_18064;
wire n_16959;
wire n_17848;
wire n_11734;
wire n_18272;
wire n_14222;
wire n_15054;
wire n_511;
wire n_358;
wire n_16352;
wire n_8354;
wire n_4326;
wire n_6695;
wire n_18402;
wire n_5383;
wire n_14598;
wire n_14446;
wire n_4305;
wire n_14747;
wire n_14909;
wire n_5781;
wire n_19110;
wire n_1407;
wire n_12010;
wire n_19781;
wire n_21359;
wire n_21244;
wire n_19531;
wire n_19121;
wire n_11427;
wire n_16365;
wire n_21820;
wire n_911;
wire n_9746;
wire n_9680;
wire n_1430;
wire n_4802;
wire n_9633;
wire n_513;
wire n_16499;
wire n_10884;
wire n_18718;
wire n_3029;
wire n_19297;
wire n_7586;
wire n_6719;
wire n_17333;
wire n_11475;
wire n_18820;
wire n_14191;
wire n_490;
wire n_18398;
wire n_21546;
wire n_2243;
wire n_13092;
wire n_13888;
wire n_8974;
wire n_16464;
wire n_14561;
wire n_2929;
wire n_3751;
wire n_10821;
wire n_1611;
wire n_8983;
wire n_19708;
wire n_9338;
wire n_19267;
wire n_6884;
wire n_2554;
wire n_8013;
wire n_19810;
wire n_3927;
wire n_1630;
wire n_6513;
wire n_12524;
wire n_21781;
wire n_7841;
wire n_391;
wire n_17072;
wire n_701;
wire n_20193;
wire n_1092;
wire n_16980;
wire n_12173;
wire n_6516;
wire n_10358;
wire n_7792;
wire n_6924;
wire n_21286;
wire n_12168;
wire n_12349;
wire n_19107;
wire n_5606;
wire n_4830;
wire n_20792;
wire n_11736;
wire n_5237;
wire n_20918;
wire n_21641;
wire n_1206;
wire n_17092;
wire n_7073;
wire n_21497;
wire n_11393;
wire n_5093;
wire n_4946;
wire n_21232;
wire n_20567;
wire n_21016;
wire n_14718;
wire n_9098;
wire n_4663;
wire n_1060;
wire n_5347;
wire n_9861;
wire n_3298;
wire n_3033;
wire n_6788;
wire n_13638;
wire n_14869;
wire n_19367;
wire n_18435;
wire n_1386;
wire n_19647;
wire n_17878;
wire n_12282;
wire n_19192;
wire n_20497;
wire n_2916;
wire n_6249;
wire n_483;
wire n_6849;
wire n_13268;
wire n_12431;
wire n_1066;
wire n_18219;
wire n_14595;
wire n_11281;
wire n_15218;
wire n_18065;
wire n_20491;
wire n_14215;
wire n_15437;
wire n_2870;
wire n_12830;
wire n_15991;
wire n_378;
wire n_6572;
wire n_4791;
wire n_11372;
wire n_14781;
wire n_5151;
wire n_7003;
wire n_18727;
wire n_21645;
wire n_7897;
wire n_4773;
wire n_17160;
wire n_14954;
wire n_21555;
wire n_7962;
wire n_4497;
wire n_8113;
wire n_5982;
wire n_1768;
wire n_21721;
wire n_10308;
wire n_17640;
wire n_1719;
wire n_4658;
wire n_15711;
wire n_19591;
wire n_5827;
wire n_15298;
wire n_21161;
wire n_15409;
wire n_4306;
wire n_18958;
wire n_3209;
wire n_3504;
wire n_19995;
wire n_1953;
wire n_2589;
wire n_7094;
wire n_16320;
wire n_10605;
wire n_8944;
wire n_21677;
wire n_12385;
wire n_17128;
wire n_537;
wire n_14937;
wire n_19699;
wire n_10464;
wire n_1504;
wire n_10034;
wire n_15130;
wire n_14249;
wire n_17884;
wire n_7790;
wire n_250;
wire n_3375;
wire n_12735;
wire n_12475;
wire n_260;
wire n_15375;
wire n_15461;
wire n_16186;
wire n_21020;
wire n_18636;
wire n_18340;
wire n_3167;
wire n_5558;
wire n_14022;
wire n_13800;
wire n_19883;
wire n_5350;
wire n_2362;
wire n_14105;
wire n_21154;
wire n_15120;
wire n_21790;
wire n_540;
wire n_8992;
wire n_13032;
wire n_19055;
wire n_11224;
wire n_20608;
wire n_10762;
wire n_10490;
wire n_14357;
wire n_894;
wire n_9078;
wire n_21037;
wire n_7207;
wire n_21368;
wire n_7454;
wire n_9012;
wire n_12794;
wire n_5830;
wire n_4812;
wire n_21399;
wire n_9233;
wire n_9217;
wire n_13576;
wire n_5760;
wire n_234;
wire n_18694;
wire n_20528;
wire n_15893;
wire n_1881;
wire n_2749;
wire n_17219;
wire n_3451;
wire n_8926;
wire n_4657;
wire n_2971;
wire n_14662;
wire n_2311;
wire n_5765;
wire n_14341;
wire n_6596;
wire n_14159;
wire n_5613;
wire n_4756;
wire n_5104;
wire n_4860;
wire n_4359;
wire n_21053;
wire n_20456;
wire n_20428;
wire n_20046;
wire n_19494;
wire n_10468;
wire n_12894;
wire n_10906;
wire n_4573;
wire n_19119;
wire n_5513;
wire n_12276;
wire n_15925;
wire n_4803;
wire n_19298;
wire n_12594;
wire n_10905;
wire n_7029;
wire n_13030;
wire n_2002;
wire n_5145;
wire n_12529;
wire n_21823;
wire n_2371;
wire n_6444;
wire n_6333;
wire n_13704;
wire n_5869;
wire n_5925;
wire n_749;
wire n_19220;
wire n_5359;
wire n_17325;
wire n_1134;
wire n_20730;
wire n_15427;
wire n_10361;
wire n_11269;
wire n_9955;
wire n_12402;
wire n_19998;
wire n_8921;
wire n_21493;
wire n_20309;
wire n_11314;
wire n_15359;
wire n_2016;
wire n_2711;
wire n_14963;
wire n_17035;
wire n_8286;
wire n_990;
wire n_2867;
wire n_9765;
wire n_1894;
wire n_975;
wire n_11130;
wire n_16530;
wire n_3124;
wire n_6737;
wire n_6454;
wire n_4253;
wire n_151;
wire n_14175;
wire n_19359;
wire n_15919;
wire n_770;
wire n_13656;
wire n_2852;
wire n_11035;
wire n_8925;
wire n_18556;
wire n_3100;
wire n_15986;
wire n_17740;
wire n_12901;
wire n_7505;
wire n_3758;
wire n_3356;
wire n_8047;
wire n_17875;
wire n_21899;
wire n_16658;
wire n_14562;
wire n_1736;
wire n_8268;
wire n_12564;
wire n_18989;
wire n_5858;
wire n_20840;
wire n_9840;
wire n_5723;
wire n_21602;
wire n_5295;
wire n_6137;
wire n_217;
wire n_4679;
wire n_12204;
wire n_6201;
wire n_7113;
wire n_20720;
wire n_14684;
wire n_2988;
wire n_21132;
wire n_15055;
wire n_15852;
wire n_21561;
wire n_11895;
wire n_15291;
wire n_7872;
wire n_1970;
wire n_13895;
wire n_12888;
wire n_4167;
wire n_8845;
wire n_19514;
wire n_12013;
wire n_17098;
wire n_21946;
wire n_5016;
wire n_20380;
wire n_12741;
wire n_8022;
wire n_3902;
wire n_4730;
wire n_7228;
wire n_15092;
wire n_19609;
wire n_19155;
wire n_6380;
wire n_9091;
wire n_18290;
wire n_5996;
wire n_11977;
wire n_2232;
wire n_19852;
wire n_11215;
wire n_9932;
wire n_15274;
wire n_1774;
wire n_19933;
wire n_15814;
wire n_13726;
wire n_11530;
wire n_7702;
wire n_9542;
wire n_15000;
wire n_12889;
wire n_15765;
wire n_17862;
wire n_17669;
wire n_8791;
wire n_4204;
wire n_6772;
wire n_6823;
wire n_732;
wire n_5906;
wire n_20459;
wire n_16036;
wire n_20118;
wire n_16944;
wire n_14549;
wire n_3825;
wire n_21479;
wire n_8048;
wire n_15058;
wire n_20155;
wire n_10802;
wire n_2008;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_19129;
wire n_18515;
wire n_1213;
wire n_13280;
wire n_20476;
wire n_19653;
wire n_3792;
wire n_8506;
wire n_11289;
wire n_8465;
wire n_16433;
wire n_12277;
wire n_4269;
wire n_4695;
wire n_5736;
wire n_3312;
wire n_1352;
wire n_12250;
wire n_5069;
wire n_10574;
wire n_6543;
wire n_16480;
wire n_20145;
wire n_11622;
wire n_19152;
wire n_11763;
wire n_20970;
wire n_5052;
wire n_6091;
wire n_664;
wire n_10155;
wire n_16930;
wire n_14585;
wire n_21416;
wire n_15964;
wire n_9751;
wire n_14866;
wire n_916;
wire n_13134;
wire n_13399;
wire n_7085;
wire n_20242;
wire n_9579;
wire n_3606;
wire n_6652;
wire n_18974;
wire n_5004;
wire n_8366;
wire n_16137;
wire n_20298;
wire n_8101;
wire n_14065;
wire n_18181;
wire n_17198;
wire n_19586;
wire n_5880;
wire n_15082;
wire n_12211;
wire n_17162;
wire n_5713;
wire n_1683;
wire n_10212;
wire n_17528;
wire n_8052;
wire n_997;
wire n_19314;
wire n_11143;
wire n_18674;
wire n_9729;
wire n_5105;
wire n_15367;
wire n_18438;
wire n_13886;
wire n_15934;
wire n_1268;
wire n_17855;
wire n_7856;
wire n_4050;
wire n_17320;
wire n_15250;
wire n_5623;
wire n_10005;
wire n_17433;
wire n_17760;
wire n_14798;
wire n_981;
wire n_18680;
wire n_7399;
wire n_867;
wire n_19166;
wire n_2422;
wire n_5256;
wire n_21797;
wire n_12545;
wire n_11621;
wire n_6814;
wire n_16943;
wire n_2057;
wire n_9825;
wire n_10093;
wire n_18231;
wire n_905;
wire n_17377;
wire n_7472;
wire n_10850;
wire n_8371;
wire n_5872;
wire n_18688;
wire n_15984;
wire n_3858;
wire n_8231;
wire n_4502;
wire n_20669;
wire n_20475;
wire n_4851;
wire n_5735;
wire n_12119;
wire n_21942;
wire n_8164;
wire n_6944;
wire n_7384;
wire n_14280;
wire n_3081;
wire n_3313;
wire n_8870;
wire n_6193;
wire n_10614;
wire n_20432;
wire n_934;
wire n_8422;
wire n_1618;
wire n_12094;
wire n_12730;
wire n_5049;
wire n_6757;
wire n_19351;
wire n_654;
wire n_5953;
wire n_2726;
wire n_20116;
wire n_4723;
wire n_5176;
wire n_6779;
wire n_17772;
wire n_14094;
wire n_7938;
wire n_8253;
wire n_12534;
wire n_5820;
wire n_9028;
wire n_14722;
wire n_2456;
wire n_2678;
wire n_11383;
wire n_16386;
wire n_16168;
wire n_2451;
wire n_11655;
wire n_12553;
wire n_7812;
wire n_5051;
wire n_930;
wire n_181;
wire n_9724;
wire n_8292;
wire n_21499;
wire n_2854;
wire n_1701;
wire n_18113;
wire n_8611;
wire n_19390;
wire n_20335;
wire n_682;
wire n_9826;
wire n_19391;
wire n_4153;
wire n_13118;
wire n_15271;
wire n_20394;
wire n_839;
wire n_2964;
wire n_12283;
wire n_17672;
wire n_4530;
wire n_8123;
wire n_2292;
wire n_3865;
wire n_7092;
wire n_6971;
wire n_9938;
wire n_21672;
wire n_8424;
wire n_9776;
wire n_8859;
wire n_21473;
wire n_16539;
wire n_11914;
wire n_19447;
wire n_3428;
wire n_17829;
wire n_2961;
wire n_9212;
wire n_13431;
wire n_236;
wire n_1396;
wire n_1752;
wire n_21157;
wire n_13082;
wire n_7904;
wire n_21411;
wire n_4182;
wire n_12683;
wire n_12108;
wire n_15267;
wire n_20644;
wire n_5120;
wire n_17135;
wire n_11625;
wire n_10416;
wire n_18401;
wire n_21809;
wire n_14933;
wire n_7922;
wire n_8618;
wire n_11787;
wire n_14024;
wire n_8285;
wire n_15790;
wire n_10396;
wire n_12899;
wire n_14252;
wire n_10123;
wire n_5772;
wire n_474;
wire n_3575;
wire n_17898;
wire n_6964;
wire n_20835;
wire n_6202;
wire n_11364;
wire n_12713;
wire n_9445;
wire n_18261;
wire n_4097;
wire n_14031;
wire n_13089;
wire n_5392;
wire n_9930;
wire n_17278;
wire n_19946;
wire n_15755;
wire n_17038;
wire n_21007;
wire n_12757;
wire n_7371;
wire n_6962;
wire n_17783;
wire n_10347;
wire n_6455;
wire n_9727;
wire n_4273;
wire n_3024;
wire n_18159;
wire n_15895;
wire n_13879;
wire n_16975;
wire n_6644;
wire n_13848;
wire n_14633;
wire n_14475;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_6160;
wire n_11486;
wire n_1540;
wire n_10650;
wire n_11777;
wire n_6031;
wire n_720;
wire n_2500;
wire n_7653;
wire n_20894;
wire n_5656;
wire n_863;
wire n_8531;
wire n_20956;
wire n_2695;
wire n_3480;
wire n_6280;
wire n_11941;
wire n_10048;
wire n_15372;
wire n_3662;
wire n_7383;
wire n_18031;
wire n_9396;
wire n_17504;
wire n_9234;
wire n_10364;
wire n_17402;
wire n_5752;
wire n_17824;
wire n_4726;
wire n_1879;
wire n_4222;
wire n_8341;
wire n_19842;
wire n_20431;
wire n_13995;
wire n_16263;
wire n_2274;
wire n_8521;
wire n_811;
wire n_6077;
wire n_11718;
wire n_4119;
wire n_7743;
wire n_17407;
wire n_14128;
wire n_12762;
wire n_5217;
wire n_1004;
wire n_242;
wire n_1681;
wire n_10502;
wire n_2975;
wire n_5029;
wire n_19350;
wire n_16377;
wire n_19302;
wire n_10674;
wire n_16721;
wire n_4884;
wire n_21612;
wire n_4009;
wire n_19929;
wire n_16273;
wire n_4580;
wire n_6792;
wire n_1263;
wire n_12980;
wire n_4999;
wire n_18237;
wire n_11418;
wire n_20078;
wire n_13795;
wire n_4112;
wire n_18994;
wire n_17018;
wire n_4337;
wire n_18118;
wire n_14052;
wire n_16562;
wire n_552;
wire n_5335;
wire n_12650;
wire n_20787;
wire n_7300;
wire n_423;
wire n_9566;
wire n_18928;
wire n_19131;
wire n_17426;
wire n_8483;
wire n_14820;
wire n_5960;
wire n_8605;
wire n_18014;
wire n_14778;
wire n_5002;
wire n_11750;
wire n_11038;
wire n_13363;
wire n_19193;
wire n_1947;
wire n_2114;
wire n_19813;
wire n_11894;
wire n_16305;
wire n_13689;
wire n_8374;
wire n_19323;
wire n_4635;
wire n_7118;
wire n_8006;
wire n_6285;
wire n_8723;
wire n_6025;
wire n_18695;
wire n_10944;
wire n_19885;
wire n_16999;
wire n_15809;
wire n_2543;
wire n_19026;
wire n_10140;
wire n_10013;
wire n_3180;
wire n_13909;
wire n_16234;
wire n_8220;
wire n_1705;
wire n_20224;
wire n_11356;
wire n_19414;
wire n_3107;
wire n_13045;
wire n_7910;
wire n_1261;
wire n_4955;
wire n_15985;
wire n_20066;
wire n_14147;
wire n_9394;
wire n_3650;
wire n_8991;
wire n_6343;
wire n_10186;
wire n_11938;
wire n_15505;
wire n_16404;
wire n_18205;
wire n_21885;
wire n_6049;
wire n_2515;
wire n_2466;
wire n_6052;
wire n_17565;
wire n_11412;
wire n_13522;
wire n_10700;
wire n_4197;
wire n_21941;
wire n_7069;
wire n_13208;
wire n_1949;
wire n_1946;
wire n_14219;
wire n_12169;
wire n_11249;
wire n_12838;
wire n_775;
wire n_19395;
wire n_13847;
wire n_15006;
wire n_13559;
wire n_10758;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_7252;
wire n_20723;
wire n_20987;
wire n_15450;
wire n_1831;
wire n_4394;
wire n_9051;
wire n_7133;
wire n_21287;
wire n_10345;
wire n_243;
wire n_12809;
wire n_9908;
wire n_12748;
wire n_13639;
wire n_350;
wire n_7061;
wire n_17516;
wire n_15297;
wire n_4065;
wire n_19263;
wire n_8660;
wire n_5187;
wire n_18202;
wire n_21639;
wire n_7216;
wire n_6601;
wire n_475;
wire n_9687;
wire n_20651;
wire n_11984;
wire n_6839;
wire n_13053;
wire n_9519;
wire n_7711;
wire n_958;
wire n_15431;
wire n_18471;
wire n_12137;
wire n_3744;
wire n_17569;
wire n_11651;
wire n_21231;
wire n_6051;
wire n_4716;
wire n_18445;
wire n_19045;
wire n_164;
wire n_2432;
wire n_7972;
wire n_1521;
wire n_21518;
wire n_17602;
wire n_6532;
wire n_13517;
wire n_214;
wire n_18759;
wire n_17817;
wire n_12644;
wire n_7458;
wire n_7614;
wire n_20541;
wire n_2337;
wire n_17422;
wire n_19913;
wire n_11696;
wire n_3907;
wire n_16730;
wire n_6526;
wire n_8142;
wire n_13455;
wire n_17451;
wire n_2932;
wire n_17424;
wire n_18368;
wire n_2980;
wire n_5225;
wire n_1784;
wire n_16061;
wire n_14213;
wire n_10447;
wire n_10022;
wire n_18263;
wire n_5265;
wire n_10305;
wire n_14769;
wire n_15777;
wire n_460;
wire n_16880;
wire n_21505;
wire n_12877;
wire n_4753;
wire n_19820;
wire n_18882;
wire n_3885;
wire n_9405;
wire n_19321;
wire n_13892;
wire n_19941;
wire n_13636;
wire n_16489;
wire n_14317;
wire n_16866;
wire n_5574;
wire n_20049;
wire n_18508;
wire n_20112;
wire n_16272;
wire n_1039;
wire n_6508;
wire n_15820;
wire n_11116;
wire n_16346;
wire n_3320;
wire n_7052;
wire n_5009;
wire n_21064;
wire n_2688;
wire n_17793;
wire n_10510;
wire n_13934;
wire n_13905;
wire n_13240;
wire n_15915;
wire n_17097;
wire n_21253;
wire n_18032;
wire n_10993;
wire n_15353;
wire n_14132;
wire n_21341;
wire n_16918;
wire n_12844;
wire n_4375;
wire n_13868;
wire n_9902;
wire n_16430;
wire n_17537;
wire n_9621;
wire n_21237;
wire n_9604;
wire n_3580;
wire n_18144;
wire n_4609;
wire n_20278;
wire n_9821;
wire n_5876;
wire n_19126;
wire n_17042;
wire n_12076;
wire n_6704;
wire n_6409;
wire n_1565;
wire n_4088;
wire n_6876;
wire n_1809;
wire n_19523;
wire n_21478;
wire n_5540;
wire n_19752;
wire n_3305;
wire n_15784;
wire n_4148;
wire n_20859;
wire n_12702;
wire n_18879;
wire n_6938;
wire n_12050;
wire n_4373;
wire n_14577;
wire n_4934;
wire n_9952;
wire n_12473;
wire n_20819;
wire n_4475;
wire n_3989;
wire n_10076;
wire n_3804;
wire n_8168;
wire n_1775;
wire n_14837;
wire n_17043;
wire n_7038;
wire n_4683;
wire n_728;
wire n_272;
wire n_13649;
wire n_12956;
wire n_18145;
wire n_2603;
wire n_11203;
wire n_18314;
wire n_9447;
wire n_1905;
wire n_18190;
wire n_2195;
wire n_20300;
wire n_9592;
wire n_14111;
wire n_931;
wire n_11416;
wire n_17398;
wire n_1544;
wire n_11809;
wire n_15187;
wire n_19277;
wire n_1629;
wire n_12038;
wire n_5901;
wire n_21298;
wire n_16989;
wire n_14359;
wire n_17530;
wire n_21729;
wire n_17513;
wire n_21228;
wire n_4905;
wire n_17733;
wire n_360;
wire n_19255;
wire n_19831;
wire n_10772;
wire n_21779;
wire n_16895;
wire n_4278;
wire n_1635;
wire n_13184;
wire n_15641;
wire n_4910;
wire n_15330;
wire n_12297;
wire n_9874;
wire n_7392;
wire n_2215;
wire n_8245;
wire n_6239;
wire n_706;
wire n_15050;
wire n_3978;
wire n_14281;
wire n_7583;
wire n_14876;
wire n_4809;
wire n_5226;
wire n_7657;
wire n_1925;
wire n_5867;
wire n_13318;
wire n_5590;
wire n_14515;
wire n_8390;
wire n_15252;
wire n_11480;
wire n_11874;
wire n_12115;
wire n_1415;
wire n_19711;
wire n_2592;
wire n_15324;
wire n_2838;
wire n_3133;
wire n_10181;
wire n_17988;
wire n_11862;
wire n_3725;
wire n_4972;
wire n_18299;
wire n_3128;
wire n_18077;
wire n_15496;
wire n_14370;
wire n_7896;
wire n_2178;
wire n_19559;
wire n_10481;
wire n_7176;
wire n_14194;
wire n_15770;
wire n_10220;
wire n_13917;
wire n_17324;
wire n_5625;
wire n_9218;
wire n_20354;
wire n_21955;
wire n_10634;
wire n_3942;
wire n_2736;
wire n_14489;
wire n_21566;
wire n_15321;
wire n_7826;
wire n_3000;
wire n_252;
wire n_20828;
wire n_3108;
wire n_3111;
wire n_1837;
wire n_5646;
wire n_18538;
wire n_21317;
wire n_9164;
wire n_3844;
wire n_4054;
wire n_5448;
wire n_20878;
wire n_13732;
wire n_259;
wire n_448;
wire n_11985;
wire n_3003;
wire n_6995;
wire n_7185;
wire n_1158;
wire n_6254;
wire n_11020;
wire n_15233;
wire n_18112;
wire n_8134;
wire n_14542;
wire n_8694;
wire n_8965;
wire n_13288;
wire n_17704;
wire n_908;
wire n_15350;
wire n_6128;
wire n_11587;
wire n_17046;
wire n_2084;
wire n_5749;
wire n_11697;
wire n_8427;
wire n_20804;
wire n_16554;
wire n_5108;
wire n_959;
wire n_9156;
wire n_14591;
wire n_16832;
wire n_19146;
wire n_11435;
wire n_3243;
wire n_21617;
wire n_16765;
wire n_1169;
wire n_13236;
wire n_6848;
wire n_15590;
wire n_8345;
wire n_10414;
wire n_9708;
wire n_11644;
wire n_17165;
wire n_20065;
wire n_20485;
wire n_17498;
wire n_1640;
wire n_7775;
wire n_2162;
wire n_21825;
wire n_2051;
wire n_19519;
wire n_5072;
wire n_3629;
wire n_17667;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_20646;
wire n_9473;
wire n_1171;
wire n_12341;
wire n_20400;
wire n_8038;
wire n_15525;
wire n_8949;
wire n_14248;
wire n_19410;
wire n_14928;
wire n_10612;
wire n_5619;
wire n_2048;
wire n_9244;
wire n_14878;
wire n_9584;
wire n_1921;
wire n_10797;
wire n_13320;
wire n_9439;
wire n_11915;
wire n_355;
wire n_20464;
wire n_8655;
wire n_1286;
wire n_3276;
wire n_6728;
wire n_18567;
wire n_15313;
wire n_17430;
wire n_9768;
wire n_18788;
wire n_8777;
wire n_6133;
wire n_14951;
wire n_8852;
wire n_20185;
wire n_10114;
wire n_613;
wire n_7407;
wire n_1119;
wire n_1240;
wire n_21917;
wire n_8185;
wire n_19761;
wire n_2519;
wire n_8513;
wire n_6670;
wire n_20454;
wire n_8365;
wire n_14229;
wire n_361;
wire n_17562;
wire n_6038;
wire n_19648;
wire n_4818;
wire n_20930;
wire n_19985;
wire n_10599;
wire n_4514;
wire n_4800;
wire n_3960;
wire n_9836;
wire n_2277;
wire n_18217;
wire n_8035;
wire n_11399;
wire n_18824;
wire n_8874;
wire n_11542;
wire n_2474;
wire n_7334;
wire n_10623;
wire n_1591;
wire n_2033;
wire n_7755;
wire n_19142;
wire n_4341;
wire n_9187;
wire n_1682;
wire n_11276;
wire n_4312;
wire n_2628;
wire n_10511;
wire n_1249;
wire n_1111;
wire n_15180;
wire n_18472;
wire n_9406;
wire n_13604;
wire n_9342;
wire n_1909;
wire n_14119;
wire n_4277;
wire n_13323;
wire n_14321;
wire n_19606;
wire n_18087;
wire n_17678;
wire n_14808;
wire n_16946;
wire n_18139;
wire n_19627;
wire n_12755;
wire n_8644;
wire n_12306;
wire n_10516;
wire n_20564;
wire n_3779;
wire n_18999;
wire n_19722;
wire n_7200;
wire n_13068;
wire n_1456;
wire n_9860;
wire n_18924;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_3037;
wire n_18709;
wire n_16938;
wire n_17547;
wire n_10548;
wire n_6743;
wire n_10547;
wire n_2176;
wire n_1816;
wire n_14011;
wire n_13958;
wire n_19650;
wire n_12603;
wire n_14230;
wire n_15907;
wire n_2455;
wire n_7877;
wire n_1849;
wire n_8945;
wire n_1131;
wire n_11857;
wire n_15886;
wire n_5631;
wire n_8028;
wire n_21135;
wire n_7243;
wire n_20619;
wire n_4063;
wire n_11193;
wire n_6617;
wire n_1209;
wire n_602;
wire n_4888;
wire n_21958;
wire n_4874;
wire n_7608;
wire n_3793;
wire n_4669;
wire n_19585;
wire n_12244;
wire n_16971;
wire n_13851;
wire n_14209;
wire n_4060;
wire n_996;
wire n_1717;
wire n_14177;
wire n_2128;
wire n_18186;
wire n_21352;
wire n_327;
wire n_21865;
wire n_14485;
wire n_18704;
wire n_1438;
wire n_7373;
wire n_20129;
wire n_2534;
wire n_15009;
wire n_6186;
wire n_5153;
wire n_16574;
wire n_21311;
wire n_2198;
wire n_11285;
wire n_12618;
wire n_20818;
wire n_11513;
wire n_1424;
wire n_16142;
wire n_4266;
wire n_11250;
wire n_7874;
wire n_15992;
wire n_11340;
wire n_19186;
wire n_199;
wire n_4248;
wire n_5915;
wire n_5452;
wire n_7226;
wire n_8930;
wire n_20151;
wire n_18015;
wire n_6609;
wire n_20237;
wire n_19803;
wire n_13592;
wire n_18630;
wire n_3548;
wire n_418;
wire n_19548;
wire n_8405;
wire n_14558;
wire n_7913;
wire n_4383;
wire n_397;
wire n_5535;
wire n_17453;
wire n_20972;
wire n_3875;
wire n_15598;
wire n_13967;
wire n_7891;
wire n_6391;
wire n_20408;
wire n_8088;
wire n_5299;
wire n_20281;
wire n_4586;
wire n_4048;
wire n_1844;
wire n_13546;
wire n_20964;
wire n_13978;
wire n_11771;
wire n_4784;
wire n_17224;
wire n_18177;
wire n_7203;
wire n_9757;
wire n_15121;
wire n_18995;
wire n_2999;
wire n_18583;
wire n_5082;
wire n_2086;
wire n_5209;
wire n_7215;
wire n_10246;
wire n_16146;
wire n_16662;
wire n_20985;
wire n_15347;
wire n_14295;
wire n_21931;
wire n_1179;
wire n_753;
wire n_11185;
wire n_18572;
wire n_11498;
wire n_10299;
wire n_330;
wire n_20153;
wire n_692;
wire n_18757;
wire n_20499;
wire n_1911;
wire n_15494;
wire n_20557;
wire n_5868;
wire n_6538;
wire n_17517;
wire n_15946;
wire n_1688;
wire n_6633;
wire n_9371;
wire n_15662;
wire n_6172;
wire n_18273;
wire n_5275;
wire n_10702;
wire n_4689;
wire n_20534;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_11768;
wire n_17385;
wire n_21075;
wire n_17173;
wire n_14748;
wire n_20699;
wire n_6574;
wire n_11683;
wire n_9484;
wire n_7996;
wire n_449;
wire n_20926;
wire n_1400;
wire n_1342;
wire n_8588;
wire n_20852;
wire n_3574;
wire n_19011;
wire n_16564;
wire n_4201;
wire n_10366;
wire n_12207;
wire n_14168;
wire n_896;
wire n_17754;
wire n_6766;
wire n_356;
wire n_20294;
wire n_1730;
wire n_14575;
wire n_4123;
wire n_6330;
wire n_5520;
wire n_8896;
wire n_14695;
wire n_964;
wire n_16706;
wire n_4479;
wire n_17462;
wire n_19851;
wire n_9452;
wire n_16771;
wire n_1307;
wire n_3372;
wire n_814;
wire n_17085;
wire n_9974;
wire n_15221;
wire n_5920;
wire n_17030;
wire n_8256;
wire n_14578;
wire n_14003;
wire n_17710;
wire n_15692;
wire n_17336;
wire n_7916;
wire n_6450;
wire n_16990;
wire n_17665;
wire n_1204;
wire n_13776;
wire n_21496;
wire n_12878;
wire n_4690;
wire n_10174;
wire n_12879;
wire n_3780;
wire n_783;
wire n_12601;
wire n_6775;
wire n_5274;
wire n_18564;
wire n_10873;
wire n_3848;
wire n_4284;
wire n_11582;
wire n_20356;
wire n_8207;
wire n_3919;
wire n_13688;
wire n_6445;
wire n_19952;
wire n_19806;
wire n_20341;
wire n_510;
wire n_16922;
wire n_17341;
wire n_9615;
wire n_4053;
wire n_7759;
wire n_11180;
wire n_21515;
wire n_9945;
wire n_15574;
wire n_5587;
wire n_6855;
wire n_2444;
wire n_5789;
wire n_8217;
wire n_241;
wire n_13911;
wire n_6585;
wire n_19491;
wire n_13124;
wire n_10659;
wire n_866;
wire n_9295;
wire n_18746;
wire n_6252;
wire n_20253;
wire n_10239;
wire n_577;
wire n_4005;
wire n_1687;
wire n_11630;
wire n_8051;
wire n_3578;
wire n_3812;
wire n_20353;
wire n_14303;
wire n_15998;
wire n_17346;
wire n_15714;
wire n_7757;
wire n_5865;
wire n_13019;
wire n_1375;
wire n_15275;
wire n_17811;
wire n_14848;
wire n_3774;
wire n_14989;
wire n_19811;
wire n_10276;
wire n_3093;
wire n_15332;
wire n_12533;
wire n_7138;
wire n_8544;
wire n_21345;
wire n_2431;
wire n_9789;
wire n_9299;
wire n_7284;
wire n_14693;
wire n_1190;
wire n_18861;
wire n_17596;
wire n_12573;
wire n_15047;
wire n_966;
wire n_14839;
wire n_5786;
wire n_4987;
wire n_11113;
wire n_1212;
wire n_2074;
wire n_19073;
wire n_21461;
wire n_19836;
wire n_20521;
wire n_2217;
wire n_13116;
wire n_5658;
wire n_899;
wire n_18740;
wire n_13968;
wire n_4823;
wire n_17003;
wire n_9427;
wire n_1628;
wire n_19748;
wire n_20381;
wire n_8698;
wire n_19638;
wire n_12530;
wire n_13718;
wire n_15671;
wire n_1005;
wire n_607;
wire n_2437;
wire n_20620;
wire n_6813;
wire n_5564;
wire n_2445;
wire n_17485;
wire n_1835;
wire n_7644;
wire n_12494;
wire n_1853;
wire n_13147;
wire n_8986;
wire n_11905;
wire n_12488;
wire n_19064;
wire n_4529;
wire n_12229;
wire n_3034;
wire n_8200;
wire n_19492;
wire n_20387;
wire n_8528;
wire n_529;
wire n_17749;
wire n_10764;
wire n_16894;
wire n_16177;
wire n_14333;
wire n_19639;
wire n_202;
wire n_15490;
wire n_19890;
wire n_791;
wire n_3467;
wire n_8267;
wire n_2830;
wire n_4354;
wire n_4653;
wire n_17507;
wire n_21394;
wire n_16042;
wire n_9734;
wire n_9505;
wire n_2246;
wire n_7199;
wire n_17527;
wire n_3901;
wire n_715;
wire n_18270;
wire n_14085;
wire n_16932;
wire n_18056;
wire n_21251;
wire n_19433;
wire n_12946;
wire n_13397;
wire n_17214;
wire n_10707;
wire n_12613;
wire n_13882;
wire n_21120;
wire n_17423;
wire n_9336;
wire n_9360;
wire n_21611;
wire n_18490;
wire n_6024;
wire n_7866;
wire n_18172;
wire n_13252;
wire n_18317;
wire n_2814;
wire n_15553;
wire n_17784;
wire n_3826;
wire n_12978;
wire n_2211;
wire n_7638;
wire n_20366;
wire n_14857;
wire n_7988;
wire n_3337;
wire n_855;
wire n_3204;
wire n_7259;
wire n_13050;
wire n_2136;
wire n_13384;
wire n_12289;
wire n_1273;
wire n_10862;
wire n_21296;
wire n_18397;
wire n_5157;
wire n_980;
wire n_698;
wire n_20397;
wire n_1282;
wire n_3043;
wire n_19213;
wire n_998;
wire n_12596;
wire n_9478;
wire n_4880;
wire n_9266;
wire n_9813;
wire n_19818;
wire n_501;
wire n_3892;
wire n_1417;
wire n_5061;
wire n_5572;
wire n_20276;
wire n_11573;
wire n_11703;
wire n_11671;
wire n_7576;
wire n_21943;
wire n_19173;
wire n_6795;
wire n_18403;
wire n_20936;
wire n_21098;
wire n_21041;
wire n_16090;
wire n_20133;
wire n_4193;
wire n_5873;
wire n_9666;
wire n_10112;
wire n_15200;
wire n_7734;
wire n_18271;
wire n_15046;
wire n_3647;
wire n_10056;
wire n_15680;
wire n_506;
wire n_737;
wire n_19596;
wire n_17277;
wire n_17722;
wire n_3609;
wire n_15498;
wire n_12423;
wire n_18241;
wire n_10105;
wire n_13008;
wire n_16577;
wire n_6663;
wire n_20570;
wire n_20371;
wire n_15022;
wire n_3959;
wire n_7327;
wire n_18084;
wire n_5763;
wire n_18442;
wire n_9987;
wire n_20383;
wire n_8124;
wire n_20871;
wire n_12518;
wire n_15519;
wire n_12764;
wire n_5246;
wire n_5964;
wire n_11065;
wire n_13812;
wire n_13751;
wire n_15143;
wire n_11447;
wire n_12427;
wire n_17908;
wire n_14217;
wire n_4592;
wire n_16700;
wire n_3069;
wire n_18921;
wire n_20032;
wire n_1900;
wire n_20074;
wire n_11676;
wire n_11319;
wire n_8478;
wire n_6075;
wire n_7082;
wire n_9569;
wire n_18030;
wire n_13513;
wire n_2735;
wire n_2497;
wire n_15808;
wire n_11018;
wire n_18212;
wire n_9707;
wire n_19530;
wire n_14664;
wire n_13858;
wire n_2014;
wire n_11537;
wire n_19814;
wire n_8996;
wire n_15949;
wire n_16112;
wire n_4828;
wire n_9797;
wire n_17713;
wire n_19739;
wire n_9053;
wire n_6478;
wire n_6066;
wire n_19692;
wire n_12437;
wire n_7034;
wire n_21564;
wire n_20438;
wire n_8303;
wire n_3626;
wire n_19859;
wire n_13859;
wire n_10661;
wire n_12026;
wire n_16442;
wire n_9089;
wire n_10505;
wire n_21680;
wire n_21619;
wire n_3908;
wire n_6175;
wire n_15387;
wire n_2423;
wire n_3671;
wire n_17687;
wire n_9493;
wire n_14364;
wire n_6410;
wire n_12607;
wire n_12958;
wire n_16185;
wire n_21904;
wire n_3302;
wire n_17143;
wire n_20453;
wire n_15713;
wire n_8914;
wire n_5162;
wire n_8520;
wire n_3842;
wire n_18780;
wire n_16991;
wire n_4482;
wire n_2041;
wire n_631;
wire n_14780;
wire n_1797;
wire n_9119;
wire n_11903;
wire n_12226;
wire n_8682;
wire n_7331;
wire n_8775;
wire n_18681;
wire n_11476;
wire n_8696;
wire n_16002;
wire n_6957;
wire n_7514;
wire n_11966;
wire n_20531;
wire n_11115;
wire n_17186;
wire n_15113;
wire n_17354;
wire n_5946;
wire n_2744;
wire n_6711;
wire n_7445;
wire n_6847;
wire n_21086;
wire n_9131;
wire n_10522;
wire n_11200;
wire n_16072;
wire n_10752;
wire n_15426;
wire n_6384;
wire n_333;
wire n_1298;
wire n_1652;
wire n_10768;
wire n_16806;
wire n_258;
wire n_15352;
wire n_6298;
wire n_11170;
wire n_11337;
wire n_13987;
wire n_17300;
wire n_9032;
wire n_14982;
wire n_188;
wire n_7361;
wire n_12929;
wire n_8890;
wire n_16979;
wire n_5710;
wire n_7453;
wire n_463;
wire n_14010;
wire n_5566;
wire n_19845;
wire n_19175;
wire n_20590;
wire n_2438;
wire n_465;
wire n_17487;
wire n_2296;
wire n_20372;
wire n_13988;
wire n_3181;
wire n_2278;
wire n_10412;
wire n_5450;
wire n_6834;
wire n_20703;
wire n_11975;
wire n_5313;
wire n_13073;
wire n_20858;
wire n_9374;
wire n_20033;
wire n_21178;
wire n_6723;
wire n_14008;
wire n_1408;
wire n_494;
wire n_12763;
wire n_14597;
wire n_11402;
wire n_8342;
wire n_17985;
wire n_15549;
wire n_795;
wire n_5188;
wire n_180;
wire n_3281;
wire n_6078;
wire n_8571;
wire n_9308;
wire n_20264;
wire n_4318;
wire n_10721;
wire n_20477;
wire n_20763;
wire n_7921;
wire n_8877;
wire n_16247;
wire n_8862;
wire n_4797;
wire n_10823;
wire n_1526;
wire n_10176;
wire n_1275;
wire n_20744;
wire n_7538;
wire n_712;
wire n_11778;
wire n_17343;
wire n_1042;
wire n_7077;
wire n_21889;
wire n_12561;
wire n_19594;
wire n_13382;
wire n_20626;
wire n_15528;
wire n_4124;
wire n_15276;
wire n_17093;
wire n_4994;
wire n_13353;
wire n_4245;
wire n_4364;
wire n_2383;
wire n_597;
wire n_3406;
wire n_16158;
wire n_9847;
wire n_20957;
wire n_19488;
wire n_10227;
wire n_11096;
wire n_17554;
wire n_1558;
wire n_8805;
wire n_18652;
wire n_1704;
wire n_15219;
wire n_3721;
wire n_12635;
wire n_6507;
wire n_20640;
wire n_2013;
wire n_14819;
wire n_1032;
wire n_15137;
wire n_2991;
wire n_10409;
wire n_2752;
wire n_19191;
wire n_10709;
wire n_21324;
wire n_18845;
wire n_3699;
wire n_13047;
wire n_13049;
wire n_3360;
wire n_18208;
wire n_15668;
wire n_16735;
wire n_17968;
wire n_8111;
wire n_13903;
wire n_9194;
wire n_3241;
wire n_6546;
wire n_13683;
wire n_9655;
wire n_18728;
wire n_2899;
wire n_790;
wire n_18706;
wire n_3541;
wire n_3622;
wire n_11326;
wire n_19017;
wire n_14036;
wire n_13241;
wire n_13217;
wire n_16007;
wire n_13927;
wire n_18151;
wire n_7303;
wire n_13112;
wire n_9083;
wire n_16276;
wire n_14631;
wire n_17821;
wire n_13779;
wire n_8383;
wire n_5035;
wire n_21429;
wire n_1960;
wire n_11583;
wire n_551;
wire n_13499;
wire n_20363;
wire n_1466;
wire n_14203;
wire n_13768;
wire n_3202;
wire n_8002;
wire n_18648;
wire n_4977;
wire n_8594;
wire n_6276;
wire n_18858;
wire n_6072;
wire n_3587;
wire n_5033;
wire n_10883;
wire n_7686;
wire n_4211;
wire n_16152;
wire n_12328;
wire n_8603;
wire n_12493;
wire n_6742;
wire n_9769;
wire n_16454;
wire n_15411;
wire n_3776;
wire n_7616;
wire n_2530;
wire n_2483;
wire n_4950;
wire n_11450;
wire n_8244;
wire n_16963;
wire n_1107;
wire n_2076;
wire n_6580;
wire n_17857;
wire n_18550;
wire n_17895;
wire n_21765;
wire n_21791;
wire n_17947;
wire n_19150;
wire n_2147;
wire n_16013;
wire n_19001;
wire n_11801;
wire n_14435;
wire n_13415;
wire n_4131;
wire n_18152;
wire n_2584;
wire n_5851;
wire n_21605;
wire n_15797;
wire n_3082;
wire n_2189;
wire n_1242;
wire n_9363;
wire n_13906;
wire n_12012;
wire n_12462;
wire n_5744;
wire n_18713;
wire n_17526;
wire n_11947;
wire n_14411;
wire n_281;
wire n_4499;
wire n_8413;
wire n_731;
wire n_5648;
wire n_13748;
wire n_18100;
wire n_7667;
wire n_1512;
wire n_6931;
wire n_1490;
wire n_17833;
wire n_9811;
wire n_12970;
wire n_6618;
wire n_18942;
wire n_4311;
wire n_5922;
wire n_12100;
wire n_1449;
wire n_20274;
wire n_15990;
wire n_15484;
wire n_18109;
wire n_10399;
wire n_21402;
wire n_219;
wire n_157;
wire n_17124;
wire n_20435;
wire n_20989;
wire n_12819;
wire n_7421;
wire n_14403;
wire n_16311;
wire n_3183;
wire n_8089;
wire n_13401;
wire n_19344;
wire n_4203;
wire n_9382;
wire n_16558;
wire n_16275;
wire n_3376;
wire n_15256;
wire n_11497;
wire n_5037;
wire n_16598;
wire n_11541;
wire n_8885;
wire n_3653;
wire n_10437;
wire n_10430;
wire n_4976;
wire n_2648;
wire n_10177;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_18431;
wire n_2439;
wire n_4811;
wire n_6096;
wire n_12767;
wire n_1165;
wire n_12754;
wire n_5144;
wire n_1034;
wire n_9422;
wire n_16942;
wire n_14892;
wire n_21278;
wire n_4758;
wire n_16326;
wire n_9795;
wire n_8380;
wire n_845;
wire n_528;
wire n_5577;
wire n_395;
wire n_7592;
wire n_15697;
wire n_3668;
wire n_21004;
wire n_14579;
wire n_15312;
wire n_6512;
wire n_11272;
wire n_13096;
wire n_2934;
wire n_3550;
wire n_15154;
wire n_1626;
wire n_1405;
wire n_12101;
wire n_13753;
wire n_10316;
wire n_9033;
wire n_20572;
wire n_21816;
wire n_7613;
wire n_16683;
wire n_9429;
wire n_3395;
wire n_12576;
wire n_17265;
wire n_7083;
wire n_4917;
wire n_13610;
wire n_16687;
wire n_15343;
wire n_6464;
wire n_2863;
wire n_11962;
wire n_5825;
wire n_1585;
wire n_6820;
wire n_1599;
wire n_12237;
wire n_18531;
wire n_17230;
wire n_16876;
wire n_2730;
wire n_21925;
wire n_2251;
wire n_6561;
wire n_21468;
wire n_18504;
wire n_4532;
wire n_3339;
wire n_228;
wire n_3735;
wire n_14605;
wire n_2248;
wire n_17998;
wire n_19706;
wire n_3007;
wire n_6769;
wire n_21957;
wire n_13131;
wire n_6592;
wire n_11150;
wire n_5686;
wire n_2622;
wire n_12298;
wire n_5463;
wire n_310;
wire n_12299;
wire n_2258;
wire n_9625;
wire n_10980;
wire n_279;
wire n_1014;
wire n_12232;
wire n_19884;
wire n_8064;
wire n_18604;
wire n_19439;
wire n_15564;
wire n_2140;
wire n_9694;
wire n_19881;
wire n_20656;
wire n_15544;
wire n_17427;
wire n_16341;
wire n_19740;
wire n_7701;
wire n_3611;
wire n_2862;
wire n_18081;
wire n_19227;
wire n_8214;
wire n_6793;
wire n_15762;
wire n_2828;
wire n_13620;
wire n_5397;
wire n_4471;
wire n_10575;
wire n_11746;
wire n_20794;
wire n_3430;
wire n_7568;
wire n_15331;
wire n_3208;
wire n_5695;
wire n_2379;
wire n_14227;
wire n_14345;
wire n_11330;
wire n_15896;
wire n_7965;
wire n_6928;
wire n_13283;
wire n_15857;
wire n_20110;
wire n_13555;
wire n_20241;
wire n_4786;
wire n_7026;
wire n_326;
wire n_5854;
wire n_16376;
wire n_16731;
wire n_7002;
wire n_8898;
wire n_8410;
wire n_7141;
wire n_14019;
wire n_21819;
wire n_13809;
wire n_1199;
wire n_11102;
wire n_15622;
wire n_20832;
wire n_1841;
wire n_18732;
wire n_20685;
wire n_21261;
wire n_6027;
wire n_9254;
wire n_15345;
wire n_9529;
wire n_20722;
wire n_2581;
wire n_19003;
wire n_21358;
wire n_3752;
wire n_14627;
wire n_6638;
wire n_1891;
wire n_10651;
wire n_21737;
wire n_5254;
wire n_19464;
wire n_2546;
wire n_21769;
wire n_12731;
wire n_13644;
wire n_11686;
wire n_9726;
wire n_8823;
wire n_10851;
wire n_16486;
wire n_12383;
wire n_4613;
wire n_15041;
wire n_20150;
wire n_14709;
wire n_1963;
wire n_5902;
wire n_7768;
wire n_13294;
wire n_20745;
wire n_16669;
wire n_12902;
wire n_16723;
wire n_7357;
wire n_5083;
wire n_6927;
wire n_9627;
wire n_7975;
wire n_1194;
wire n_13380;
wire n_8172;
wire n_4186;
wire n_7310;
wire n_18645;
wire n_7521;
wire n_2190;
wire n_7593;
wire n_4742;
wire n_6256;
wire n_3620;
wire n_1260;
wire n_5870;
wire n_13884;
wire n_4295;
wire n_14415;
wire n_16778;
wire n_15594;
wire n_10451;
wire n_12718;
wire n_21102;
wire n_10201;
wire n_12249;
wire n_11814;
wire n_20048;
wire n_20714;
wire n_20324;
wire n_12932;
wire n_9465;
wire n_8456;
wire n_9970;
wire n_13719;
wire n_5081;
wire n_10278;
wire n_5124;
wire n_17161;
wire n_17500;
wire n_5807;
wire n_20141;
wire n_4244;
wire n_16203;
wire n_9129;
wire n_14616;
wire n_4697;
wire n_7137;
wire n_9957;
wire n_10915;
wire n_9558;
wire n_11292;
wire n_15642;
wire n_11487;
wire n_18828;
wire n_17119;
wire n_949;
wire n_8514;
wire n_14628;
wire n_14117;
wire n_5954;
wire n_3263;
wire n_1001;
wire n_10773;
wire n_10621;
wire n_5047;
wire n_11600;
wire n_15506;
wire n_16143;
wire n_7125;
wire n_2577;
wire n_5109;
wire n_757;
wire n_13912;
wire n_15307;
wire n_9095;
wire n_2937;
wire n_8337;
wire n_11781;
wire n_11550;
wire n_7983;
wire n_18479;
wire n_2805;
wire n_12786;
wire n_13467;
wire n_4918;
wire n_16069;
wire n_3856;
wire n_9246;
wire n_16304;
wire n_7624;
wire n_12117;
wire n_14716;
wire n_19218;
wire n_20361;
wire n_18250;
wire n_21176;
wire n_14683;
wire n_2406;
wire n_18044;
wire n_14373;
wire n_20611;
wire n_3773;
wire n_8950;
wire n_2398;
wire n_13982;
wire n_21983;
wire n_13577;
wire n_6351;
wire n_4822;
wire n_17521;
wire n_2155;
wire n_11502;
wire n_4299;
wire n_4801;
wire n_13300;
wire n_1665;
wire n_12456;
wire n_11424;
wire n_2886;
wire n_13405;
wire n_3378;
wire n_14735;
wire n_1431;
wire n_4279;
wire n_14584;
wire n_17321;
wire n_660;
wire n_21876;
wire n_20161;
wire n_7139;
wire n_14655;
wire n_8640;
wire n_4294;
wire n_16947;
wire n_9332;
wire n_4232;
wire n_17432;
wire n_2941;
wire n_459;
wire n_18798;
wire n_15132;
wire n_17328;
wire n_723;
wire n_18475;
wire n_2536;
wire n_16531;
wire n_18954;
wire n_16902;
wire n_12464;
wire n_5321;
wire n_3058;
wire n_20014;
wire n_7964;
wire n_13135;
wire n_13721;
wire n_18507;
wire n_21560;
wire n_6019;
wire n_6222;
wire n_3505;
wire n_8838;
wire n_20455;
wire n_17813;
wire n_6486;
wire n_8766;
wire n_4992;
wire n_13628;
wire n_3001;
wire n_20560;
wire n_13326;
wire n_4542;
wire n_2261;
wire n_19673;
wire n_10897;
wire n_15894;
wire n_19561;
wire n_15151;
wire n_10287;
wire n_1612;
wire n_9321;
wire n_21021;
wire n_5857;
wire n_20641;
wire n_16204;
wire n_8173;
wire n_17055;
wire n_15283;
wire n_6087;
wire n_9951;
wire n_19536;
wire n_4597;
wire n_4329;
wire n_17036;
wire n_15416;
wire n_20847;
wire n_5756;
wire n_12294;
wire n_11336;
wire n_8851;
wire n_15069;
wire n_3453;
wire n_11262;
wire n_9359;
wire n_10402;
wire n_15083;
wire n_19797;
wire n_15280;
wire n_18669;
wire n_22006;
wire n_1041;
wire n_1562;
wire n_383;
wire n_7194;
wire n_17825;
wire n_20490;
wire n_11661;
wire n_3984;
wire n_11889;
wire n_15066;
wire n_239;
wire n_5927;
wire n_19253;
wire n_17206;
wire n_2716;
wire n_18132;
wire n_11756;
wire n_13153;
wire n_20135;
wire n_11419;
wire n_3888;
wire n_9975;
wire n_13763;
wire n_18251;
wire n_12778;
wire n_17004;
wire n_14994;
wire n_9942;
wire n_11081;
wire n_2803;
wire n_13304;
wire n_13711;
wire n_1846;
wire n_21717;
wire n_8952;
wire n_11654;
wire n_1903;
wire n_19197;
wire n_10209;
wire n_18174;
wire n_17750;
wire n_21436;
wire n_19467;
wire n_12011;
wire n_19734;
wire n_11978;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_2645;
wire n_340;
wire n_2240;
wire n_11595;
wire n_16201;
wire n_574;
wire n_13305;
wire n_8299;
wire n_18204;
wire n_7245;
wire n_15303;
wire n_11235;
wire n_1327;
wire n_4763;
wire n_16776;
wire n_18120;
wire n_366;
wire n_13837;
wire n_11906;
wire n_21453;
wire n_18500;
wire n_10790;
wire n_5970;
wire n_13955;
wire n_12505;
wire n_8657;
wire n_4076;
wire n_21968;
wire n_4776;
wire n_2122;
wire n_18055;
wire n_2512;
wire n_9287;
wire n_20919;
wire n_18613;
wire n_16892;
wire n_17279;
wire n_14500;
wire n_18411;
wire n_21129;
wire n_2786;
wire n_13974;
wire n_15158;
wire n_6671;
wire n_10449;
wire n_645;
wire n_12164;
wire n_21777;
wire n_6591;
wire n_18782;
wire n_17944;
wire n_14929;
wire n_8609;
wire n_21752;
wire n_18644;
wire n_15640;
wire n_21627;
wire n_21012;
wire n_1893;
wire n_12140;
wire n_19780;
wire n_10920;
wire n_3546;
wire n_6893;
wire n_16626;
wire n_14261;
wire n_17368;
wire n_256;
wire n_11082;
wire n_10224;
wire n_2443;
wire n_3012;
wire n_21085;
wire n_17693;
wire n_419;
wire n_8476;
wire n_3244;
wire n_6028;
wire n_20470;
wire n_19598;
wire n_389;
wire n_3130;
wire n_5629;
wire n_4452;
wire n_13890;
wire n_5634;
wire n_376;
wire n_8137;
wire n_4355;
wire n_8469;
wire n_13270;
wire n_10808;
wire n_6798;
wire n_19629;
wire n_351;
wire n_5702;
wire n_5050;
wire n_5229;
wire n_2125;
wire n_11430;
wire n_1051;
wire n_20077;
wire n_13476;
wire n_4572;
wire n_3073;
wire n_12395;
wire n_13176;
wire n_1608;
wire n_20583;
wire n_18268;
wire n_9436;
wire n_18912;
wire n_9562;
wire n_11516;
wire n_11005;
wire n_5977;
wire n_6875;
wire n_19248;
wire n_2341;
wire n_16215;
wire n_16969;
wire n_15763;
wire n_17105;
wire n_6853;
wire n_15020;
wire n_17409;
wire n_5767;
wire n_6324;
wire n_18124;
wire n_5640;
wire n_8284;
wire n_12259;
wire n_20302;
wire n_991;
wire n_8810;
wire n_21127;
wire n_3255;
wire n_15778;
wire n_17437;
wire n_10443;
wire n_16923;
wire n_19436;
wire n_17532;
wire n_2997;
wire n_9946;
wire n_14383;
wire n_5168;
wire n_21699;
wire n_21233;
wire n_16492;
wire n_10274;
wire n_8373;
wire n_21036;
wire n_13525;
wire n_20093;
wire n_16197;
wire n_17694;
wire n_325;
wire n_17397;
wire n_16775;
wire n_5322;
wire n_14782;
wire n_20340;
wire n_1793;
wire n_14694;
wire n_7519;
wire n_17549;
wire n_12465;
wire n_1804;
wire n_20642;
wire n_17652;
wire n_4347;
wire n_10791;
wire n_2533;
wire n_14895;
wire n_11236;
wire n_14183;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_12852;
wire n_21239;
wire n_195;
wire n_20680;
wire n_1636;
wire n_13162;
wire n_3601;
wire n_6997;
wire n_11629;
wire n_10286;
wire n_12511;
wire n_1350;
wire n_1575;
wire n_20812;
wire n_10913;
wire n_18498;
wire n_9890;
wire n_14736;
wire n_10273;
wire n_16011;
wire n_12014;
wire n_2043;
wire n_8163;
wire n_13980;
wire n_17053;
wire n_10806;
wire n_1934;
wire n_5933;
wire n_15759;
wire n_20844;
wire n_12305;
wire n_17152;
wire n_4948;
wire n_21616;
wire n_1446;
wire n_472;
wire n_7023;
wire n_1807;
wire n_17555;
wire n_10694;
wire n_11509;
wire n_4010;
wire n_9832;
wire n_20328;
wire n_14480;
wire n_14663;
wire n_555;
wire n_4607;
wire n_9954;
wire n_14091;
wire n_2441;
wire n_1802;
wire n_17606;
wire n_3083;
wire n_21467;
wire n_21189;
wire n_15144;
wire n_21027;
wire n_9334;
wire n_20413;
wire n_2795;
wire n_8252;
wire n_15052;
wire n_14088;
wire n_13446;
wire n_17169;
wire n_8450;
wire n_21975;
wire n_9284;
wire n_16394;
wire n_14318;
wire n_19244;
wire n_9147;
wire n_8367;
wire n_3538;
wire n_21863;
wire n_8834;
wire n_6869;
wire n_16713;
wire n_11571;
wire n_4849;
wire n_17922;
wire n_5424;
wire n_3198;
wire n_13916;
wire n_19541;
wire n_20321;
wire n_14812;
wire n_588;
wire n_8471;
wire n_11904;
wire n_12324;
wire n_4247;
wire n_17189;
wire n_17262;
wire n_18179;
wire n_19841;
wire n_4018;
wire n_12643;
wire n_20401;
wire n_3900;
wire n_16397;
wire n_10185;
wire n_4902;
wire n_17820;
wire n_11656;
wire n_4409;
wire n_17285;
wire n_15412;
wire n_6569;
wire n_18216;
wire n_20494;
wire n_15356;
wire n_16916;
wire n_19468;
wire n_1908;
wire n_2259;
wire n_9614;
wire n_17551;
wire n_12948;
wire n_16589;
wire n_21742;
wire n_458;
wire n_2995;
wire n_13694;
wire n_3547;
wire n_9154;
wire n_1102;
wire n_20017;
wire n_16089;
wire n_19944;
wire n_6961;
wire n_4954;
wire n_12697;
wire n_2435;
wire n_9437;
wire n_5460;
wire n_9276;
wire n_6761;
wire n_9346;
wire n_20873;
wire n_11636;
wire n_6767;
wire n_19432;
wire n_19268;
wire n_18777;
wire n_4805;
wire n_18739;
wire n_14118;
wire n_10343;
wire n_17236;
wire n_5983;
wire n_5910;
wire n_13591;
wire n_19922;
wire n_16491;
wire n_18265;
wire n_9162;
wire n_861;
wire n_21648;
wire n_7752;
wire n_1904;
wire n_13631;
wire n_10807;
wire n_15166;
wire n_17573;
wire n_15265;
wire n_9401;
wire n_16171;
wire n_19879;
wire n_6921;
wire n_16502;
wire n_2219;
wire n_7845;
wire n_13122;
wire n_10750;
wire n_1726;
wire n_4631;
wire n_15628;
wire n_20308;
wire n_21598;
wire n_5464;
wire n_6565;
wire n_19237;
wire n_12679;
wire n_8261;
wire n_754;
wire n_3639;
wire n_7302;
wire n_8201;
wire n_19372;
wire n_7180;
wire n_1915;
wire n_1109;
wire n_20746;
wire n_12605;
wire n_16233;
wire n_1399;
wire n_21173;
wire n_2924;
wire n_10472;
wire n_20822;
wire n_14180;
wire n_808;
wire n_797;
wire n_1025;
wire n_4587;
wire n_20399;
wire n_21803;
wire n_13578;
wire n_18679;
wire n_13870;
wire n_14958;
wire n_7247;
wire n_17556;
wire n_13600;
wire n_536;
wire n_13843;
wire n_14707;
wire n_19098;
wire n_5204;
wire n_21582;
wire n_18533;
wire n_4094;
wire n_17574;
wire n_2866;
wire n_1418;
wire n_10184;
wire n_20621;
wire n_9057;
wire n_12497;
wire n_2425;
wire n_21074;
wire n_21051;
wire n_14544;
wire n_8861;
wire n_18026;
wire n_11749;
wire n_18312;
wire n_3934;
wire n_18388;
wire n_11490;
wire n_21519;
wire n_8191;
wire n_11704;
wire n_318;
wire n_2160;
wire n_21547;
wire n_2697;
wire n_3074;
wire n_14157;
wire n_20606;
wire n_8836;
wire n_6676;
wire n_3673;
wire n_6492;
wire n_18787;
wire n_12161;
wire n_3768;
wire n_605;
wire n_21262;
wire n_8446;
wire n_7742;
wire n_19900;
wire n_5795;
wire n_17743;
wire n_4022;
wire n_9989;
wire n_1531;
wire n_1334;
wire n_4869;
wire n_4035;
wire n_16277;
wire n_3294;
wire n_554;
wire n_11932;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_6648;
wire n_7880;
wire n_4601;
wire n_8857;
wire n_714;
wire n_909;
wire n_9667;
wire n_18988;
wire n_13159;
wire n_10815;
wire n_12928;
wire n_17221;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_2884;
wire n_21727;
wire n_7513;
wire n_12321;
wire n_11274;
wire n_11770;
wire n_3126;
wire n_4403;
wire n_17812;
wire n_3700;
wire n_5504;
wire n_19726;
wire n_20345;
wire n_147;
wire n_4223;
wire n_9885;
wire n_19379;
wire n_12698;
wire n_17980;
wire n_19475;
wire n_209;
wire n_21433;
wire n_5025;
wire n_8565;
wire n_6362;
wire n_14509;
wire n_20041;
wire n_21283;
wire n_16784;
wire n_8141;
wire n_6491;
wire n_10015;
wire n_17900;
wire n_18866;
wire n_9306;
wire n_2898;
wire n_7151;
wire n_11652;
wire n_6229;
wire n_10362;
wire n_16921;
wire n_1867;
wire n_481;
wire n_11331;
wire n_11640;
wire n_2573;
wire n_2939;
wire n_3807;
wire n_5884;
wire n_271;
wire n_2447;
wire n_5653;
wire n_10095;
wire n_19986;
wire n_5394;
wire n_17382;
wire n_6755;
wire n_2774;
wire n_20070;
wire n_1707;
wire n_7942;
wire n_853;
wire n_4655;
wire n_12477;
wire n_16777;
wire n_13156;
wire n_15531;
wire n_9644;
wire n_14051;
wire n_392;
wire n_3477;
wire n_5421;
wire n_8527;
wire n_704;
wire n_4399;
wire n_11681;
wire n_2781;
wire n_14724;
wire n_11522;
wire n_9750;
wire n_2778;
wire n_13164;
wire n_12145;
wire n_16888;
wire n_8988;
wire n_7368;
wire n_13624;
wire n_5889;
wire n_11578;
wire n_10916;
wire n_10208;
wire n_13714;
wire n_13655;
wire n_15142;
wire n_9616;
wire n_8004;
wire n_2167;
wire n_16609;
wire n_9291;
wire n_6442;
wire n_19025;
wire n_21309;
wire n_17737;
wire n_13606;
wire n_8908;
wire n_4259;
wire n_15067;
wire n_16003;
wire n_10384;
wire n_5543;
wire n_816;
wire n_10237;
wire n_18535;
wire n_14453;
wire n_4564;
wire n_17048;
wire n_3840;
wire n_7677;
wire n_8569;
wire n_19705;
wire n_18386;
wire n_328;
wire n_10118;
wire n_15260;
wire n_17819;
wire n_1842;
wire n_685;
wire n_6162;
wire n_4526;
wire n_1555;
wire n_11268;
wire n_20827;
wire n_6278;
wire n_11066;
wire n_21826;
wire n_4899;
wire n_6208;
wire n_20943;
wire n_14642;
wire n_2552;
wire n_20089;
wire n_9310;
wire n_19303;
wire n_14246;
wire n_7027;
wire n_8001;
wire n_5671;
wire n_8322;
wire n_8403;
wire n_2182;
wire n_13140;
wire n_3251;
wire n_19145;
wire n_2931;
wire n_13573;
wire n_17444;
wire n_8999;
wire n_5185;
wire n_8596;
wire n_10291;
wire n_3511;
wire n_18678;
wire n_20653;
wire n_7763;
wire n_21412;
wire n_7498;
wire n_3336;
wire n_3521;
wire n_8555;
wire n_15769;
wire n_21256;
wire n_13796;
wire n_16308;
wire n_13314;
wire n_8610;
wire n_13195;
wire n_21801;
wire n_14456;
wire n_12993;
wire n_19340;
wire n_10324;
wire n_20031;
wire n_12663;
wire n_7945;
wire n_6744;
wire n_3114;
wire n_12039;
wire n_20558;
wire n_8615;
wire n_18987;
wire n_9714;
wire n_19763;
wire n_4081;
wire n_3132;
wire n_4407;
wire n_648;
wire n_7291;
wire n_20466;
wire n_14840;
wire n_18876;
wire n_18375;
wire n_9753;
wire n_20796;
wire n_19387;
wire n_19076;
wire n_13017;
wire n_11137;
wire n_11607;
wire n_2036;
wire n_12930;
wire n_18725;
wire n_20094;
wire n_10649;
wire n_18390;
wire n_13529;
wire n_20163;
wire n_11265;
wire n_20566;
wire n_1642;
wire n_2279;
wire n_4446;
wire n_6475;
wire n_3884;
wire n_8470;
wire n_18029;
wire n_11739;
wire n_16919;
wire n_20158;
wire n_10060;
wire n_17690;
wire n_6496;
wire n_20167;
wire n_18883;
wire n_2892;
wire n_2907;
wire n_15230;
wire n_17051;
wire n_2049;
wire n_2273;
wire n_12885;
wire n_18871;
wire n_15204;
wire n_1160;
wire n_1258;
wire n_1074;
wire n_7980;
wire n_11617;
wire n_2113;
wire n_14952;
wire n_11581;
wire n_10981;
wire n_14626;
wire n_7695;
wire n_13850;
wire n_17564;
wire n_6357;
wire n_12616;
wire n_2256;
wire n_15845;
wire n_12287;
wire n_12217;
wire n_5106;
wire n_11867;
wire n_17903;
wire n_8642;
wire n_6985;
wire n_5319;
wire n_13552;
wire n_8624;
wire n_6238;
wire n_17474;
wire n_1622;
wire n_13495;
wire n_1180;
wire n_15030;
wire n_10441;
wire n_17762;
wire n_9149;
wire n_9174;
wire n_11175;
wire n_17243;
wire n_3705;
wire n_6548;
wire n_14755;
wire n_4705;
wire n_19269;
wire n_5455;
wire n_8894;
wire n_19625;
wire n_2268;
wire n_5706;
wire n_6366;
wire n_5337;
wire n_20484;
wire n_18066;
wire n_3912;
wire n_9835;
wire n_2771;
wire n_17625;
wire n_15663;
wire n_20569;
wire n_10934;
wire n_4477;
wire n_7560;
wire n_11291;
wire n_16618;
wire n_18658;
wire n_1501;
wire n_3086;
wire n_13139;
wire n_564;
wire n_6529;
wire n_17257;
wire n_8803;
wire n_9515;
wire n_8801;
wire n_17140;
wire n_14258;
wire n_21811;
wire n_7169;
wire n_15779;
wire n_7140;
wire n_11311;
wire n_2302;
wire n_15869;
wire n_9948;
wire n_7134;
wire n_292;
wire n_12234;
wire n_16657;
wire n_3434;
wire n_1806;
wire n_6892;
wire n_15653;
wire n_17267;
wire n_9423;
wire n_11378;
wire n_9660;
wire n_14472;
wire n_9108;
wire n_20613;
wire n_11222;
wire n_16917;
wire n_19823;
wire n_9631;
wire n_16130;
wire n_4330;
wire n_6683;
wire n_556;
wire n_2677;
wire n_13254;
wire n_16211;
wire n_18562;
wire n_20327;
wire n_15305;
wire n_19880;
wire n_19807;
wire n_902;
wire n_5352;
wire n_19228;
wire n_4991;
wire n_8138;
wire n_8990;
wire n_15616;
wire n_16529;
wire n_16698;
wire n_19665;
wire n_12988;
wire n_1098;
wire n_17973;
wire n_8190;
wire n_320;
wire n_15247;
wire n_1135;
wire n_8092;
wire n_3048;
wire n_6124;
wire n_2203;
wire n_1243;
wire n_12609;
wire n_14494;
wire n_14503;
wire n_9531;
wire n_7893;
wire n_4208;
wire n_17144;
wire n_7090;
wire n_20986;
wire n_21708;
wire n_21603;
wire n_17849;
wire n_14174;
wire n_5992;
wire n_16244;
wire n_4177;
wire n_6199;
wire n_11584;
wire n_5958;
wire n_7749;
wire n_19850;
wire n_12053;
wire n_19775;
wire n_10880;
wire n_17850;
wire n_10810;
wire n_7681;
wire n_308;
wire n_2149;
wire n_1078;
wire n_19935;
wire n_11920;
wire n_4276;
wire n_13388;
wire n_9944;
wire n_19401;
wire n_16245;
wire n_5170;
wire n_20814;
wire n_8304;
wire n_13915;
wire n_18869;
wire n_8586;
wire n_5107;
wire n_339;
wire n_16184;
wire n_347;
wire n_10835;
wire n_6100;
wire n_14815;
wire n_9521;
wire n_1414;
wire n_8212;
wire n_4975;
wire n_9759;
wire n_18843;
wire n_12781;
wire n_13204;
wire n_1852;
wire n_13085;
wire n_16497;
wire n_9378;
wire n_5602;
wire n_13778;
wire n_422;
wire n_15164;
wire n_8933;
wire n_14805;
wire n_2470;
wire n_16321;
wire n_17890;
wire n_7244;
wire n_5405;
wire n_9485;
wire n_4760;
wire n_4652;
wire n_18737;
wire n_12842;
wire n_1587;
wire n_19738;
wire n_8690;
wire n_1284;
wire n_16933;
wire n_3440;
wire n_15214;
wire n_17200;
wire n_6510;
wire n_1748;
wire n_9440;
wire n_12366;
wire n_2615;
wire n_446;
wire n_5842;
wire n_691;
wire n_14419;
wire n_5722;
wire n_19527;
wire n_11357;
wire n_7287;
wire n_363;
wire n_1582;
wire n_13383;
wire n_11386;
wire n_1836;
wire n_5492;
wire n_12122;
wire n_14600;
wire n_21977;
wire n_8835;
wire n_15038;
wire n_16145;
wire n_3936;
wire n_17401;
wire n_21572;
wire n_3821;
wire n_21181;
wire n_16859;
wire n_2700;
wire n_11221;
wire n_9807;
wire n_21571;
wire n_8963;
wire n_20532;
wire n_18730;
wire n_21990;
wire n_19792;
wire n_16958;
wire n_16474;
wire n_8353;
wire n_9390;
wire n_17577;
wire n_18889;
wire n_21799;
wire n_7773;
wire n_17735;
wire n_13333;
wire n_9518;
wire n_13826;
wire n_586;
wire n_12233;
wire n_20336;
wire n_18323;
wire n_11885;
wire n_4218;
wire n_10966;
wire n_5165;
wire n_18890;
wire n_19389;
wire n_954;
wire n_14761;
wire n_11380;
wire n_17805;
wire n_14420;
wire n_17858;
wire n_17104;
wire n_14059;
wire n_1623;
wire n_20011;
wire n_15854;
wire n_11539;
wire n_4161;
wire n_9373;
wire n_17896;
wire n_8606;
wire n_2462;
wire n_1532;
wire n_10351;
wire n_3625;
wire n_8868;
wire n_10408;
wire n_13340;
wire n_11731;
wire n_12760;
wire n_2331;
wire n_10656;
wire n_16622;
wire n_4844;
wire n_6296;
wire n_12318;
wire n_11531;
wire n_18476;
wire n_10639;
wire n_2979;
wire n_21139;
wire n_6288;
wire n_14517;
wire n_8718;
wire n_19649;
wire n_20503;
wire n_14512;
wire n_822;
wire n_5645;
wire n_11392;
wire n_13490;
wire n_13754;
wire n_21424;
wire n_11627;
wire n_4388;
wire n_12340;
wire n_12478;
wire n_8597;
wire n_4738;
wire n_6211;
wire n_13998;
wire n_20727;
wire n_16261;
wire n_8430;
wire n_19002;
wire n_8600;
wire n_6860;
wire n_16384;
wire n_20108;
wire n_2804;
wire n_8978;
wire n_414;
wire n_17611;
wire n_20579;
wire n_21854;
wire n_9848;
wire n_19198;
wire n_14911;
wire n_12689;
wire n_20932;
wire n_15021;
wire n_8278;
wire n_6645;
wire n_17045;
wire n_12271;
wire n_14006;
wire n_3150;
wire n_13780;
wire n_2413;
wire n_17289;
wire n_10090;
wire n_615;
wire n_15681;
wire n_10937;
wire n_13278;
wire n_16583;
wire n_705;
wire n_13836;
wire n_21117;
wire n_14181;
wire n_19686;
wire n_10568;
wire n_2518;
wire n_9464;
wire n_367;
wire n_4481;
wire n_3416;
wire n_2181;
wire n_10053;
wire n_13856;
wire n_17738;
wire n_10359;
wire n_14961;
wire n_15619;
wire n_7436;
wire n_15726;
wire n_20578;
wire n_7502;
wire n_1128;
wire n_7335;
wire n_7103;
wire n_10648;
wire n_10151;
wire n_6246;
wire n_14602;
wire n_19052;
wire n_590;
wire n_11194;
wire n_11804;
wire n_3770;
wire n_19963;
wire n_15976;
wire n_9717;
wire n_7020;
wire n_11244;
wire n_8175;
wire n_21383;
wire n_5336;
wire n_17927;
wire n_8850;
wire n_20508;
wire n_14865;
wire n_3220;
wire n_18611;
wire n_10589;
wire n_13501;
wire n_2054;
wire n_11991;
wire n_1559;
wire n_12150;
wire n_5693;
wire n_1744;
wire n_11183;
wire n_295;
wire n_3113;
wire n_2718;
wire n_17350;
wire n_20574;
wire n_19104;
wire n_16542;
wire n_19239;
wire n_18387;
wire n_19400;
wire n_4360;
wire n_7825;
wire n_9001;
wire n_17213;
wire n_3828;
wire n_10218;
wire n_13482;
wire n_17874;
wire n_18430;
wire n_12964;
wire n_5514;
wire n_8578;
wire n_1509;
wire n_2613;
wire n_6626;
wire n_6563;
wire n_10775;
wire n_17441;
wire n_3558;
wire n_11114;
wire n_17536;
wire n_16637;
wire n_14771;
wire n_15834;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_6473;
wire n_10637;
wire n_15043;
wire n_20320;
wire n_1492;
wire n_15728;
wire n_592;
wire n_9397;
wire n_11775;
wire n_2481;
wire n_10834;
wire n_18063;
wire n_6688;
wire n_19482;
wire n_18306;
wire n_21938;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_9179;
wire n_2339;
wire n_6714;
wire n_7462;
wire n_603;
wire n_16285;
wire n_16710;
wire n_10619;
wire n_19154;
wire n_3426;
wire n_13801;
wire n_11322;
wire n_19398;
wire n_18048;
wire n_18874;
wire n_7401;
wire n_20367;
wire n_9169;
wire n_16603;
wire n_5298;
wire n_16660;
wire n_13996;
wire n_4413;
wire n_16889;
wire n_18337;
wire n_16798;
wire n_662;
wire n_4493;
wire n_218;
wire n_3475;
wire n_8181;
wire n_21213;
wire n_1592;
wire n_20292;
wire n_11467;
wire n_7288;
wire n_7124;
wire n_12668;
wire n_16995;
wire n_21089;
wire n_14969;
wire n_20201;
wire n_9166;
wire n_10265;
wire n_486;
wire n_20675;
wire n_12435;
wire n_13367;
wire n_17307;
wire n_21331;
wire n_13123;
wire n_1159;
wire n_15459;
wire n_5928;
wire n_3845;
wire n_18670;
wire n_15693;
wire n_11455;
wire n_299;
wire n_13930;
wire n_7386;
wire n_2156;
wire n_5101;
wire n_5019;
wire n_5911;
wire n_12029;
wire n_12548;
wire n_18569;
wire n_9641;
wire n_7187;
wire n_7544;
wire n_11087;
wire n_21520;
wire n_4606;
wire n_21371;
wire n_13108;
wire n_13948;
wire n_18719;
wire n_21922;
wire n_3887;
wire n_17335;
wire n_7255;
wire n_16056;
wire n_4672;
wire n_15016;
wire n_4174;
wire n_2367;
wire n_309;
wire n_10249;
wire n_19700;
wire n_9645;
wire n_16786;
wire n_4766;
wire n_8045;
wire n_17019;
wire n_21567;
wire n_5633;
wire n_8697;
wire n_21413;
wire n_8077;
wire n_1927;
wire n_8026;
wire n_3645;
wire n_6064;
wire n_18792;
wire n_7196;
wire n_10390;
wire n_2272;
wire n_14861;
wire n_21440;
wire n_19455;
wire n_5501;
wire n_20225;
wire n_21868;
wire n_12112;
wire n_5377;
wire n_18452;
wire n_13168;
wire n_874;
wire n_13574;
wire n_12346;
wire n_20984;
wire n_11853;
wire n_7081;
wire n_9307;
wire n_19508;
wire n_10795;
wire n_2066;
wire n_7968;
wire n_7832;
wire n_9238;
wire n_13581;
wire n_12732;
wire n_13138;
wire n_18307;
wire n_20983;
wire n_7584;
wire n_21671;
wire n_3366;
wire n_12863;
wire n_12347;
wire n_15188;
wire n_1534;
wire n_11898;
wire n_4863;
wire n_1205;
wire n_12041;
wire n_19830;
wire n_11710;
wire n_6808;
wire n_16854;
wire n_20407;
wire n_15460;
wire n_10878;
wire n_2405;
wire n_2953;
wire n_14169;
wire n_14086;
wire n_16511;
wire n_15074;
wire n_15470;
wire n_6251;
wire n_14309;
wire n_12088;
wire n_16688;
wire n_14204;
wire n_3483;
wire n_17308;
wire n_13202;
wire n_2740;
wire n_15930;
wire n_8056;
wire n_20540;
wire n_17823;
wire n_1274;
wire n_7623;
wire n_8954;
wire n_13590;
wire n_20329;
wire n_426;
wire n_20748;
wire n_8840;
wire n_6467;
wire n_13456;
wire n_20207;
wire n_10477;
wire n_562;
wire n_13321;
wire n_18700;
wire n_14306;
wire n_20370;
wire n_11834;
wire n_20303;
wire n_21908;
wire n_16149;
wire n_12772;
wire n_2281;
wire n_10559;
wire n_17889;
wire n_11141;
wire n_12539;
wire n_13007;
wire n_8346;
wire n_9697;
wire n_4230;
wire n_16260;
wire n_18833;
wire n_7882;
wire n_8827;
wire n_13196;
wire n_9060;
wire n_12775;
wire n_3941;
wire n_20939;
wire n_21355;
wire n_16362;
wire n_19899;
wire n_17721;
wire n_16676;
wire n_18687;
wire n_10572;
wire n_1808;
wire n_316;
wire n_2650;
wire n_16091;
wire n_5003;
wire n_10139;
wire n_17263;
wire n_10230;
wire n_14294;
wire n_21380;
wire n_16594;
wire n_17120;
wire n_21188;
wire n_20121;
wire n_19210;
wire n_15597;
wire n_16755;
wire n_4122;
wire n_11144;
wire n_7365;
wire n_9653;
wire n_6277;
wire n_7395;
wire n_17302;
wire n_13373;
wire n_17807;
wire n_19697;
wire n_12957;
wire n_13014;
wire n_19621;
wire n_10255;
wire n_3162;
wire n_20404;
wire n_15881;
wire n_5720;
wire n_21293;
wire n_13022;
wire n_17460;
wire n_2304;
wire n_762;
wire n_5325;
wire n_15380;
wire n_2637;
wire n_17763;
wire n_17664;
wire n_20522;
wire n_4384;
wire n_17830;
wire n_17990;
wire n_4423;
wire n_10063;
wire n_18962;
wire n_19334;
wire n_6616;
wire n_1203;
wire n_13136;
wire n_14690;
wire n_15288;
wire n_14532;
wire n_7871;
wire n_4996;
wire n_4598;
wire n_14944;
wire n_9215;
wire n_2646;
wire n_20695;
wire n_13630;
wire n_16053;
wire n_9407;
wire n_13269;
wire n_21243;
wire n_14570;
wire n_21543;
wire n_20961;
wire n_16523;
wire n_11897;
wire n_10368;
wire n_3921;
wire n_828;
wire n_13031;
wire n_5738;
wire n_7649;
wire n_17524;
wire n_17429;
wire n_21295;
wire n_5215;
wire n_9153;
wire n_945;
wire n_19108;
wire n_21090;
wire n_10173;
wire n_11554;
wire n_10644;
wire n_10323;
wire n_694;
wire n_17731;
wire n_17204;
wire n_1983;
wire n_10229;
wire n_9737;
wire n_11688;
wire n_1594;
wire n_19397;
wire n_6379;
wire n_3529;
wire n_7358;
wire n_10622;
wire n_1147;
wire n_21673;
wire n_18049;
wire n_9026;
wire n_9710;
wire n_15665;
wire n_8710;
wire n_13512;
wire n_19634;
wire n_16837;
wire n_14557;
wire n_16526;
wire n_18600;
wire n_21638;
wire n_14436;
wire n_16954;
wire n_2901;
wire n_14524;
wire n_17148;
wire n_13375;
wire n_13852;
wire n_3998;
wire n_14378;
wire n_11158;
wire n_7270;
wire n_13473;
wire n_8893;
wire n_14923;
wire n_12317;
wire n_5121;
wire n_9479;
wire n_3386;
wire n_12724;
wire n_4667;
wire n_16310;
wire n_15155;
wire n_3488;
wire n_18440;
wire n_1035;
wire n_14891;
wire n_11161;
wire n_5784;
wire n_6272;
wire n_7699;
wire n_6236;
wire n_8620;
wire n_8298;
wire n_11614;
wire n_4953;
wire n_6958;
wire n_21693;
wire n_10270;
wire n_8235;
wire n_21266;
wire n_430;
wire n_9294;
wire n_13773;
wire n_11263;
wire n_13066;
wire n_20816;
wire n_15109;
wire n_17196;
wire n_13469;
wire n_10992;
wire n_2377;
wire n_17218;
wire n_11257;
wire n_16844;
wire n_18162;
wire n_16904;
wire n_12664;
wire n_15885;
wire n_2361;
wire n_13450;
wire n_12206;
wire n_1603;
wire n_15081;
wire n_21847;
wire n_969;
wire n_19646;
wire n_4113;
wire n_16517;
wire n_20053;
wire n_8097;
wire n_10327;
wire n_18860;
wire n_8902;
wire n_10365;
wire n_18714;
wire n_15435;
wire n_5506;
wire n_3966;
wire n_15061;
wire n_9819;
wire n_13725;
wire n_21786;
wire n_18166;
wire n_4872;
wire n_16005;
wire n_7283;
wire n_18758;
wire n_5038;
wire n_11323;
wire n_6448;
wire n_12982;
wire n_7304;
wire n_10143;
wire n_14872;
wire n_15705;
wire n_1187;
wire n_7756;
wire n_13150;
wire n_8580;
wire n_3324;
wire n_3914;
wire n_18235;
wire n_3742;
wire n_17581;
wire n_17088;
wire n_1685;
wire n_1714;
wire n_9341;
wire n_14164;
wire n_14165;
wire n_6242;
wire n_10681;
wire n_12942;
wire n_12750;
wire n_17435;
wire n_12729;
wire n_19465;
wire n_6206;
wire n_2373;
wire n_19743;
wire n_17033;
wire n_17296;
wire n_14239;
wire n_3817;
wire n_1253;
wire n_13805;
wire n_1059;
wire n_11169;
wire n_11041;
wire n_17707;
wire n_21813;
wire n_7230;
wire n_8700;
wire n_11160;
wire n_10957;
wire n_5011;
wire n_3318;
wire n_16028;
wire n_4282;
wire n_16799;
wire n_4180;
wire n_19421;
wire n_1440;
wire n_16763;
wire n_9482;
wire n_3333;
wire n_8637;
wire n_5651;
wire n_8757;
wire n_4143;
wire n_14794;
wire n_5819;
wire n_205;
wire n_18461;
wire n_9193;
wire n_1812;
wire n_12069;
wire n_17570;
wire n_9527;
wire n_20892;
wire n_3791;
wire n_3368;
wire n_14028;
wire n_13170;
wire n_14368;
wire n_18830;
wire n_19560;
wire n_14374;
wire n_2994;
wire n_3135;
wire n_1457;
wire n_8709;
wire n_10825;
wire n_20803;
wire n_17937;
wire n_6722;
wire n_3573;
wire n_9943;
wire n_17717;
wire n_18075;
wire n_6428;
wire n_20056;
wire n_3534;
wire n_12818;
wire n_17764;
wire n_11132;
wire n_12531;
wire n_594;
wire n_200;
wire n_20422;
wire n_8108;
wire n_21855;
wire n_17681;
wire n_985;
wire n_5850;
wire n_10014;
wire n_13454;
wire n_5111;
wire n_17070;
wire n_18971;
wire n_15968;
wire n_20067;
wire n_3973;
wire n_3670;
wire n_13758;
wire n_10830;
wire n_17025;
wire n_2023;
wire n_2351;
wire n_17127;
wire n_8490;
wire n_21042;
wire n_5113;
wire n_9491;
wire n_4698;
wire n_642;
wire n_17583;
wire n_1602;
wire n_1178;
wire n_18396;
wire n_19072;
wire n_16299;
wire n_19329;
wire n_4966;
wire n_503;
wire n_18282;
wire n_18690;
wire n_20364;
wire n_8808;
wire n_3397;
wire n_3740;
wire n_11811;
wire n_19689;
wire n_8685;
wire n_13877;
wire n_703;
wire n_19799;
wire n_780;
wire n_8701;
wire n_11212;
wire n_6303;
wire n_6182;
wire n_16114;
wire n_15118;
wire n_21537;
wire n_12984;
wire n_2836;
wire n_5682;
wire n_15170;
wire n_16194;
wire n_20826;
wire n_14330;
wire n_8875;
wire n_6392;
wire n_898;
wire n_3239;
wire n_5117;
wire n_3686;
wire n_11477;
wire n_7999;
wire n_14347;
wire n_21696;
wire n_1791;
wire n_18491;
wire n_12086;
wire n_8389;
wire n_3982;
wire n_15289;
wire n_17203;
wire n_14823;
wire n_20901;
wire n_20478;
wire n_18105;
wire n_4559;
wire n_12703;
wire n_12411;
wire n_4368;
wire n_7382;
wire n_13337;
wire n_8814;
wire n_13867;
wire n_5301;
wire n_9286;
wire n_4642;
wire n_11313;
wire n_5898;
wire n_3576;
wire n_11206;
wire n_7298;
wire n_1792;
wire n_6641;
wire n_3495;
wire n_17131;
wire n_10696;
wire n_7074;
wire n_20232;
wire n_21049;
wire n_11223;
wire n_16872;
wire n_4724;
wire n_5832;
wire n_18721;
wire n_16614;
wire n_1238;
wire n_11515;
wire n_16747;
wire n_9265;
wire n_19014;
wire n_19835;
wire n_21205;
wire n_282;
wire n_752;
wire n_9080;
wire n_1108;
wire n_12645;
wire n_6367;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_9770;
wire n_2889;
wire n_20386;
wire n_9463;
wire n_7001;
wire n_5593;
wire n_10580;
wire n_16759;
wire n_1675;
wire n_1924;
wire n_19704;
wire n_9939;
wire n_21456;
wire n_11390;
wire n_5211;
wire n_10122;
wire n_17106;
wire n_14320;
wire n_19041;
wire n_3056;
wire n_17915;
wire n_9691;
wire n_5110;
wire n_16223;
wire n_379;
wire n_3295;
wire n_4178;
wire n_18898;
wire n_13803;
wire n_7450;
wire n_14455;
wire n_10532;
wire n_15583;
wire n_5737;
wire n_16544;
wire n_786;
wire n_15178;
wire n_2579;
wire n_15889;
wire n_18008;
wire n_1716;
wire n_14113;
wire n_7439;
wire n_5560;
wire n_9155;
wire n_21883;
wire n_6399;
wire n_8623;
wire n_12109;
wire n_11438;
wire n_1087;
wire n_6575;
wire n_7924;
wire n_16338;
wire n_7732;
wire n_7040;
wire n_7325;
wire n_4968;
wire n_17155;
wire n_9201;
wire n_5961;
wire n_7459;
wire n_19532;
wire n_7191;
wire n_1247;
wire n_11051;
wire n_591;
wire n_12519;
wire n_13872;
wire n_3050;
wire n_17280;
wire n_19023;
wire n_9227;
wire n_21000;
wire n_5361;
wire n_369;
wire n_10939;
wire n_5847;
wire n_6678;
wire n_5068;
wire n_9025;
wire n_1460;
wire n_16543;
wire n_18039;
wire n_13086;
wire n_8282;
wire n_21372;
wire n_2702;
wire n_7697;
wire n_11685;
wire n_17982;
wire n_10955;
wire n_10824;
wire n_6748;
wire n_903;
wire n_20042;
wire n_4749;
wire n_17854;
wire n_1794;
wire n_9749;
wire n_9972;
wire n_10058;
wire n_20514;
wire n_7652;
wire n_14533;
wire n_21374;
wire n_6500;
wire n_9214;
wire n_2797;
wire n_13299;
wire n_11443;
wire n_9271;
wire n_12661;
wire n_18553;
wire n_5905;
wire n_1601;
wire n_10658;
wire n_16908;
wire n_2841;
wire n_19000;
wire n_7952;
wire n_10912;
wire n_4576;
wire n_19368;
wire n_2427;
wire n_16052;
wire n_18805;
wire n_3250;
wire n_2594;
wire n_5798;
wire n_14701;
wire n_12489;
wire n_4767;
wire n_7998;
wire n_17125;
wire n_10160;
wire n_1379;
wire n_4676;
wire n_17235;
wire n_11495;
wire n_14259;
wire n_12480;
wire n_13265;
wire n_13273;
wire n_4544;
wire n_17013;
wire n_2170;
wire n_8516;
wire n_1091;
wire n_641;
wire n_5676;
wire n_7307;
wire n_10631;
wire n_8237;
wire n_13372;
wire n_20971;
wire n_15897;
wire n_10852;
wire n_18024;
wire n_16469;
wire n_16800;
wire n_20609;
wire n_11406;
wire n_13121;
wire n_6370;
wire n_15634;
wire n_15836;
wire n_7039;
wire n_12624;
wire n_9107;
wire n_6859;
wire n_16461;
wire n_14574;
wire n_17146;
wire n_21344;
wire n_20807;
wire n_16014;
wire n_12771;
wire n_7443;
wire n_13262;
wire n_20307;
wire n_19974;
wire n_7811;
wire n_5341;
wire n_4320;
wire n_19274;
wire n_5930;
wire n_21614;
wire n_17418;
wire n_3613;
wire n_15806;
wire n_16538;
wire n_12544;
wire n_4012;
wire n_5518;
wire n_10125;
wire n_17102;
wire n_14810;
wire n_12931;
wire n_13940;
wire n_3910;
wire n_835;
wire n_17446;
wire n_7348;
wire n_18716;
wire n_4680;
wire n_2044;
wire n_13873;
wire n_3259;
wire n_5482;
wire n_2010;
wire n_8938;
wire n_21892;
wire n_8787;
wire n_21474;
wire n_10017;
wire n_6535;
wire n_14987;
wire n_18859;
wire n_1827;
wire n_16724;
wire n_16665;
wire n_8335;
wire n_13449;
wire n_14974;
wire n_5041;
wire n_13395;
wire n_14463;
wire n_1423;
wire n_5431;
wire n_19287;
wire n_2200;
wire n_16255;
wire n_14151;
wire n_5026;
wire n_15609;
wire n_10842;
wire n_2746;
wire n_18042;
wire n_8150;
wire n_5059;
wire n_12009;
wire n_5505;
wire n_3127;
wire n_9486;
wire n_226;
wire n_9134;
wire n_1055;
wire n_19500;
wire n_18209;
wire n_12481;
wire n_21184;
wire n_20252;
wire n_14307;
wire n_14407;
wire n_14715;
wire n_15595;
wire n_14563;
wire n_13558;
wire n_12562;
wire n_11494;
wire n_9182;
wire n_19757;
wire n_5908;
wire n_6018;
wire n_19524;
wire n_12744;
wire n_5212;
wire n_14107;
wire n_9591;
wire n_10033;
wire n_7177;
wire n_13027;
wire n_3766;
wire n_12615;
wire n_1353;
wire n_10886;
wire n_18454;
wire n_9261;
wire n_7379;
wire n_1666;
wire n_4165;
wire n_4866;
wire n_5931;
wire n_19506;
wire n_7435;
wire n_4109;
wire n_7813;
wire n_16278;
wire n_19070;
wire n_20006;
wire n_16996;
wire n_6654;
wire n_20173;
wire n_6740;
wire n_20184;
wire n_17787;
wire n_18796;
wire n_8379;
wire n_18128;
wire n_2538;
wire n_2105;
wire n_21980;
wire n_16484;
wire n_307;
wire n_5891;
wire n_1230;
wire n_18153;
wire n_17732;
wire n_10876;
wire n_20170;
wire n_11852;
wire n_6452;
wire n_3379;
wire n_4374;
wire n_14020;
wire n_6791;
wire n_21091;
wire n_18885;
wire n_8671;
wire n_7110;
wire n_19698;
wire n_19888;
wire n_1294;
wire n_21013;
wire n_10831;
wire n_18761;
wire n_7791;
wire n_8484;
wire n_18750;
wire n_2963;
wire n_11492;
wire n_7232;
wire n_11544;
wire n_21357;
wire n_18182;
wire n_8703;
wire n_21788;
wire n_20083;
wire n_16615;
wire n_10206;
wire n_21818;
wire n_4315;
wire n_12880;
wire n_6364;
wire n_6451;
wire n_14205;
wire n_15168;
wire n_2193;
wire n_5140;
wire n_7827;
wire n_11646;
wire n_19176;
wire n_18211;
wire n_8127;
wire n_21489;
wire n_3810;
wire n_15751;
wire n_17510;
wire n_18717;
wire n_12458;
wire n_10319;
wire n_21860;
wire n_5598;
wire n_11900;
wire n_9470;
wire n_18227;
wire n_17860;
wire n_12132;
wire n_14434;
wire n_5306;
wire n_19714;
wire n_12037;
wire n_9328;
wire n_19102;
wire n_16156;
wire n_9245;
wire n_10739;
wire n_8232;
wire n_18037;
wire n_2561;
wire n_7363;
wire n_18682;
wire n_3446;
wire n_9455;
wire n_4806;
wire n_9744;
wire n_8842;
wire n_5533;
wire n_11871;
wire n_18647;
wire n_17311;
wire n_6866;
wire n_18426;
wire n_19115;
wire n_20683;
wire n_12621;
wire n_11674;
wire n_1931;
wire n_10718;
wire n_4166;
wire n_7093;
wire n_17949;
wire n_1071;
wire n_15249;
wire n_20440;
wire n_14153;
wire n_1513;
wire n_15101;
wire n_4937;
wire n_13324;
wire n_10513;
wire n_18301;
wire n_21812;
wire n_4258;
wire n_4498;
wire n_16396;
wire n_14953;
wire n_1590;
wire n_10194;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_675;
wire n_17901;
wire n_15537;
wire n_8308;
wire n_4936;
wire n_13406;
wire n_5387;
wire n_9630;
wire n_13071;
wire n_8378;
wire n_4770;
wire n_881;
wire n_21162;
wire n_4907;
wire n_10021;
wire n_12381;
wire n_8500;
wire n_17809;
wire n_16820;
wire n_17384;
wire n_5018;
wire n_10457;
wire n_9934;
wire n_16762;
wire n_973;
wire n_13364;
wire n_8548;
wire n_3193;
wire n_1971;
wire n_14340;
wire n_20967;
wire n_15526;
wire n_12064;
wire n_12503;
wire n_10111;
wire n_1447;
wire n_11921;
wire n_13358;
wire n_5159;
wire n_15248;
wire n_18565;
wire n_3954;
wire n_14621;
wire n_16367;
wire n_20414;
wire n_20379;
wire n_7823;
wire n_7467;
wire n_19245;
wire n_14555;
wire n_21956;
wire n_19957;
wire n_2750;
wire n_7550;
wire n_21466;
wire n_9937;
wire n_15754;
wire n_18801;
wire n_10545;
wire n_7717;
wire n_5300;
wire n_10595;
wire n_13883;
wire n_18940;
wire n_4912;
wire n_9082;
wire n_11366;
wire n_14279;
wire n_9424;
wire n_9453;
wire n_13757;
wire n_16199;
wire n_1882;
wire n_9637;
wire n_6706;
wire n_14190;
wire n_4256;
wire n_21833;
wire n_14185;
wire n_6999;
wire n_7054;
wire n_19453;
wire n_6403;
wire n_9183;
wire n_13935;
wire n_13325;
wire n_6228;
wire n_11315;
wire n_19088;
wire n_20688;
wire n_14188;
wire n_21388;
wire n_4415;
wire n_6888;
wire n_4457;
wire n_17781;
wire n_9030;
wire n_20968;
wire n_18633;
wire n_20756;
wire n_1393;
wire n_9380;
wire n_5481;
wire n_8744;
wire n_2808;
wire n_6070;
wire n_2676;
wire n_1709;
wire n_11524;
wire n_5821;
wire n_4491;
wire n_6647;
wire n_5733;
wire n_8765;
wire n_15183;
wire n_17138;
wire n_5871;
wire n_16951;
wire n_4261;
wire n_15424;
wire n_11514;
wire n_12438;
wire n_18011;
wire n_4886;
wire n_21683;
wire n_7507;
wire n_1662;
wire n_15509;
wire n_5707;
wire n_13907;
wire n_9211;
wire n_5836;
wire n_18165;
wire n_914;
wire n_5281;
wire n_12887;
wire n_4473;
wire n_12898;
wire n_9677;
wire n_13464;
wire n_5048;
wire n_11954;
wire n_19144;
wire n_13611;
wire n_1479;
wire n_4480;
wire n_8195;
wire n_1892;
wire n_806;
wire n_1766;
wire n_7033;
wire n_9881;
wire n_324;
wire n_8462;
wire n_5561;
wire n_10391;
wire n_8377;
wire n_14390;
wire n_12509;
wire n_20271;
wire n_15666;
wire n_18865;
wire n_21770;
wire n_15208;
wire n_12365;
wire n_5875;
wire n_8103;
wire n_20330;
wire n_9682;
wire n_1790;
wire n_4720;
wire n_11540;
wire n_15397;
wire n_19420;
wire n_18822;
wire n_6101;
wire n_9415;
wire n_2563;
wire n_16426;
wire n_9845;
wire n_1830;
wire n_16506;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_6106;
wire n_9822;
wire n_17499;
wire n_7688;
wire n_2336;
wire n_17965;
wire n_11101;
wire n_254;
wire n_14313;
wire n_17777;
wire n_18931;
wire n_4175;
wire n_8288;
wire n_10613;
wire n_14719;
wire n_19207;
wire n_244;
wire n_1333;
wire n_11612;
wire n_5006;
wire n_14288;
wire n_7806;
wire n_10085;
wire n_14833;
wire n_12599;
wire n_1539;
wire n_5734;
wire n_21656;
wire n_21066;
wire n_8806;
wire n_16274;
wire n_10560;
wire n_21366;
wire n_16160;
wire n_20817;
wire n_1866;
wire n_8601;
wire n_21881;
wire n_14097;
wire n_4486;
wire n_9722;
wire n_2960;
wire n_9791;
wire n_633;
wire n_9229;
wire n_11603;
wire n_21119;
wire n_9603;
wire n_18378;
wire n_11060;
wire n_17345;
wire n_7448;
wire n_6244;
wire n_2290;
wire n_16212;
wire n_8768;
wire n_19945;
wire n_19035;
wire n_20117;
wire n_14388;
wire n_9309;
wire n_12418;
wire n_13853;
wire n_7852;
wire n_13762;
wire n_1049;
wire n_2145;
wire n_5725;
wire n_3030;
wire n_16054;
wire n_9454;
wire n_11744;
wire n_4961;
wire n_10352;
wire n_14962;
wire n_20069;
wire n_21829;
wire n_2035;
wire n_5190;
wire n_8433;
wire n_19313;
wire n_2509;
wire n_4317;
wire n_1362;
wire n_14413;
wire n_10911;
wire n_20996;
wire n_4154;
wire n_14050;
wire n_15587;
wire n_19821;
wire n_15179;
wire n_9256;
wire n_9706;
wire n_13044;
wire n_12448;
wire n_7900;
wire n_13723;
wire n_7136;
wire n_13923;
wire n_6055;
wire n_5138;
wire n_21576;
wire n_21155;
wire n_13472;
wire n_12129;
wire n_9133;
wire n_8115;
wire n_1434;
wire n_6165;
wire n_18751;
wire n_17475;
wire n_1045;
wire n_5349;
wire n_2038;
wire n_20240;
wire n_7810;
wire n_9109;
wire n_4640;
wire n_17468;
wire n_636;
wire n_18835;
wire n_16416;
wire n_21550;
wire n_6731;
wire n_5485;
wire n_19950;
wire n_10484;
wire n_21428;
wire n_5766;
wire n_16004;
wire n_13183;
wire n_9673;
wire n_13601;
wire n_8891;
wire n_1989;
wire n_17838;
wire n_2523;
wire n_255;
wire n_21415;
wire n_18141;
wire n_16881;
wire n_17466;
wire n_4453;
wire n_6881;
wire n_1578;
wire n_7665;
wire n_8131;
wire n_9230;
wire n_14947;
wire n_7764;
wire n_10198;
wire n_6216;
wire n_21762;
wire n_2585;
wire n_10638;
wire n_7170;
wire n_7314;
wire n_21570;
wire n_6509;
wire n_15882;
wire n_21008;
wire n_11657;
wire n_10483;
wire n_20073;
wire n_11717;
wire n_8844;
wire n_16312;
wire n_4660;
wire n_4392;
wire n_5611;
wire n_4661;
wire n_16438;
wire n_15002;
wire n_2111;
wire n_21319;
wire n_19290;
wire n_9786;
wire n_8584;
wire n_8932;
wire n_21768;
wire n_9467;
wire n_9372;
wire n_329;
wire n_7850;
wire n_15592;
wire n_1390;
wire n_6401;
wire n_6227;
wire n_8480;
wire n_12095;
wire n_10094;
wire n_18731;
wire n_19139;
wire n_21920;
wire n_12432;
wire n_17999;
wire n_16371;
wire n_21697;
wire n_14293;
wire n_8398;
wire n_19866;
wire n_4361;
wire n_14884;
wire n_4614;
wire n_9480;
wire n_12156;
wire n_9158;
wire n_18992;
wire n_14441;
wire n_15827;
wire n_13264;
wire n_15965;
wire n_11517;
wire n_11022;
wire n_10162;
wire n_12302;
wire n_8466;
wire n_12190;
wire n_10353;
wire n_8813;
wire n_1101;
wire n_5447;
wire n_18904;
wire n_6127;
wire n_2851;
wire n_7883;
wire n_1455;
wire n_6600;
wire n_767;
wire n_13869;
wire n_3692;
wire n_10724;
wire n_5747;
wire n_19058;
wire n_20180;
wire n_16740;
wire n_18448;
wire n_5969;
wire n_13350;
wire n_9114;
wire n_18748;
wire n_1961;
wire n_13615;
wire n_9469;
wire n_12746;
wire n_15452;
wire n_4139;
wire n_6746;
wire n_4031;
wire n_10780;
wire n_9501;
wire n_7720;
wire n_15417;
wire n_19054;
wire n_12973;
wire n_11385;
wire n_6506;
wire n_12916;
wire n_8650;
wire n_16202;
wire n_10870;
wire n_21019;
wire n_10267;
wire n_19163;
wire n_10379;
wire n_18586;
wire n_21805;
wire n_2368;
wire n_19140;
wire n_6687;
wire n_9075;
wire n_1082;
wire n_3961;
wire n_21783;
wire n_6780;
wire n_20868;
wire n_16928;
wire n_10497;
wire n_10354;
wire n_5603;
wire n_539;
wire n_10888;
wire n_21945;
wire n_19057;
wire n_18443;
wire n_9409;
wire n_14140;
wire n_3993;
wire n_10138;
wire n_4940;
wire n_5208;
wire n_1056;
wire n_15902;
wire n_13745;
wire n_10948;
wire n_14339;
wire n_14804;
wire n_4664;
wire n_15007;
wire n_3160;
wire n_18793;
wire n_21902;
wire n_18559;
wire n_10386;
wire n_6040;
wire n_1346;
wire n_4906;
wire n_20686;
wire n_17643;
wire n_20054;
wire n_15686;
wire n_17058;
wire n_11660;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_10448;
wire n_14985;
wire n_5115;
wire n_14110;
wire n_19223;
wire n_6393;
wire n_2333;
wire n_8566;
wire n_8086;
wire n_4297;
wire n_1632;
wire n_19940;
wire n_18173;
wire n_17399;
wire n_21706;
wire n_11841;
wire n_11658;
wire n_19399;
wire n_9703;
wire n_19680;
wire n_19660;
wire n_21740;
wire n_20854;
wire n_14920;
wire n_4536;
wire n_5967;
wire n_7569;
wire n_8942;
wire n_5345;
wire n_5357;
wire n_13179;
wire n_13429;
wire n_20018;
wire n_10320;
wire n_17946;
wire n_2472;
wire n_6812;
wire n_4755;
wire n_20022;
wire n_4960;
wire n_14216;
wire n_17971;
wire n_8652;
wire n_16032;
wire n_3864;
wire n_2732;
wire n_17758;
wire n_11545;
wire n_12974;
wire n_14078;
wire n_13717;
wire n_14314;
wire n_11465;
wire n_4362;
wire n_10304;
wire n_16243;
wire n_13804;
wire n_6123;
wire n_7500;
wire n_1301;
wire n_11394;
wire n_17081;
wire n_6082;
wire n_13660;
wire n_9232;
wire n_18825;
wire n_804;
wire n_16768;
wire n_11191;
wire n_2827;
wire n_9167;
wire n_5228;
wire n_10596;
wire n_11068;
wire n_20627;
wire n_19637;
wire n_5758;
wire n_4215;
wire n_17108;
wire n_10875;
wire n_15287;
wire n_4047;
wire n_5471;
wire n_5434;
wire n_19670;
wire n_21757;
wire n_16794;
wire n_22007;
wire n_20670;
wire n_18983;
wire n_19735;
wire n_13959;
wire n_2609;
wire n_11483;
wire n_5669;
wire n_11073;
wire n_18083;
wire n_14637;
wire n_12265;
wire n_1077;
wire n_19870;
wire n_15546;
wire n_17662;
wire n_14703;
wire n_6979;
wire n_17231;
wire n_6203;
wire n_17601;
wire n_3363;
wire n_18119;
wire n_12890;
wire n_1511;
wire n_14644;
wire n_6368;
wire n_20111;
wire n_6556;
wire n_2020;
wire n_19565;
wire n_10974;
wire n_5878;
wire n_5588;
wire n_11692;
wire n_3950;
wire n_11344;
wire n_4458;
wire n_12926;
wire n_4121;
wire n_5090;
wire n_7639;
wire n_12881;
wire n_4476;
wire n_10914;
wire n_13710;
wire n_11510;
wire n_14082;
wire n_19388;
wire n_7251;
wire n_21589;
wire n_19829;
wire n_20130;
wire n_20562;
wire n_21245;
wire n_6080;
wire n_13287;
wire n_20909;
wire n_21995;
wire n_8255;
wire n_14752;
wire n_21738;
wire n_17493;
wire n_4118;
wire n_14632;
wire n_17483;
wire n_5972;
wire n_681;
wire n_5916;
wire n_5984;
wire n_14636;
wire n_19610;
wire n_15036;
wire n_12001;
wire n_5132;
wire n_15879;
wire n_16103;
wire n_3085;
wire n_8130;
wire n_13627;
wire n_9412;
wire n_18779;
wire n_939;
wire n_482;
wire n_7438;
wire n_11270;
wire n_20265;
wire n_7574;
wire n_17911;
wire n_17357;
wire n_4524;
wire n_3971;
wire n_19869;
wire n_16381;
wire n_9418;
wire n_7868;
wire n_6973;
wire n_2949;
wire n_7285;
wire n_1653;
wire n_18164;
wire n_20927;
wire n_15802;
wire n_21323;
wire n_19180;
wire n_20855;
wire n_2794;
wire n_3145;
wire n_18357;
wire n_5369;
wire n_11935;
wire n_2657;
wire n_14423;
wire n_11822;
wire n_12805;
wire n_7008;
wire n_10404;
wire n_1441;
wire n_15318;
wire n_8432;
wire n_6111;
wire n_21441;
wire n_617;
wire n_18513;
wire n_1572;
wire n_16993;
wire n_12971;
wire n_15636;
wire n_9783;
wire n_14568;
wire n_2409;
wire n_11501;
wire n_10317;
wire n_3402;
wire n_9909;
wire n_21326;
wire n_10453;
wire n_18692;
wire n_12543;
wire n_16972;
wire n_2117;
wire n_13854;
wire n_1993;
wire n_5155;
wire n_14467;
wire n_1335;
wire n_11662;
wire n_14706;
wire n_15703;
wire n_3401;
wire n_6908;
wire n_7819;
wire n_20393;
wire n_14362;
wire n_19295;
wire n_9112;
wire n_6498;
wire n_6692;
wire n_11500;
wire n_17709;
wire n_3654;
wire n_10892;
wire n_17806;
wire n_18360;
wire n_10049;
wire n_9180;
wire n_16737;
wire n_4713;
wire n_14535;
wire n_6505;
wire n_18138;
wire n_20687;
wire n_14770;
wire n_9474;
wire n_7598;
wire n_14406;
wire n_17465;
wire n_19361;
wire n_895;
wire n_8192;
wire n_2121;
wire n_17366;
wire n_6877;
wire n_7426;
wire n_15355;
wire n_8350;
wire n_20731;
wire n_12526;
wire n_17412;
wire n_14410;
wire n_500;
wire n_1067;
wire n_3805;
wire n_19762;
wire n_10395;
wire n_3928;
wire n_9781;
wire n_12068;
wire n_538;
wire n_4654;
wire n_20870;
wire n_8254;
wire n_6374;
wire n_19991;
wire n_12784;
wire n_16259;
wire n_6017;
wire n_16624;
wire n_3974;
wire n_2283;
wire n_6937;
wire n_16695;
wire n_2197;
wire n_13554;
wire n_16253;
wire n_7442;
wire n_20734;
wire n_5700;
wire n_19415;
wire n_19969;
wire n_18516;
wire n_11784;
wire n_16934;
wire n_16144;
wire n_19012;
wire n_4704;
wire n_14269;
wire n_268;
wire n_2421;
wire n_17701;
wire n_6674;
wire n_17845;
wire n_15683;
wire n_21495;
wire n_2363;
wire n_13413;
wire n_21967;
wire n_7098;
wire n_11321;
wire n_15980;
wire n_16342;
wire n_7611;
wire n_20373;
wire n_9925;
wire n_10655;
wire n_3055;
wire n_12187;
wire n_3315;
wire n_15963;
wire n_3172;
wire n_6895;
wire n_4450;
wire n_8384;
wire n_13035;
wire n_5642;
wire n_14299;
wire n_7224;
wire n_14114;
wire n_11133;
wire n_7524;
wire n_15100;
wire n_8023;
wire n_13770;
wire n_11001;
wire n_7627;
wire n_9998;
wire n_932;
wire n_10654;
wire n_5118;
wire n_14112;
wire n_1409;
wire n_788;
wire n_20148;
wire n_2996;
wire n_559;
wire n_17367;
wire n_16055;
wire n_12640;
wire n_2315;
wire n_3228;
wire n_15302;
wire n_12699;
wire n_13696;
wire n_14834;
wire n_16915;
wire n_11780;
wire n_11421;
wire n_9856;
wire n_20402;
wire n_21789;
wire n_6118;
wire n_2950;
wire n_11793;
wire n_18465;
wire n_18359;
wire n_5220;
wire n_12814;
wire n_5732;
wire n_548;
wire n_5178;
wire n_15436;
wire n_16380;
wire n_19600;
wire n_518;
wire n_4008;
wire n_8014;
wire n_13783;
wire n_15493;
wire n_21033;
wire n_8564;
wire n_11969;
wire n_12685;
wire n_5077;
wire n_782;
wire n_18192;
wire n_1901;
wire n_6858;
wire n_11948;
wire n_18366;
wire n_8558;
wire n_3032;
wire n_10275;
wire n_7254;
wire n_20542;
wire n_7837;
wire n_20036;
wire n_3924;
wire n_769;
wire n_9831;
wire n_2006;
wire n_14395;
wire n_11064;
wire n_14187;
wire n_17682;
wire n_5314;
wire n_826;
wire n_2343;
wire n_12096;
wire n_21970;
wire n_12202;
wire n_6518;
wire n_4229;
wire n_4739;
wire n_13692;
wire n_16466;
wire n_12120;
wire n_3017;
wire n_5718;
wire n_11866;
wire n_19601;
wire n_21477;
wire n_8563;
wire n_15988;
wire n_4838;
wire n_2872;
wire n_14906;
wire n_12816;
wire n_522;
wire n_14486;
wire n_11552;
wire n_14807;
wire n_10010;
wire n_10226;
wire n_1577;
wire n_14964;
wire n_18279;
wire n_14640;
wire n_21018;
wire n_4181;
wire n_14412;
wire n_14391;
wire n_2764;
wire n_7046;
wire n_12720;
wire n_13365;
wire n_18566;
wire n_19499;
wire n_922;
wire n_3627;
wire n_8011;
wire n_19169;
wire n_14431;
wire n_12535;
wire n_13279;
wire n_15497;
wire n_3769;
wire n_16678;
wire n_6589;
wire n_16424;
wire n_12046;
wire n_10720;
wire n_7173;
wire n_21107;
wire n_6197;
wire n_7460;
wire n_18997;
wire n_3117;
wire n_9605;
wire n_14731;
wire n_10868;
wire n_11047;
wire n_14841;
wire n_9417;
wire n_8730;
wire n_13945;
wire n_3527;
wire n_9721;
wire n_14789;
wire n_10615;
wire n_20365;
wire n_14504;
wire n_15884;
wire n_11004;
wire n_11287;
wire n_5701;
wire n_4440;
wire n_11208;
wire n_7079;
wire n_11860;
wire n_462;
wire n_17595;
wire n_17970;
wire n_3300;
wire n_4303;
wire n_5797;
wire n_20107;
wire n_11181;
wire n_471;
wire n_5743;
wire n_1028;
wire n_4016;
wire n_20212;
wire n_1546;
wire n_8782;
wire n_5801;
wire n_14331;
wire n_17961;
wire n_7279;
wire n_18785;
wire n_3165;
wire n_19825;
wire n_15585;
wire n_12522;
wire n_170;
wire n_4461;
wire n_3234;
wire n_21052;
wire n_2381;
wire n_6661;
wire n_3303;
wire n_1654;
wire n_13411;
wire n_10731;
wire n_4101;
wire n_11074;
wire n_11063;
wire n_3591;
wire n_15034;
wire n_12025;
wire n_10926;
wire n_6963;
wire n_3930;
wire n_4448;
wire n_16712;
wire n_6832;
wire n_16823;
wire n_7836;
wire n_16224;
wire n_14473;
wire n_7564;
wire n_12158;
wire n_8673;
wire n_20667;
wire n_2503;
wire n_20766;
wire n_17295;
wire n_20883;
wire n_14083;
wire n_17906;
wire n_21080;
wire n_5502;
wire n_2027;
wire n_453;
wire n_9421;
wire n_2642;
wire n_8577;
wire n_15835;
wire n_19106;
wire n_1918;
wire n_16858;
wire n_4831;
wire n_2513;
wire n_18457;
wire n_3057;
wire n_10116;
wire n_12937;
wire n_8485;
wire n_21055;
wire n_13596;
wire n_20204;
wire n_2229;
wire n_13609;
wire n_6758;
wire n_13715;
wire n_13398;
wire n_251;
wire n_6874;
wire n_18451;
wire n_13235;
wire n_21914;
wire n_20897;
wire n_6030;
wire n_13091;
wire n_12976;
wire n_18222;
wire n_19241;
wire n_21026;
wire n_8005;
wire n_175;
wire n_4474;
wire n_20122;
wire n_9639;
wire n_9102;
wire n_10003;
wire n_2511;
wire n_8283;
wire n_13016;
wire n_13048;
wire n_19311;
wire n_3585;
wire n_438;
wire n_20467;
wire n_4214;
wire n_8176;
wire n_21169;
wire n_17129;
wire n_5158;
wire n_14942;
wire n_6708;
wire n_16696;
wire n_13939;
wire n_12221;
wire n_14389;
wire n_12851;
wire n_11431;
wire n_12691;
wire n_20935;
wire n_11177;
wire n_4129;
wire n_17842;
wire n_21764;
wire n_13985;
wire n_11454;
wire n_12989;
wire n_9221;
wire n_12739;
wire n_7389;
wire n_13074;
wire n_12791;
wire n_5472;
wire n_7602;
wire n_21187;
wire n_19480;
wire n_14483;
wire n_2955;
wire n_6002;
wire n_14696;
wire n_7554;
wire n_16471;
wire n_14903;
wire n_7693;
wire n_1198;
wire n_15661;
wire n_15391;
wire n_6557;
wire n_18013;
wire n_15515;
wire n_17550;
wire n_12692;
wire n_12403;
wire n_19528;
wire n_9578;
wire n_18122;
wire n_2185;
wire n_13451;
wire n_3270;
wire n_2143;
wire n_14124;
wire n_18249;
wire n_3595;
wire n_11572;
wire n_18238;
wire n_1347;
wire n_7532;
wire n_21623;
wire n_5143;
wire n_7724;
wire n_20105;
wire n_18002;
wire n_14838;
wire n_16833;
wire n_2374;
wire n_18948;
wire n_4734;
wire n_10004;
wire n_8928;
wire n_18422;
wire n_3501;
wire n_14540;
wire n_16509;
wire n_11806;
wire n_21601;
wire n_11504;
wire n_6778;
wire n_7946;
wire n_14622;
wire n_21460;
wire n_13769;
wire n_8957;
wire n_3851;
wire n_17774;
wire n_12600;
wire n_7933;
wire n_1896;
wire n_21367;
wire n_5283;
wire n_7669;
wire n_14720;
wire n_17126;
wire n_20144;
wire n_10133;
wire n_9471;
wire n_9048;
wire n_18052;
wire n_3880;
wire n_5122;
wire n_12005;
wire n_13426;
wire n_21898;
wire n_3186;
wire n_20473;
wire n_4501;
wire n_406;
wire n_15153;
wire n_12953;
wire n_15159;
wire n_21701;
wire n_546;
wire n_1280;
wire n_21916;
wire n_15432;
wire n_291;
wire n_5840;
wire n_19320;
wire n_3157;
wire n_17557;
wire n_20360;
wire n_6919;
wire n_7423;
wire n_17773;
wire n_17673;
wire n_20219;
wire n_18705;
wire n_5330;
wire n_15690;
wire n_4829;
wire n_8326;
wire n_13538;
wire n_10521;
wire n_15465;
wire n_12325;
wire n_20460;
wire n_1484;
wire n_21643;
wire n_5378;
wire n_20877;
wire n_17241;
wire n_6883;
wire n_21506;
wire n_13065;
wire n_5519;
wire n_1749;
wire n_18123;
wire n_16691;
wire n_196;
wire n_8155;
wire n_20457;
wire n_16592;
wire n_11633;
wire n_1394;
wire n_13221;
wire n_10232;
wire n_17182;
wire n_4944;
wire n_15581;
wire n_12054;
wire n_21767;
wire n_14552;
wire n_17222;
wire n_9828;
wire n_14355;
wire n_14448;
wire n_2908;
wire n_19394;
wire n_10089;
wire n_15538;
wire n_1862;
wire n_21744;
wire n_1239;
wire n_4942;
wire n_13671;
wire n_5844;
wire n_15610;
wire n_15075;
wire n_17815;
wire n_20504;
wire n_17187;
wire n_6250;
wire n_1167;
wire n_10632;
wire n_1384;
wire n_8050;
wire n_6736;
wire n_19943;
wire n_18837;
wire n_19463;
wire n_923;
wire n_10820;
wire n_6339;
wire n_14594;
wire n_7013;
wire n_12892;
wire n_1069;
wire n_3306;
wire n_5662;
wire n_17371;
wire n_4857;
wire n_3136;
wire n_12373;
wire n_4080;
wire n_2101;
wire n_14184;
wire n_17211;
wire n_12855;
wire n_3986;
wire n_10031;
wire n_15730;
wire n_14576;
wire n_15944;
wire n_12388;
wire n_6845;
wire n_14647;
wire n_9302;
wire n_21915;
wire n_12836;
wire n_21528;
wire n_5181;
wire n_18766;
wire n_1197;
wire n_11888;
wire n_3008;
wire n_15024;
wire n_3709;
wire n_11879;
wire n_11054;
wire n_20857;
wire n_1403;
wire n_15370;
wire n_5553;
wire n_4176;
wire n_15220;
wire n_8246;
wire n_21390;
wire n_7771;
wire n_13742;
wire n_9322;
wire n_11937;
wire n_5368;
wire n_18522;
wire n_10098;
wire n_18381;
wire n_10042;
wire n_8349;
wire n_14073;
wire n_19867;
wire n_6576;
wire n_7943;
wire n_13838;
wire n_7208;
wire n_21700;
wire n_12992;
wire n_349;
wire n_21032;
wire n_5499;
wire n_18287;
wire n_4788;
wire n_4986;
wire n_2152;
wire n_10444;
wire n_10054;
wire n_627;
wire n_21840;
wire n_16726;
wire n_19183;
wire n_7202;
wire n_9140;
wire n_5291;
wire n_10540;
wire n_14444;
wire n_16230;
wire n_11943;
wire n_19917;
wire n_10178;
wire n_11995;
wire n_12790;
wire n_12979;
wire n_16191;
wire n_12659;
wire n_3682;
wire n_9343;
wire n_18512;
wire n_4462;
wire n_7313;
wire n_5288;
wire n_21271;
wire n_561;
wire n_11568;
wire n_14384;
wire n_21038;
wire n_1712;
wire n_16350;
wire n_21488;
wire n_5218;
wire n_8785;
wire n_2625;
wire n_12606;
wire n_7337;
wire n_6989;
wire n_8512;
wire n_21870;
wire n_4630;
wire n_10971;
wire n_4643;
wire n_4331;
wire n_13051;
wire n_4846;
wire n_3296;
wire n_14064;
wire n_21301;
wire n_19289;
wire n_14745;
wire n_18503;
wire n_10282;
wire n_10900;
wire n_6146;
wire n_6270;
wire n_599;
wire n_4696;
wire n_1978;
wire n_19346;
wire n_8419;
wire n_16280;
wire n_639;
wire n_10858;
wire n_6353;
wire n_20762;
wire n_10769;
wire n_16739;
wire n_9446;
wire n_2763;
wire n_10023;
wire n_11877;
wire n_3643;
wire n_4876;
wire n_6345;
wire n_16336;
wire n_14324;
wire n_15939;
wire n_15361;
wire n_19256;
wire n_14567;
wire n_746;
wire n_16931;
wire n_7919;
wire n_3660;
wire n_14129;
wire n_1815;
wire n_15382;
wire n_8985;
wire n_18098;
wire n_5079;
wire n_913;
wire n_3833;
wire n_697;
wire n_19156;
wire n_1679;
wire n_4841;
wire n_19832;
wire n_6336;
wire n_20952;
wire n_19066;
wire n_17096;
wire n_4842;
wire n_7370;
wire n_3513;
wire n_11104;
wire n_11952;
wire n_6174;
wire n_1833;
wire n_13322;
wire n_6023;
wire n_2517;
wire n_284;
wire n_14894;
wire n_9947;
wire n_15758;
wire n_744;
wire n_15423;
wire n_629;
wire n_19449;
wire n_19190;
wire n_10962;
wire n_20166;
wire n_14624;
wire n_21265;
wire n_14868;
wire n_18488;
wire n_12332;
wire n_2469;
wire n_21862;
wire n_13317;
wire n_10642;
wire n_604;
wire n_17816;
wire n_3917;
wire n_6669;
wire n_9096;
wire n_20030;
wire n_10170;
wire n_10142;
wire n_18862;
wire n_21590;
wire n_498;
wire n_624;
wire n_5429;
wire n_11044;
wire n_6940;
wire n_4557;
wire n_4451;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3280;
wire n_14977;
wire n_5432;
wire n_16606;
wire n_3205;
wire n_13545;
wire n_3610;
wire n_8208;
wire n_15117;
wire n_1933;
wire n_1656;
wire n_9730;
wire n_13246;
wire n_16209;
wire n_20928;
wire n_21208;
wire n_204;
wire n_16444;
wire n_10374;
wire n_14367;
wire n_4324;
wire n_21665;
wire n_11892;
wire n_8647;
wire n_11013;
wire n_3271;
wire n_7332;
wire n_6660;
wire n_10529;
wire n_13823;
wire n_12396;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_12081;
wire n_13157;
wire n_724;
wire n_15982;
wire n_17449;
wire n_18329;
wire n_3173;
wire n_18349;
wire n_21199;
wire n_9596;
wire n_7409;
wire n_4692;
wire n_10667;
wire n_7258;
wire n_11916;
wire n_21146;
wire n_17064;
wire n_18747;
wire n_17607;
wire n_21658;
wire n_2171;
wire n_7765;
wire n_17666;
wire n_13310;
wire n_10340;
wire n_18225;
wire n_21438;
wire n_20577;
wire n_17761;
wire n_17477;
wire n_12701;
wire n_17886;
wire n_6400;
wire n_2299;
wire n_12342;
wire n_10256;
wire n_21580;
wire n_742;
wire n_5436;
wire n_3021;
wire n_17374;
wire n_20845;
wire n_20747;
wire n_16736;
wire n_10917;
wire n_13933;
wire n_6470;
wire n_14619;
wire n_3015;
wire n_10727;
wire n_20908;
wire n_1920;
wire n_1065;
wire n_10938;
wire n_18741;
wire n_9175;
wire n_4925;
wire n_15444;
wire n_13210;
wire n_1548;
wire n_8705;
wire n_9043;
wire n_11306;
wire n_3787;
wire n_15334;
wire n_9037;
wire n_12434;
wire n_20976;
wire n_17790;
wire n_12998;
wire n_13427;
wire n_12248;
wire n_11007;
wire n_21689;
wire n_19170;
wire n_12405;
wire n_700;
wire n_18521;
wire n_15320;
wire n_7727;
wire n_388;
wire n_1366;
wire n_11231;
wire n_3248;
wire n_1568;
wire n_2110;
wire n_20537;
wire n_8505;
wire n_19077;
wire n_10008;
wire n_15742;
wire n_512;
wire n_7684;
wire n_15629;
wire n_6178;
wire n_11575;
wire n_2132;
wire n_609;
wire n_15146;
wire n_7787;
wire n_19782;
wire n_20123;
wire n_4140;
wire n_8067;
wire n_12421;
wire n_14950;
wire n_13106;
wire n_17349;
wire n_891;
wire n_7849;
wire n_5186;
wire n_13126;
wire n_17520;
wire n_7367;
wire n_9851;
wire n_14818;
wire n_19914;
wire n_8679;
wire n_11982;
wire n_18574;
wire n_2464;
wire n_6715;
wire n_11395;
wire n_2831;
wire n_16668;
wire n_21984;
wire n_11887;
wire n_11301;
wire n_19563;
wire n_4545;
wire n_261;
wire n_19141;
wire n_8332;
wire n_11010;
wire n_15182;
wire n_8632;
wire n_7745;
wire n_19773;
wire n_10733;
wire n_14646;
wire n_9240;
wire n_11666;
wire n_18115;
wire n_11506;
wire n_21900;
wire n_8918;
wire n_19418;
wire n_7673;
wire n_21100;
wire n_18425;
wire n_16925;
wire n_17239;
wire n_16035;
wire n_1094;
wire n_9345;
wire n_12439;
wire n_15920;
wire n_8968;
wire n_8404;
wire n_12199;
wire n_11214;
wire n_14495;
wire n_2895;
wire n_11362;
wire n_17597;
wire n_11409;
wire n_15091;
wire n_3097;
wire n_12996;
wire n_16283;
wire n_12873;
wire n_3824;
wire n_16129;
wire n_6289;
wire n_5267;
wire n_21544;
wire n_4494;
wire n_20948;
wire n_1316;
wire n_17415;
wire n_3589;
wire n_20665;
wire n_18523;
wire n_11031;
wire n_2610;
wire n_14080;
wire n_20516;
wire n_6852;
wire n_11346;
wire n_21615;
wire n_5044;
wire n_5809;
wire n_17802;
wire n_162;
wire n_5365;
wire n_14888;
wire n_17116;
wire n_19006;
wire n_13729;
wire n_5045;
wire n_14739;
wire n_17609;
wire n_9635;
wire n_6818;
wire n_11190;
wire n_4754;
wire n_13992;
wire n_12736;
wire n_11818;
wire n_6753;
wire n_9581;
wire n_3053;
wire n_14625;
wire n_1141;
wire n_4585;
wire n_16970;
wire n_451;
wire n_18838;
wire n_1699;
wire n_17299;
wire n_2541;
wire n_8492;
wire n_6764;
wire n_14569;
wire n_1432;
wire n_4003;
wire n_16093;
wire n_11785;
wire n_841;
wire n_1954;
wire n_17040;
wire n_15960;
wire n_13061;
wire n_19956;
wire n_6627;
wire n_10027;
wire n_5761;
wire n_19893;
wire n_17940;
wire n_8854;
wire n_12333;
wire n_11912;
wire n_20758;
wire n_4046;
wire n_20709;
wire n_1974;
wire n_10426;
wire n_11284;
wire n_13500;
wire n_6636;
wire n_19404;
wire n_4199;
wire n_10617;
wire n_21971;
wire n_10909;
wire n_20586;
wire n_5478;
wire n_11298;
wire n_15733;
wire n_6243;
wire n_19644;
wire n_6022;
wire n_8686;
wire n_2236;
wire n_17312;
wire n_12904;
wire n_16900;
wire n_18684;
wire n_20831;
wire n_2460;
wire n_13520;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_8887;
wire n_3417;
wire n_1579;
wire n_14680;
wire n_21869;
wire n_20418;
wire n_11496;
wire n_19097;
wire n_6187;
wire n_20051;
wire n_15196;
wire n_13572;
wire n_17864;
wire n_19209;
wire n_12085;
wire n_18818;
wire n_3237;
wire n_9008;
wire n_8929;
wire n_6395;
wire n_17932;
wire n_3400;
wire n_6233;
wire n_4550;
wire n_8776;
wire n_18313;
wire n_3382;
wire n_7488;
wire n_21267;
wire n_10165;
wire n_1557;
wire n_13242;
wire n_13194;
wire n_14915;
wire n_16076;
wire n_13871;
wire n_9904;
wire n_9157;
wire n_21634;
wire n_18197;
wire n_5242;
wire n_15978;
wire n_21147;
wire n_17310;
wire n_19254;
wire n_7950;
wire n_13741;
wire n_2670;
wire n_19114;
wire n_11210;
wire n_20005;
wire n_1646;
wire n_15539;
wire n_8837;
wire n_7031;
wire n_20448;
wire n_2707;
wire n_8907;
wire n_19582;
wire n_14514;
wire n_19972;
wire n_14149;
wire n_21527;
wire n_16417;
wire n_14454;
wire n_13245;
wire n_6672;
wire n_2471;
wire n_1472;
wire n_17851;
wire n_21206;
wire n_10087;
wire n_18220;
wire n_17247;
wire n_5294;
wire n_20690;
wire n_16050;
wire n_10266;
wire n_10509;
wire n_20991;
wire n_21029;
wire n_5617;
wire n_4736;
wire n_1928;
wire n_5244;
wire n_16639;
wire n_8065;
wire n_6107;
wire n_9634;
wire n_17023;
wire n_20632;
wire n_11828;
wire n_12291;
wire n_13109;
wire n_10106;
wire n_336;
wire n_6232;
wire n_19354;
wire n_17955;
wire n_9903;
wire n_15712;
wire n_3608;
wire n_6932;
wire n_7036;
wire n_3177;
wire n_17425;
wire n_9748;
wire n_14072;
wire n_11876;
wire n_17392;
wire n_16165;
wire n_5787;
wire n_10954;
wire n_10388;
wire n_1088;
wire n_5249;
wire n_8849;
wire n_638;
wire n_7944;
wire n_5198;
wire n_11709;
wire n_10804;
wire n_7455;
wire n_5829;
wire n_4887;
wire n_4617;
wire n_11304;
wire n_18255;
wire n_12723;
wire n_7947;
wire n_12428;
wire n_10841;
wire n_21585;
wire n_1637;
wire n_5899;
wire n_13339;
wire n_13478;
wire n_17580;
wire n_4792;
wire n_11461;
wire n_18742;
wire n_1886;
wire n_19331;
wire n_4980;
wire n_12520;
wire n_11994;
wire n_13918;
wire n_17117;
wire n_9316;
wire n_13526;
wire n_17386;
wire n_20520;
wire n_5317;
wire n_1843;
wire n_11024;
wire n_3061;
wire n_8749;
wire n_7290;
wire n_15419;
wire n_13524;
wire n_8249;
wire n_8496;
wire n_19357;
wire n_7625;
wire n_5822;
wire n_18415;
wire n_12251;
wire n_4947;
wire n_11715;
wire n_19623;
wire n_16266;
wire n_5182;
wire n_4971;
wire n_2000;
wire n_206;
wire n_15310;
wire n_12542;
wire n_19135;
wire n_17834;
wire n_20914;
wire n_12585;
wire n_2307;
wire n_3408;
wire n_2722;
wire n_11613;
wire n_13942;
wire n_4875;
wire n_8695;
wire n_1771;
wire n_15789;
wire n_15864;
wire n_710;
wire n_3090;
wire n_17292;
wire n_18911;
wire n_3762;
wire n_15720;
wire n_20821;
wire n_15918;
wire n_16490;
wire n_1988;
wire n_14799;
wire n_8472;
wire n_9535;
wire n_6042;
wire n_18901;
wire n_1787;
wire n_4137;
wire n_19251;
wire n_10055;
wire n_7907;
wire n_11926;
wire n_8188;
wire n_13041;
wire n_14879;
wire n_6207;
wire n_20134;
wire n_12630;
wire n_6524;
wire n_10787;
wire n_17964;
wire n_6225;
wire n_4322;
wire n_8920;
wire n_7297;
wire n_16587;
wire n_12883;
wire n_9664;
wire n_2354;
wire n_12672;
wire n_17094;
wire n_21104;
wire n_17916;
wire n_10826;
wire n_13828;
wire n_4677;
wire n_17676;
wire n_5261;
wire n_6520;
wire n_14162;
wire n_21224;
wire n_18088;
wire n_9863;
wire n_9199;
wire n_3381;
wire n_5193;
wire n_20113;
wire n_12706;
wire n_4909;
wire n_10556;
wire n_15374;
wire n_17303;
wire n_810;
wire n_1144;
wire n_7487;
wire n_20236;
wire n_16293;
wire n_5993;
wire n_8833;
wire n_15169;
wire n_21141;
wire n_4634;
wire n_21720;
wire n_6432;
wire n_16104;
wire n_14354;
wire n_20079;
wire n_12583;
wire n_4380;
wire n_9893;
wire n_2601;
wire n_11928;
wire n_17339;
wire n_12551;
wire n_6760;
wire n_1907;
wire n_13817;
wire n_2686;
wire n_15700;
wire n_15929;
wire n_10338;
wire n_10205;
wire n_1985;
wire n_14275;
wire n_2906;
wire n_382;
wire n_14692;
wire n_8608;
wire n_1013;
wire n_13946;
wire n_17142;
wire n_12498;
wire n_10285;
wire n_14040;
wire n_5881;
wire n_8079;
wire n_12378;
wire n_6261;
wire n_4075;
wire n_3104;
wire n_19028;
wire n_17408;
wire n_5755;
wire n_825;
wire n_9274;
wire n_2819;
wire n_18947;
wire n_8702;
wire n_15999;
wire n_4136;
wire n_7858;
wire n_15172;
wire n_7385;
wire n_8662;
wire n_1922;
wire n_15694;
wire n_4794;
wire n_20951;
wire n_8436;
wire n_11154;
wire n_17803;
wire n_20655;
wire n_19672;
wire n_8033;
wire n_16599;
wire n_12417;
wire n_21145;
wire n_12209;
wire n_505;
wire n_3011;
wire n_7266;
wire n_4196;
wire n_17786;
wire n_6969;
wire n_18302;
wire n_8741;
wire n_13894;
wire n_1425;
wire n_5665;
wire n_21664;
wire n_15012;
wire n_4370;
wire n_14541;
wire n_1620;
wire n_15439;
wire n_18524;
wire n_6659;
wire n_6750;
wire n_15685;
wire n_14477;
wire n_1046;
wire n_13663;
wire n_22011;
wire n_15674;
wire n_18549;
wire n_7132;
wire n_8763;
wire n_13361;
wire n_12707;
wire n_21834;
wire n_1641;
wire n_1361;
wire n_9007;
wire n_13132;
wire n_20374;
wire n_6003;
wire n_13662;
wire n_10670;
wire n_9121;
wire n_4722;
wire n_6224;
wire n_10789;
wire n_1129;
wire n_18601;
wire n_10387;
wire n_10629;
wire n_13898;
wire n_276;
wire n_21649;
wire n_7293;
wire n_1225;
wire n_20889;
wire n_4092;
wire n_10860;
wire n_6891;
wire n_8860;
wire n_16927;
wire n_8003;
wire n_21798;
wire n_3344;
wire n_16746;
wire n_17283;
wire n_4465;
wire n_17471;
wire n_14849;
wire n_19895;
wire n_1223;
wire n_8524;
wire n_21688;
wire n_16200;
wire n_20040;
wire n_1567;
wire n_13650;
wire n_10524;
wire n_12737;
wire n_10376;
wire n_145;
wire n_1857;
wire n_18638;
wire n_479;
wire n_6267;
wire n_11523;
wire n_9525;
wire n_21533;
wire n_10697;
wire n_2357;
wire n_21776;
wire n_21806;
wire n_6437;
wire n_6610;
wire n_608;
wire n_10259;
wire n_19299;
wire n_20452;
wire n_15371;
wire n_3260;
wire n_4926;
wire n_1589;
wire n_14742;
wire n_15600;
wire n_19953;
wire n_14658;
wire n_5704;
wire n_7620;
wire n_18481;
wire n_2815;
wire n_5473;
wire n_18437;
wire n_4612;
wire n_10197;
wire n_19654;
wire n_19501;
wire n_8464;
wire n_13313;
wire n_16847;
wire n_9790;
wire n_16291;
wire n_5177;
wire n_3617;
wire n_11332;
wire n_7123;
wire n_10854;
wire n_17380;
wire n_7959;
wire n_7563;
wire n_19778;
wire n_20678;
wire n_20829;
wire n_1277;
wire n_14218;
wire n_22001;
wire n_9428;
wire n_3384;
wire n_9990;
wire n_16062;
wire n_16029;
wire n_4602;
wire n_18062;
wire n_9705;
wire n_19366;
wire n_7322;
wire n_17326;
wire n_18321;
wire n_12022;
wire n_12358;
wire n_12242;
wire n_4445;
wire n_17775;
wire n_18374;
wire n_20310;
wire n_18468;
wire n_10419;
wire n_21761;
wire n_4870;
wire n_2832;
wire n_362;
wire n_1975;
wire n_16427;
wire n_616;
wire n_18210;
wire n_4915;
wire n_6129;
wire n_20427;
wire n_3323;
wire n_16421;
wire n_16536;
wire n_16419;
wire n_14960;
wire n_7261;
wire n_2823;
wire n_1761;
wire n_10294;
wire n_10687;
wire n_18369;
wire n_9771;
wire n_10480;
wire n_354;
wire n_12627;
wire n_5270;
wire n_7834;
wire n_9905;
wire n_656;
wire n_9163;
wire n_1220;
wire n_18126;
wire n_2655;
wire n_4185;
wire n_16178;
wire n_20190;
wire n_20693;
wire n_16414;
wire n_18701;
wire n_19079;
wire n_20677;
wire n_17356;
wire n_5823;
wire n_13687;
wire n_9387;
wire n_21621;
wire n_12492;
wire n_19069;
wire n_14758;
wire n_3539;
wire n_10799;
wire n_17467;
wire n_10315;
wire n_285;
wire n_412;
wire n_4343;
wire n_17692;
wire n_4212;
wire n_4492;
wire n_7346;
wire n_20594;
wire n_5148;
wire n_15076;
wire n_17065;
wire n_7333;
wire n_1996;
wire n_3604;
wire n_3853;
wire n_10932;
wire n_17099;
wire n_20601;
wire n_10951;
wire n_4309;
wire n_10646;
wire n_262;
wire n_6511;
wire n_1254;
wire n_1026;
wire n_12568;
wire n_2109;
wire n_364;
wire n_9853;
wire n_7319;
wire n_20728;
wire n_12639;
wire n_6497;
wire n_9941;
wire n_9135;
wire n_14414;
wire n_3473;
wire n_10633;
wire n_15346;
wire n_2237;
wire n_15292;
wire n_5067;
wire n_10606;
wire n_16070;
wire n_3873;
wire n_11936;
wire n_3693;
wire n_17476;
wire n_17689;
wire n_7469;
wire n_3857;
wire n_13332;
wire n_21710;
wire n_2253;
wire n_10564;
wire n_17509;
wire n_19381;
wire n_5567;
wire n_12148;
wire n_15969;
wire n_6579;
wire n_15974;
wire n_16559;
wire n_14881;
wire n_18693;
wire n_14101;
wire n_1488;
wire n_15948;
wire n_5484;
wire n_10515;
wire n_2395;
wire n_20139;
wire n_5207;
wire n_12853;
wire n_2347;
wire n_6786;
wire n_12327;
wire n_4240;
wire n_2021;
wire n_7710;
wire n_19435;
wire n_2391;
wire n_16000;
wire n_3615;
wire n_2059;
wire n_7461;
wire n_12641;
wire n_9331;
wire n_6649;
wire n_7154;
wire n_19980;
wire n_12924;
wire n_19273;
wire n_21419;
wire n_6810;
wire n_14070;
wire n_11016;
wire n_3341;
wire n_17501;
wire n_20850;
wire n_2001;
wire n_14144;
wire n_1462;
wire n_16119;
wire n_18807;
wire n_17049;
wire n_17014;
wire n_19683;
wire n_16997;
wire n_3448;
wire n_11342;
wire n_15734;
wire n_16153;
wire n_21666;
wire n_2096;
wire n_9312;
wire n_10363;
wire n_7486;
wire n_13822;
wire n_9273;
wire n_21137;
wire n_18489;
wire n_19231;
wire n_21531;
wire n_11678;
wire n_6549;
wire n_8105;
wire n_18902;
wire n_668;
wire n_7867;
wire n_301;
wire n_19552;
wire n_3010;
wire n_18424;
wire n_10761;
wire n_11299;
wire n_13146;
wire n_21163;
wire n_13775;
wire n_15311;
wire n_11077;
wire n_16602;
wire n_12861;
wire n_17191;
wire n_7468;
wire n_14721;
wire n_14714;
wire n_17244;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_4927;
wire n_15543;
wire n_19085;
wire n_10745;
wire n_13178;
wire n_13072;
wire n_8114;
wire n_15657;
wire n_21092;
wire n_17870;
wire n_9993;
wire n_9208;
wire n_21867;
wire n_14729;
wire n_2091;
wire n_16388;
wire n_17914;
wire n_16722;
wire n_17101;
wire n_8158;
wire n_15727;
wire n_19641;
wire n_2032;
wire n_156;
wire n_17912;
wire n_10420;
wire n_12575;
wire n_17436;
wire n_11635;
wire n_19440;
wire n_20347;
wire n_18117;
wire n_5406;
wire n_12501;
wire n_14408;
wire n_15805;
wire n_3947;
wire n_11505;
wire n_10535;
wire n_6214;
wire n_3437;
wire n_7804;
wire n_19987;
wire n_12078;
wire n_3353;
wire n_12175;
wire n_16383;
wire n_11615;
wire n_10307;
wire n_8262;
wire n_8290;
wire n_696;
wire n_21448;
wire n_12626;
wire n_436;
wire n_5661;
wire n_20305;
wire n_6991;
wire n_5562;
wire n_16390;
wire n_19992;
wire n_2159;
wire n_13875;
wire n_6707;
wire n_5852;
wire n_3420;
wire n_18605;
wire n_13110;
wire n_6868;
wire n_17502;
wire n_16339;
wire n_19590;
wire n_10672;
wire n_521;
wire n_21040;
wire n_15551;
wire n_9027;
wire n_12225;
wire n_8962;
wire n_7402;
wire n_4484;
wire n_11316;
wire n_19787;
wire n_9966;
wire n_19136;
wire n_5689;
wire n_13087;
wire n_10392;
wire n_144;
wire n_12670;
wire n_15336;
wire n_12152;
wire n_7992;
wire n_9161;
wire n_19027;
wire n_3418;
wire n_8556;
wire n_4901;
wire n_21698;
wire n_6725;
wire n_197;
wire n_20649;
wire n_21252;
wire n_10514;
wire n_10958;
wire n_10562;
wire n_11273;
wire n_18060;
wire n_15008;
wire n_14792;
wire n_8653;
wire n_7712;
wire n_11303;
wire n_14711;
wire n_21068;
wire n_12751;
wire n_9824;
wire n_6686;
wire n_11664;
wire n_10523;
wire n_4836;
wire n_11720;
wire n_4020;
wire n_3915;
wire n_4414;
wire n_6584;
wire n_17587;
wire n_283;
wire n_7323;
wire n_18581;
wire n_14405;
wire n_17269;
wire n_13243;
wire n_10988;
wire n_18551;
wire n_21523;
wire n_1000;
wire n_16030;
wire n_19626;
wire n_16782;
wire n_2668;
wire n_13457;
wire n_5236;
wire n_6062;
wire n_6191;
wire n_7903;
wire n_1667;
wire n_16684;
wire n_16956;
wire n_4405;
wire n_5433;
wire n_8525;
wire n_1331;
wire n_4195;
wire n_13734;
wire n_21061;
wire n_1241;
wire n_9368;
wire n_5909;
wire n_17637;
wire n_440;
wire n_18389;
wire n_13458;
wire n_15760;
wire n_19306;
wire n_2385;
wire n_11520;
wire n_1527;
wire n_13416;
wire n_8931;
wire n_9072;
wire n_9612;
wire n_2324;
wire n_9971;
wire n_7127;
wire n_182;
wire n_407;
wire n_21370;
wire n_9720;
wire n_207;
wire n_10400;
wire n_17318;
wire n_17799;
wire n_21613;
wire n_15911;
wire n_2514;
wire n_6304;
wire n_8210;
wire n_5189;
wire n_17957;
wire n_16638;
wire n_21150;
wire n_4160;
wire n_13582;
wire n_15316;
wire n_11599;
wire n_3009;
wire n_17593;
wire n_14852;
wire n_5936;
wire n_16578;
wire n_12284;
wire n_21465;
wire n_9649;
wire n_8501;
wire n_15205;
wire n_154;
wire n_11535;
wire n_1711;
wire n_16732;
wire n_3526;
wire n_8953;
wire n_18794;
wire n_21230;
wire n_14046;
wire n_21827;
wire n_7718;
wire n_17383;
wire n_16629;
wire n_1888;
wire n_13360;
wire n_6269;
wire n_17316;
wire n_4795;
wire n_21044;
wire n_15165;
wire n_21512;
wire n_1690;
wire n_15632;
wire n_21596;
wire n_9106;
wire n_21624;
wire n_2449;
wire n_8247;
wire n_15257;
wire n_21258;
wire n_8941;
wire n_8940;
wire n_13021;
wire n_12070;
wire n_19481;
wire n_2177;
wire n_17464;
wire n_3747;
wire n_5698;
wire n_7716;
wire n_2876;
wire n_7406;
wire n_7600;
wire n_11353;
wire n_10223;
wire n_2479;
wire n_11823;
wire n_1444;
wire n_13686;
wire n_18328;
wire n_18558;
wire n_12719;
wire n_10215;
wire n_4694;
wire n_18573;
wire n_4533;
wire n_11138;
wire n_19265;
wire n_9894;
wire n_10100;
wire n_2871;
wire n_15425;
wire n_5863;
wire n_17810;
wire n_20348;
wire n_2943;
wire n_16553;
wire n_4254;
wire n_15341;
wire n_3143;
wire n_14842;
wire n_3168;
wire n_6982;
wire n_7286;
wire n_12625;
wire n_4190;
wire n_3994;
wire n_18596;
wire n_11753;
wire n_4810;
wire n_10689;
wire n_12371;
wire n_7539;
wire n_1121;
wire n_16231;
wire n_8769;
wire n_433;
wire n_7229;
wire n_16232;
wire n_13487;
wire n_8334;
wire n_1503;
wire n_22010;
wire n_8639;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_14342;
wire n_14916;
wire n_19225;
wire n_4527;
wire n_15186;
wire n_11844;
wire n_2796;
wire n_10874;
wire n_7869;
wire n_6466;
wire n_18034;
wire n_12602;
wire n_16501;
wire n_20290;
wire n_18428;
wire n_1851;
wire n_19043;
wire n_16363;
wire n_6008;
wire n_15048;
wire n_15338;
wire n_20002;
wire n_3095;
wire n_8257;
wire n_8125;
wire n_1145;
wire n_14860;
wire n_16718;
wire n_17455;
wire n_1153;
wire n_9683;
wire n_12110;
wire n_2914;
wire n_18506;
wire n_1964;
wire n_6805;
wire n_14334;
wire n_3623;
wire n_19707;
wire n_17481;
wire n_15776;
wire n_9899;
wire n_5358;
wire n_20954;
wire n_4619;
wire n_13034;
wire n_6004;
wire n_6901;
wire n_11965;
wire n_19333;
wire n_11997;
wire n_9094;
wire n_5580;
wire n_5937;
wire n_18006;
wire n_3515;
wire n_8339;
wire n_15898;
wire n_267;
wire n_1208;
wire n_3287;
wire n_13641;
wire n_5435;
wire n_10867;
wire n_11361;
wire n_19779;
wire n_4769;
wire n_19990;
wire n_10741;
wire n_5373;
wire n_5745;
wire n_15223;
wire n_19847;
wire n_5279;
wire n_8351;
wire n_18708;
wire n_11499;
wire n_19808;
wire n_8196;
wire n_11580;
wire n_16753;
wire n_15084;
wire n_17604;
wire n_18400;
wire n_7857;
wire n_9054;
wire n_10150;
wire n_18916;
wire n_13028;
wire n_14896;
wire n_13613;
wire n_12389;
wire n_2952;
wire n_4847;
wire n_7338;
wire n_20230;
wire n_5096;
wire n_16024;
wire n_4365;
wire n_9661;
wire n_10861;
wire n_1878;
wire n_15672;
wire n_11070;
wire n_11245;
wire n_19733;
wire n_10635;
wire n_12874;
wire n_14749;
wire n_14871;
wire n_12990;
wire n_7235;
wire n_5210;
wire n_8488;
wire n_16095;
wire n_11286;
wire n_21774;
wire n_6083;
wire n_6844;
wire n_8969;
wire n_12240;
wire n_11631;
wire n_303;
wire n_10555;
wire n_2729;
wire n_15793;
wire n_10983;
wire n_15243;
wire n_4500;
wire n_9800;
wire n_7437;
wire n_20461;
wire n_11053;
wire n_8420;
wire n_21255;
wire n_3185;
wire n_1300;
wire n_17675;
wire n_3523;
wire n_1006;
wire n_1664;
wire n_20228;
wire n_11247;
wire n_15943;
wire n_15523;
wire n_7449;
wire n_19324;
wire n_7329;
wire n_2390;
wire n_5708;
wire n_8687;
wire n_10001;
wire n_19744;
wire n_3077;
wire n_21890;
wire n_11363;
wire n_3474;
wire n_8740;
wire n_14450;
wire n_15664;
wire n_6807;
wire n_630;
wire n_21998;
wire n_2151;
wire n_7708;
wire n_5638;
wire n_10997;
wire n_16494;
wire n_9335;
wire n_4189;
wire n_8815;
wire n_17034;
wire n_1304;
wire n_3707;
wire n_12813;
wire n_11407;
wire n_19727;
wire n_9247;
wire n_9933;
wire n_21072;
wire n_12907;
wire n_19201;
wire n_21401;
wire n_429;
wire n_8128;
wire n_11519;
wire n_4687;
wire n_18148;
wire n_17327;
wire n_17071;
wire n_5664;
wire n_11668;
wire n_18933;
wire n_10829;
wire n_7281;
wire n_10233;
wire n_11810;
wire n_9362;
wire n_15723;
wire n_10311;
wire n_3421;
wire n_2436;
wire n_11198;
wire n_14712;
wire n_20751;
wire n_19955;
wire n_9216;
wire n_11168;
wire n_5262;
wire n_11872;
wire n_21056;
wire n_3286;
wire n_5963;
wire n_12007;
wire n_10146;
wire n_1684;
wire n_5310;
wire n_9152;
wire n_17974;
wire n_15139;
wire n_16827;
wire n_4594;
wire n_6153;
wire n_16769;
wire n_20886;
wire n_21501;
wire n_14528;
wire n_19427;
wire n_13908;
wire n_15019;
wire n_16241;
wire n_19981;
wire n_19709;
wire n_13461;
wire n_18772;
wire n_21646;
wire n_12577;
wire n_17069;
wire n_16175;
wire n_3215;
wire n_11122;
wire n_4102;
wire n_9511;
wire n_21522;
wire n_19457;
wire n_8081;
wire n_20691;
wire n_3171;
wire n_10407;
wire n_1437;
wire n_6266;
wire n_10950;
wire n_14235;
wire n_14425;
wire n_7161;
wire n_14352;
wire n_7153;
wire n_5213;
wire n_3677;
wire n_14609;
wire n_18433;
wire n_3468;
wire n_17248;
wire n_14196;
wire n_5690;
wire n_1123;
wire n_13312;
wire n_9248;
wire n_17237;
wire n_1382;
wire n_10321;
wire n_7535;
wire n_424;
wire n_1311;
wire n_10506;
wire n_19403;
wire n_7178;
wire n_7480;
wire n_15212;
wire n_19855;
wire n_6501;
wire n_10157;
wire n_12200;
wire n_20843;
wire n_14603;
wire n_3822;
wire n_912;
wire n_136;
wire n_16001;
wire n_14332;
wire n_5430;
wire n_18584;
wire n_6709;
wire n_15630;
wire n_14285;
wire n_17275;
wire n_14443;
wire n_515;
wire n_885;
wire n_5063;
wire n_18878;
wire n_5199;
wire n_12023;
wire n_14673;
wire n_8423;
wire n_5527;
wire n_6986;
wire n_12239;
wire n_21470;
wire n_11279;
wire n_10975;
wire n_280;
wire n_3178;
wire n_5355;
wire n_18557;
wire n_17913;
wire n_21209;
wire n_13961;
wire n_15342;
wire n_2289;
wire n_302;
wire n_14811;
wire n_1343;
wire n_2263;
wire n_10566;
wire n_15745;
wire n_19308;
wire n_11451;
wire n_17891;
wire n_2733;
wire n_20216;
wire n_11980;
wire n_7905;
wire n_2785;
wire n_4519;
wire n_18836;
wire n_6699;
wire n_18332;
wire n_2499;
wire n_10688;
wire n_12261;
wire n_16189;
wire n_18003;
wire n_15625;
wire n_5655;
wire n_11239;
wire n_12338;
wire n_9203;
wire n_18091;
wire n_12222;
wire n_4400;
wire n_943;
wire n_3326;
wire n_20377;
wire n_650;
wire n_11740;
wire n_286;
wire n_19009;
wire n_10482;
wire n_18552;
wire n_11012;
wire n_470;
wire n_17103;
wire n_14774;
wire n_19493;
wire n_20782;
wire n_16018;
wire n_6827;
wire n_942;
wire n_13042;
wire n_18436;
wire n_189;
wire n_14592;
wire n_21280;
wire n_3196;
wire n_8846;
wire n_17293;
wire n_4593;
wire n_6312;
wire n_3492;
wire n_17068;
wire n_4043;
wire n_19910;
wire n_5418;
wire n_15910;
wire n_17751;
wire n_2973;
wire n_16868;
wire n_1096;
wire n_2094;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_9883;
wire n_19127;
wire n_9361;
wire n_6131;
wire n_4893;
wire n_19877;
wire n_13059;
wire n_4000;
wire n_13681;
wire n_2025;
wire n_1458;
wire n_8972;
wire n_2559;
wire n_11351;
wire n_4748;
wire n_1219;
wire n_16673;
wire n_11271;
wire n_14421;
wire n_20550;
wire n_1814;
wire n_5123;
wire n_8737;
wire n_3636;
wire n_7961;
wire n_10953;
wire n_1722;
wire n_11761;
wire n_7847;
wire n_9997;
wire n_21841;
wire n_7149;
wire n_10847;
wire n_11565;
wire n_2981;
wire n_2282;
wire n_21185;
wire n_15786;
wire n_7700;
wire n_16964;
wire n_311;
wire n_18543;
wire n_2098;
wire n_1296;
wire n_16720;
wire n_3460;
wire n_16432;
wire n_10922;
wire n_16647;
wire n_20661;
wire n_10738;
wire n_13197;
wire n_17052;
wire n_7914;
wire n_445;
wire n_1895;
wire n_7967;
wire n_21921;
wire n_21226;
wire n_13925;
wire n_19602;
wire n_12130;
wire n_8474;
wire n_18927;
wire n_16789;
wire n_11131;
wire n_4518;
wire n_10591;
wire n_16565;
wire n_11673;
wire n_14348;
wire n_11701;
wire n_18276;
wire n_2270;
wire n_20016;
wire n_18802;
wire n_9494;
wire n_9551;
wire n_6639;
wire n_5496;
wire n_13189;
wire n_4052;
wire n_1499;
wire n_21540;
wire n_21435;
wire n_13392;
wire n_2633;
wire n_12574;
wire n_16871;
wire n_18150;
wire n_1164;
wire n_2097;
wire n_20783;
wire n_7628;
wire n_4304;
wire n_19118;
wire n_11229;
wire n_4431;
wire n_4192;
wire n_6326;
wire n_18206;
wire n_11919;
wire n_10456;
wire n_18412;
wire n_11675;
wire n_20742;
wire n_21339;
wire n_601;
wire n_14134;
wire n_7979;
wire n_20942;
wire n_172;
wire n_15415;
wire n_19377;
wire n_10979;
wire n_10332;
wire n_18464;
wire n_9443;
wire n_18486;
wire n_6582;
wire n_1658;
wire n_21978;
wire n_19645;
wire n_9897;
wire n_11570;
wire n_176;
wire n_9301;
wire n_6974;
wire n_21690;
wire n_8388;
wire n_16821;
wire n_16701;
wire n_8321;
wire n_1003;
wire n_8091;
wire n_8486;
wire n_19796;
wire n_11592;
wire n_11466;
wire n_5194;
wire n_6898;
wire n_5717;
wire n_19160;
wire n_18059;
wire n_13232;
wire n_17340;
wire n_8841;
wire n_6533;
wire n_3079;
wire n_4965;
wire n_18893;
wire n_5610;
wire n_20097;
wire n_11043;
wire n_8947;
wire n_9671;
wire n_6972;
wire n_4111;
wire n_19747;
wire n_11415;
wire n_2946;
wire n_14773;
wire n_6344;
wire n_5305;
wire n_6093;
wire n_10499;
wire n_15096;
wire n_8093;
wire n_19664;
wire n_19396;
wire n_1117;
wire n_2754;
wire n_10435;
wire n_12220;
wire n_10066;
wire n_13605;
wire n_2012;
wire n_1291;
wire n_21913;
wire n_19872;
wire n_3503;
wire n_8811;
wire n_7150;
wire n_20159;
wire n_7687;
wire n_13599;
wire n_12867;
wire n_18229;
wire n_19504;
wire n_14173;
wire n_3661;
wire n_4878;
wire n_1703;
wire n_14875;
wire n_1137;
wire n_11417;
wire n_19521;
wire n_6988;
wire n_8755;
wire n_12401;
wire n_20998;
wire n_18385;
wire n_21511;
wire n_5897;
wire n_653;
wire n_14777;
wire n_19617;
wire n_15065;
wire n_9809;
wire n_18955;
wire n_16041;
wire n_13518;
wire n_17782;
wire n_19857;
wire n_1999;
wire n_16475;
wire n_13540;
wire n_1372;
wire n_2861;
wire n_18339;
wire n_3943;
wire n_16220;
wire n_10577;
wire n_19243;
wire n_15085;
wire n_8916;
wire n_3293;
wire n_19993;
wire n_17566;
wire n_10037;
wire n_13370;
wire n_16385;
wire n_15844;
wire n_10234;
wire n_21985;
wire n_14801;
wire n_11766;
wire n_7547;
wire n_14802;
wire n_2528;
wire n_4700;
wire n_11457;
wire n_4426;
wire n_17561;
wire n_21375;
wire n_5292;
wire n_2598;
wire n_18910;
wire n_13937;
wire n_14298;
wire n_14623;
wire n_11275;
wire n_14253;
wire n_198;
wire n_8587;
wire n_12337;
wire n_17215;
wire n_10030;
wire n_10676;
wire n_11819;
wire n_18642;
wire n_3431;
wire n_3169;
wire n_11589;
wire n_11309;
wire n_17496;
wire n_19016;
wire n_12927;
wire n_15161;
wire n_15401;
wire n_17227;
wire n_19296;
wire n_11174;
wire n_8646;
wire n_1718;
wire n_4509;
wire n_9866;
wire n_9602;
wire n_509;
wire n_1281;
wire n_19949;
wire n_6219;
wire n_13343;
wire n_18571;
wire n_8315;
wire n_9260;
wire n_16063;
wire n_21653;
wire n_1376;
wire n_2326;
wire n_12048;
wire n_6720;
wire n_8149;
wire n_2188;
wire n_16169;
wire n_186;
wire n_8581;
wire n_16654;
wire n_13932;
wire n_14668;
wire n_1429;
wire n_4644;
wire n_5060;
wire n_17250;
wire n_5334;
wire n_19844;
wire n_7816;
wire n_21140;
wire n_3311;
wire n_7282;
wire n_13198;
wire n_20433;
wire n_19948;
wire n_1861;
wire n_9978;
wire n_16116;
wire n_5731;
wire n_8612;
wire n_5581;
wire n_18308;
wire n_7446;
wire n_16139;
wire n_20743;
wire n_20790;
wire n_17686;
wire n_10171;
wire n_7473;
wire n_20279;
wire n_4435;
wire n_10471;
wire n_6419;
wire n_6039;
wire n_15304;
wire n_11601;
wire n_14400;
wire n_9279;
wire n_8922;
wire n_886;
wire n_1221;
wire n_21606;
wire n_9563;
wire n_7276;
wire n_7351;
wire n_20039;
wire n_3161;
wire n_4827;
wire n_12740;
wire n_7412;
wire n_6436;
wire n_7666;
wire n_12089;
wire n_16328;
wire n_2476;
wire n_10154;
wire n_20013;
wire n_18702;
wire n_5309;
wire n_7901;
wire n_18201;
wire n_19402;
wire n_9980;
wire n_18663;
wire n_18909;
wire n_16476;
wire n_10818;
wire n_4363;
wire n_12721;
wire n_16839;
wire n_21421;
wire n_16681;
wire n_17691;
wire n_15420;
wire n_12541;
wire n_21500;
wire n_4335;
wire n_11849;
wire n_13484;
wire n_6389;
wire n_19020;
wire n_8375;
wire n_10403;
wire n_5764;
wire n_10260;
wire n_9092;
wire n_16870;
wire n_18311;
wire n_16473;
wire n_13438;
wire n_6441;
wire n_10372;
wire n_9283;
wire n_1536;
wire n_13498;
wire n_16842;
wire n_5085;
wire n_20738;
wire n_13661;
wire n_19416;
wire n_21172;
wire n_5950;
wire n_2173;
wire n_17029;
wire n_21845;
wire n_10691;
wire n_16060;
wire n_18579;
wire n_19383;
wire n_19911;
wire n_16864;
wire n_2018;
wire n_13674;
wire n_3245;
wire n_6109;
wire n_499;
wire n_20417;
wire n_12655;
wire n_18957;
wire n_6787;
wire n_796;
wire n_2119;
wire n_2157;
wire n_13133;
wire n_18200;
wire n_21850;
wire n_20736;
wire n_21784;
wire n_740;
wire n_3509;
wire n_3352;
wire n_12862;
wire n_6349;
wire n_20638;
wire n_1061;
wire n_7631;
wire n_15111;
wire n_21362;
wire n_21450;
wire n_16068;
wire n_18365;
wire n_10665;
wire n_10073;
wire n_13251;
wire n_14890;
wire n_8666;
wire n_11873;
wire n_15579;
wire n_8313;
wire n_1487;
wire n_781;
wire n_15149;
wire n_21327;
wire n_17771;
wire n_20913;
wire n_20021;
wire n_13679;
wire n_16648;
wire n_17419;
wire n_20759;
wire n_16402;
wire n_5945;
wire n_13667;
wire n_1739;
wire n_9323;
wire n_10765;
wire n_4835;
wire n_5811;
wire n_21168;
wire n_19932;
wire n_8677;
wire n_12938;
wire n_13772;
wire n_16348;
wire n_5565;
wire n_9540;
wire n_15859;
wire n_20920;
wire n_13033;
wire n_9105;
wire n_13746;
wire n_5643;
wire n_10149;
wire n_14530;
wire n_20941;
wire n_5846;
wire n_13914;
wire n_12722;
wire n_7870;
wire n_17390;
wire n_18691;
wire n_12042;
wire n_20199;
wire n_16671;
wire n_18848;
wire n_6104;
wire n_3373;
wire n_12469;
wire n_16641;
wire n_21392;
wire n_20846;
wire n_16810;
wire n_9574;
wire n_19442;
wire n_20249;
wire n_3726;
wire n_805;
wire n_11050;
wire n_18529;
wire n_17769;
wire n_8238;
wire n_6998;
wire n_10779;
wire n_11789;
wire n_16239;
wire n_7305;
wire n_19745;
wire n_16135;
wire n_10086;
wire n_20015;
wire n_1741;
wire n_11347;
wire n_19472;
wire n_4332;
wire n_17067;
wire n_3347;
wire n_3216;
wire n_7075;
wire n_10869;
wire n_5066;
wire n_6092;
wire n_7275;
wire n_15254;
wire n_4241;
wire n_18176;
wire n_14429;
wire n_14705;
wire n_10128;
wire n_16644;
wire n_20575;
wire n_1186;
wire n_14343;
wire n_14996;
wire n_15072;
wire n_17647;
wire n_14066;
wire n_11989;
wire n_12800;
wire n_12177;
wire n_12036;
wire n_10590;
wire n_12850;
wire n_17378;
wire n_2802;
wire n_17866;
wire n_17210;
wire n_20591;
wire n_3304;
wire n_1378;
wire n_7236;
wire n_15135;
wire n_469;
wire n_7269;
wire n_549;
wire n_20624;
wire n_21755;
wire n_6602;
wire n_4419;
wire n_6502;
wire n_15856;
wire n_13409;
wire n_7326;
wire n_13548;
wire n_7572;
wire n_17062;
wire n_4395;
wire n_12565;
wire n_2821;
wire n_20992;
wire n_9968;
wire n_5074;
wire n_16957;
wire n_2568;
wire n_16950;
wire n_8169;
wire n_15174;
wire n_11958;
wire n_21063;
wire n_20233;
wire n_1021;
wire n_8017;
wire n_5895;
wire n_14756;
wire n_5649;
wire n_5166;
wire n_13255;
wire n_14938;
wire n_2495;
wire n_10785;
wire n_1789;
wire n_21843;
wire n_5457;
wire n_19567;
wire n_15863;
wire n_5532;
wire n_12823;
wire n_18497;
wire n_247;
wire n_12422;
wire n_1494;
wire n_19566;
wire n_11528;
wire n_625;
wire n_18509;
wire n_20592;
wire n_18198;
wire n_7650;
wire n_6525;
wire n_9871;
wire n_6631;
wire n_15162;
wire n_15566;
wire n_4033;
wire n_4289;
wire n_15015;
wire n_4780;
wire n_21586;
wire n_8680;
wire n_4243;
wire n_4982;
wire n_10427;
wire n_3695;
wire n_17136;
wire n_15658;
wire n_6292;
wire n_5544;
wire n_9900;
wire n_3987;
wire n_7339;
wire n_16767;
wire n_14409;
wire n_19278;
wire n_12572;
wire n_6264;
wire n_9608;
wire n_9137;
wire n_12512;
wire n_13736;
wire n_9778;
wire n_8622;
wire n_5410;
wire n_11808;
wire n_3332;
wire n_18253;
wire n_7146;
wire n_3937;
wire n_15819;
wire n_14251;
wire n_8242;
wire n_17920;
wire n_19766;
wire n_14053;
wire n_21081;
wire n_21290;
wire n_7482;
wire n_19721;
wire n_2978;
wire n_8331;
wire n_16887;
wire n_7156;
wire n_3638;
wire n_15438;
wire n_5503;
wire n_1633;
wire n_3763;
wire n_19203;
wire n_3022;
wire n_11695;
wire n_18657;
wire n_21048;
wire n_4264;
wire n_8882;
wire n_3087;
wire n_13583;
wire n_16628;
wire n_9272;
wire n_8708;
wire n_7360;
wire n_12274;
wire n_12348;
wire n_8076;
wire n_11360;
wire n_11886;
wire n_7102;
wire n_8277;
wire n_19496;
wire n_19477;
wire n_13344;
wire n_13336;
wire n_14516;
wire n_15851;
wire n_20903;
wire n_3013;
wire n_14103;
wire n_5654;
wire n_18318;
wire n_10258;
wire n_19507;
wire n_11534;
wire n_1723;
wire n_5999;
wire n_10507;
wire n_19724;
wire n_13885;
wire n_8636;
wire n_4626;
wire n_6637;
wire n_15240;
wire n_798;
wire n_13259;
wire n_21083;
wire n_20174;
wire n_290;
wire n_20735;
wire n_17151;
wire n_6358;
wire n_14737;
wire n_16038;
wire n_16675;
wire n_18711;
wire n_11848;
wire n_8665;
wire n_9086;
wire n_11401;
wire n_9711;
wire n_18651;
wire n_21654;
wire n_13462;
wire n_3985;
wire n_5253;
wire n_21549;
wire n_1391;
wire n_11375;
wire n_4624;
wire n_20486;
wire n_14353;
wire n_9999;
wire n_10814;
wire n_19822;
wire n_813;
wire n_17663;
wire n_6171;
wire n_15366;
wire n_9613;
wire n_4897;
wire n_2769;
wire n_7788;
wire n_858;
wire n_6352;
wire n_13954;
wire n_21190;
wire n_10531;
wire n_7534;
wire n_9462;
wire n_5065;
wire n_10699;
wire n_7032;
wire n_14161;
wire n_3637;
wire n_18345;
wire n_3141;
wire n_10567;
wire n_19816;
wire n_17232;
wire n_5667;
wire n_16120;
wire n_3164;
wire n_10770;
wire n_11693;
wire n_21517;
wire n_4919;
wire n_13584;
wire n_4025;
wire n_16527;
wire n_7634;
wire n_11755;
wire n_20752;
wire n_21588;
wire n_17975;
wire n_7851;
wire n_6332;
wire n_3367;
wire n_13642;
wire n_9573;
wire n_5877;
wire n_19682;
wire n_6306;
wire n_7682;
wire n_3496;
wire n_19768;
wire n_4114;
wire n_14297;
wire n_13618;
wire n_6434;
wire n_12040;
wire n_12443;
wire n_8713;
wire n_17107;
wire n_6751;
wire n_13371;
wire n_12133;
wire n_14048;
wire n_5454;
wire n_7704;
wire n_20791;
wire n_9416;
wire n_8817;
wire n_1581;
wire n_6530;
wire n_15578;
wire n_4089;
wire n_13329;
wire n_16082;
wire n_13788;
wire n_8591;
wire n_21439;
wire n_18686;
wire n_21994;
wire n_6429;
wire n_21631;
wire n_21695;
wire n_3146;
wire n_7239;
wire n_18592;
wire n_963;
wire n_6405;
wire n_11551;
wire n_478;
wire n_18619;
wire n_6613;
wire n_4353;
wire n_2042;
wire n_15584;
wire n_1754;
wire n_20546;
wire n_7821;
wire n_1854;
wire n_5529;
wire n_10248;
wire n_14678;
wire n_19355;
wire n_143;
wire n_16734;
wire n_15224;
wire n_13257;
wire n_17061;
wire n_11976;
wire n_19039;
wire n_13063;
wire n_1906;
wire n_4466;
wire n_15702;
wire n_2262;
wire n_21158;
wire n_13834;
wire n_17827;
wire n_7915;
wire n_8121;
wire n_2945;
wire n_686;
wire n_15624;
wire n_15557;
wire n_16012;
wire n_4688;
wire n_8276;
wire n_17252;
wire n_21204;
wire n_5180;
wire n_13025;
wire n_15923;
wire n_5779;
wire n_6140;
wire n_9039;
wire n_13744;
wire n_9849;
wire n_21935;
wire n_8562;
wire n_3909;
wire n_16838;
wire n_12826;
wire n_6307;
wire n_6164;
wire n_20210;
wire n_18577;
wire n_16262;
wire n_4434;
wire n_15395;
wire n_21469;
wire n_13637;
wire n_10459;
wire n_20684;
wire n_9988;
wire n_5697;
wire n_16566;
wire n_1810;
wire n_7573;
wire n_17631;
wire n_21607;
wire n_7087;
wire n_19518;
wire n_19701;
wire n_21694;
wire n_16619;
wire n_2667;
wire n_11691;
wire n_21763;
wire n_18456;
wire n_9348;
wire n_20750;
wire n_11128;
wire n_21532;
wire n_8226;
wire n_16841;
wire n_12843;
wire n_19540;
wire n_10716;
wire n_12273;
wire n_13701;
wire n_14271;
wire n_11649;
wire n_843;
wire n_13922;
wire n_16707;
wire n_678;
wire n_4184;
wire n_5203;
wire n_17658;
wire n_9356;
wire n_6460;
wire n_1829;
wire n_15388;
wire n_7522;
wire n_19122;
wire n_18393;
wire n_7012;
wire n_11216;
wire n_19632;
wire n_15272;
wire n_17330;
wire n_13553;
wire n_8025;
wire n_1308;
wire n_6383;
wire n_15612;
wire n_16828;
wire n_19095;
wire n_12073;
wire n_15732;
wire n_9516;
wire n_8434;
wire n_17256;
wire n_12848;
wire n_12155;
wire n_13356;
wire n_14286;
wire n_9103;
wire n_18427;
wire n_16801;
wire n_20037;
wire n_16413;
wire n_21242;
wire n_19337;
wire n_2723;
wire n_5672;
wire n_13673;
wire n_20172;
wire n_5601;
wire n_7662;
wire n_14793;
wire n_3855;
wire n_12390;
wire n_12160;
wire n_11297;
wire n_10349;
wire n_20820;
wire n_4931;
wire n_1765;
wire n_18990;
wire n_21284;
wire n_8046;
wire n_19964;
wire n_13897;
wire n_8239;
wire n_4146;
wire n_21028;
wire n_12840;
wire n_8183;
wire n_8924;
wire n_13215;
wire n_20517;
wire n_16026;
wire n_1874;
wire n_2060;
wire n_8848;
wire n_13445;
wire n_10458;
wire n_21937;
wire n_9222;
wire n_15198;
wire n_12994;
wire n_5599;
wire n_18170;
wire n_7186;
wire n_19793;
wire n_8230;
wire n_10478;
wire n_20058;
wire n_21300;
wire n_19679;
wire n_16265;
wire n_8725;
wire n_658;
wire n_2061;
wire n_18817;
wire n_13680;
wire n_16561;
wire n_12951;
wire n_19522;
wire n_20862;
wire n_1586;
wire n_4291;
wire n_11956;
wire n_15996;
wire n_11805;
wire n_12280;
wire n_10698;
wire n_16835;
wire n_8202;
wire n_16852;
wire n_7906;
wire n_19544;
wire n_8678;
wire n_10783;
wire n_20272;
wire n_7658;
wire n_13439;
wire n_8905;
wire n_12051;
wire n_16808;
wire n_3410;
wire n_13789;
wire n_8812;
wire n_21062;
wire n_6828;
wire n_19091;
wire n_14200;
wire n_995;
wire n_19211;
wire n_396;
wire n_8058;
wire n_1073;
wire n_11987;
wire n_5728;
wire n_8394;
wire n_10719;
wire n_9269;
wire n_7835;
wire n_14638;
wire n_21376;
wire n_15326;
wire n_10463;
wire n_13737;
wire n_13441;
wire n_6420;
wire n_21830;
wire n_2882;
wire n_2338;
wire n_19008;
wire n_12384;
wire n_16862;
wire n_12123;
wire n_3197;
wire n_10312;
wire n_18421;
wire n_1043;
wire n_10663;
wire n_5095;
wire n_19113;
wire n_21297;
wire n_21565;
wire n_6754;
wire n_21660;
wire n_6622;
wire n_8747;
wire n_7691;
wire n_10470;
wire n_10563;
wire n_21314;
wire n_2081;
wire n_19187;
wire n_7585;
wire n_4570;
wire n_18316;
wire n_20561;
wire n_12581;
wire n_4296;
wire n_1820;
wire n_7417;
wire n_20697;
wire n_2418;
wire n_18598;
wire n_5841;
wire n_2521;
wire n_9923;
wire n_8224;
wire n_10771;
wire n_20911;
wire n_14556;
wire n_11960;
wire n_6166;
wire n_8628;
wire n_18870;
wire n_11422;
wire n_6781;
wire n_8037;
wire n_8084;
wire n_7120;
wire n_16992;
wire n_21136;
wire n_9801;
wire n_3374;
wire n_17767;
wire n_1870;
wire n_11029;
wire n_18576;
wire n_11199;
wire n_15721;
wire n_13396;
wire n_4600;
wire n_20430;
wire n_1031;
wire n_13652;
wire n_6110;
wire n_6237;
wire n_18767;
wire n_16083;
wire n_834;
wire n_19684;
wire n_19581;
wire n_9330;
wire n_20019;
wire n_15781;
wire n_17512;
wire n_6590;
wire n_9178;
wire n_16646;
wire n_17031;
wire n_10753;
wire n_13965;
wire n_9181;
wire n_7923;
wire n_14465;
wire n_2878;
wire n_6453;
wire n_7559;
wire n_1982;
wire n_20498;
wire n_15476;
wire n_21686;
wire n_10300;
wire n_10257;
wire n_19335;
wire n_12714;
wire n_11166;
wire n_2905;
wire n_18090;
wire n_11217;
wire n_14481;
wire n_3566;
wire n_15650;
wire n_20631;
wire n_19928;
wire n_1084;
wire n_6983;
wire n_7843;
wire n_13774;
wire n_18560;
wire n_10984;
wire n_20925;
wire n_1351;
wire n_17288;
wire n_495;
wire n_17880;
wire n_3486;
wire n_9547;
wire n_11238;
wire n_9895;
wire n_6724;
wire n_2088;
wire n_18199;
wire n_11608;
wire n_21164;
wire n_16407;
wire n_6571;
wire n_19165;
wire n_7470;
wire n_16059;
wire n_9548;
wire n_21475;
wire n_13410;
wire n_20044;
wire n_14432;
wire n_16998;
wire n_21058;
wire n_2656;
wire n_1080;
wire n_9538;
wire n_20390;
wire n_14984;
wire n_13230;
wire n_7597;
wire n_11996;
wire n_6733;
wire n_7071;
wire n_17552;
wire n_15029;
wire n_6035;
wire n_18920;
wire n_1436;
wire n_15967;
wire n_16067;
wire n_1691;
wire n_7109;
wire n_2075;
wire n_3658;
wire n_4807;
wire n_6150;
wire n_9176;
wire n_10461;
wire n_18275;
wire n_20299;
wire n_2131;
wire n_21361;
wire n_1919;
wire n_19997;
wire n_3419;
wire n_13113;
wire n_18819;
wire n_348;
wire n_6016;
wire n_8100;
wire n_2969;
wire n_2864;
wire n_15670;
wire n_3190;
wire n_1553;
wire n_2664;
wire n_14430;
wire n_444;
wire n_8406;
wire n_14697;
wire n_11028;
wire n_5252;
wire n_7009;
wire n_408;
wire n_15847;
wire n_20391;
wire n_21909;
wire n_15708;
wire n_19219;
wire n_2731;
wire n_8693;
wire n_5134;
wire n_3953;
wire n_10207;
wire n_12536;
wire n_11368;
wire n_16962;
wire n_15286;
wire n_7777;
wire n_2998;
wire n_4684;
wire n_15593;
wire n_11404;
wire n_16222;
wire n_7671;
wire n_15951;
wire n_8020;
wire n_20781;
wire n_13866;
wire n_2760;
wire n_3377;
wire n_15129;
wire n_3962;
wire n_5375;
wire n_12362;
wire n_8736;
wire n_16481;
wire n_21507;
wire n_3231;
wire n_10846;
wire n_16356;
wire n_16270;
wire n_621;
wire n_10195;
wire n_11847;
wire n_9718;
wire n_4478;
wire n_21557;
wire n_20420;
wire n_8909;
wire n_19215;
wire n_16033;
wire n_17376;
wire n_11968;
wire n_14127;
wire n_6317;
wire n_9762;
wire n_12903;
wire n_4890;
wire n_5691;
wire n_13103;
wire n_15865;
wire n_15771;
wire n_20496;
wire n_16708;
wire n_17661;
wire n_5647;
wire n_3203;
wire n_14971;
wire n_2903;
wire n_3717;
wire n_13646;
wire n_2743;
wire n_2675;
wire n_9953;
wire n_1439;
wire n_18800;
wire n_14154;
wire n_16332;
wire n_8786;
wire n_12673;
wire n_6734;
wire n_20931;
wire n_21069;
wire n_18923;
wire n_16463;
wire n_9571;
wire n_7135;
wire n_8263;
wire n_8884;
wire n_13062;
wire n_4721;
wire n_5597;
wire n_19233;
wire n_6382;
wire n_7328;
wire n_6404;
wire n_12063;
wire n_10693;
wire n_10493;
wire n_11125;
wire n_10554;
wire n_19966;
wire n_7703;
wire n_4496;
wire n_21751;
wire n_16176;
wire n_13144;
wire n_7277;
wire n_18760;
wire n_21849;
wire n_7265;
wire n_2287;
wire n_11126;
wire n_15958;
wire n_2056;
wire n_10019;
wire n_20248;
wire n_15591;
wire n_15719;
wire n_21529;
wire n_6440;
wire n_9725;
wire n_11953;
wire n_6417;
wire n_20277;
wire n_1735;
wire n_16503;
wire n_833;
wire n_8177;
wire n_14013;
wire n_15385;
wire n_20776;
wire n_18094;
wire n_12062;
wire n_12636;
wire n_2504;
wire n_4495;
wire n_5942;
wire n_21670;
wire n_16522;
wire n_9084;
wire n_7728;
wire n_3442;
wire n_17638;
wire n_10767;
wire n_1201;
wire n_7219;
wire n_11040;
wire n_11751;
wire n_4141;
wire n_669;
wire n_10579;
wire n_15296;
wire n_15586;
wire n_1020;
wire n_7805;
wire n_20673;
wire n_21808;
wire n_9973;
wire n_211;
wire n_19380;
wire n_1917;
wire n_16303;
wire n_2325;
wire n_8320;
wire n_15458;
wire n_12157;
wire n_2446;
wire n_18027;
wire n_11182;
wire n_10587;
wire n_19312;
wire n_7182;
wire n_4547;
wire n_2893;
wire n_4004;
wire n_2962;
wire n_10843;
wire n_6484;
wire n_661;
wire n_7674;
wire n_10755;
wire n_5466;
wire n_13645;
wire n_12649;
wire n_1786;
wire n_8370;
wire n_11908;
wire n_7951;
wire n_15190;
wire n_19839;
wire n_2080;
wire n_3552;
wire n_875;
wire n_357;
wire n_12696;
wire n_6717;
wire n_13505;
wire n_165;
wire n_8395;
wire n_11745;
wire n_13181;
wire n_10682;
wire n_5530;
wire n_12940;
wire n_19162;
wire n_6196;
wire n_15608;
wire n_21486;
wire n_18444;
wire n_18269;
wire n_10236;
wire n_1702;
wire n_5221;
wire n_6992;
wire n_20295;
wire n_4183;
wire n_12312;
wire n_15191;
wire n_10303;
wire n_3764;
wire n_11452;
wire n_15270;
wire n_19137;
wire n_19497;
wire n_5311;
wire n_2649;
wire n_7892;
wire n_11558;
wire n_17670;
wire n_9165;
wire n_21510;
wire n_13018;
wire n_13185;
wire n_14681;
wire n_15171;
wire n_21969;
wire n_18540;
wire n_5575;
wire n_7990;
wire n_7626;
wire n_10855;
wire n_8748;
wire n_4819;
wire n_11429;
wire n_7088;
wire n_6519;
wire n_16412;
wire n_1541;
wire n_4900;
wire n_8120;
wire n_6414;
wire n_1713;
wire n_1737;
wire n_10059;
wire n_10284;
wire n_4930;
wire n_5276;
wire n_6308;
wire n_14790;
wire n_6906;
wire n_14029;
wire n_19147;
wire n_6629;
wire n_18707;
wire n_16393;
wire n_17909;
wire n_4070;
wire n_11124;
wire n_665;
wire n_3839;
wire n_12734;
wire n_14032;
wire n_14760;
wire n_4659;
wire n_6188;
wire n_17727;
wire n_18915;
wire n_19264;
wire n_4579;
wire n_20773;
wire n_13709;
wire n_3014;
wire n_6398;
wire n_11586;
wire n_14660;
wire n_5023;
wire n_20075;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_18877;
wire n_9064;
wire n_3530;
wire n_18326;
wire n_14056;
wire n_2765;
wire n_3329;
wire n_18155;
wire n_10200;
wire n_12442;
wire n_14588;
wire n_2003;
wire n_12499;
wire n_9383;
wire n_10290;
wire n_15853;
wire n_15862;
wire n_16358;
wire n_13684;
wire n_18458;
wire n_6231;
wire n_11036;
wire n_872;
wire n_18420;
wire n_14826;
wire n_11927;
wire n_1297;
wire n_21043;
wire n_10306;
wire n_19503;
wire n_20628;
wire n_15445;
wire n_1972;
wire n_7862;
wire n_18373;
wire n_2806;
wire n_2184;
wire n_5312;
wire n_17933;
wire n_9986;
wire n_10355;
wire n_14967;
wire n_11118;
wire n_3249;
wire n_12496;
wire n_17347;
wire n_20137;
wire n_676;
wire n_15028;
wire n_15736;
wire n_194;
wire n_21787;
wire n_5687;
wire n_12479;
wire n_13703;
wire n_10999;
wire n_18929;
wire n_18689;
wire n_10899;
wire n_15573;
wire n_19827;
wire n_16620;
wire n_21299;
wire n_2332;
wire n_15097;
wire n_11561;
wire n_12345;
wire n_15126;
wire n_21325;
wire n_1227;
wire n_3600;
wire n_4134;
wire n_20938;
wire n_10425;
wire n_8352;
wire n_21457;
wire n_8385;
wire n_8166;
wire n_19652;
wire n_581;
wire n_11433;
wire n_2130;
wire n_2773;
wire n_17843;
wire n_17090;
wire n_1452;
wire n_5612;
wire n_6125;
wire n_15213;
wire n_4251;
wire n_6560;
wire n_14686;
wire n_17747;
wire n_1326;
wire n_10711;
wire n_8659;
wire n_20483;
wire n_8804;
wire n_19498;
wire n_16460;
wire n_2186;
wire n_8439;
wire n_18627;
wire n_21348;
wire n_8369;
wire n_11574;
wire n_18771;
wire n_5007;
wire n_16937;
wire n_2562;
wire n_7615;
wire n_1192;
wire n_15238;
wire n_19438;
wire n_21659;
wire n_3862;
wire n_5563;
wire n_5487;
wire n_6593;
wire n_19834;
wire n_2348;
wire n_6673;
wire n_7172;
wire n_10685;
wire n_5497;
wire n_8234;
wire n_18873;
wire n_18041;
wire n_21330;
wire n_7112;
wire n_16217;
wire n_19989;
wire n_8989;
wire n_13589;
wire n_16625;
wire n_14192;
wire n_3584;
wire n_3756;
wire n_381;
wire n_13481;
wire n_390;
wire n_13743;
wire n_17759;
wire n_2772;
wire n_19942;
wire n_5444;
wire n_14365;
wire n_20284;
wire n_3999;
wire n_8534;
wire n_2844;
wire n_9911;
wire n_6559;
wire n_10302;
wire n_1813;
wire n_7144;
wire n_4833;
wire n_14244;
wire n_13357;
wire n_6841;
wire n_16252;
wire n_14918;
wire n_11002;
wire n_16631;
wire n_6653;
wire n_16045;
wire n_2382;
wire n_4719;
wire n_21095;
wire n_2317;
wire n_5425;
wire n_17015;
wire n_1973;
wire n_8042;
wire n_15108;
wire n_11474;
wire n_20208;
wire n_4401;
wire n_1756;
wire n_21196;
wire n_8839;
wire n_6112;
wire n_2788;
wire n_11738;
wire n_2984;
wire n_6198;
wire n_18243;
wire n_15483;
wire n_12074;
wire n_17353;
wire n_11931;
wire n_15841;
wire n_10925;
wire n_14508;
wire n_8758;
wire n_622;
wire n_5666;
wire n_13508;
wire n_13058;
wire n_17242;
wire n_17588;
wire n_7227;
wire n_4605;
wire n_15042;
wire n_8511;
wire n_3235;
wire n_21552;
wire n_6756;
wire n_8595;
wire n_1272;
wire n_12900;
wire n_8873;
wire n_7096;
wire n_19339;
wire n_17918;
wire n_17150;
wire n_3903;
wire n_10102;
wire n_1210;
wire n_10908;
wire n_21423;
wire n_4158;
wire n_6015;
wire n_3254;
wire n_5683;
wire n_4171;
wire n_13503;
wire n_18322;
wire n_12595;
wire n_18246;
wire n_9400;
wire n_4045;
wire n_598;
wire n_3634;
wire n_16528;
wire n_2531;
wire n_10936;
wire n_17934;
wire n_413;
wire n_7485;
wire n_15673;
wire n_203;
wire n_10440;
wire n_10630;
wire n_8336;
wire n_16493;
wire n_4979;
wire n_21675;
wire n_19149;
wire n_2234;
wire n_14404;
wire n_6553;
wire n_7808;
wire n_1255;
wire n_9859;
wire n_9003;
wire n_13849;
wire n_722;
wire n_6628;
wire n_844;
wire n_3497;
wire n_20183;
wire n_5409;
wire n_7536;
wire n_20317;
wire n_17087;
wire n_20865;
wire n_4566;
wire n_9597;
wire n_6293;
wire n_8417;
wire n_9076;
wire n_18643;
wire n_8498;
wire n_7991;
wire n_7676;
wire n_11769;
wire n_19195;
wire n_12486;
wire n_585;
wire n_7553;
wire n_12623;
wire n_13698;
wire n_6381;
wire n_19889;
wire n_5307;
wire n_20266;
wire n_14122;
wire n_4328;
wire n_21962;
wire n_7095;
wire n_11794;
wire n_5415;
wire n_8880;
wire n_6577;
wire n_20346;
wire n_18189;
wire n_20010;
wire n_3175;
wire n_14546;
wire n_18262;
wire n_18236;
wire n_20096;
wire n_4429;
wire n_13079;
wire n_4591;
wire n_10500;
wire n_9805;
wire n_7210;
wire n_4646;
wire n_5769;
wire n_21202;
wire n_16051;
wire n_18134;
wire n_18298;
wire n_11428;
wire n_3247;
wire n_3091;
wire n_6309;
wire n_9520;
wire n_246;
wire n_12925;
wire n_20945;
wire n_7723;
wire n_6527;
wire n_10550;
wire n_20851;
wire n_9583;
wire n_18585;
wire n_13622;
wire n_9036;
wire n_13145;
wire n_19717;
wire n_5979;
wire n_19580;
wire n_565;
wire n_5089;
wire n_14394;
wire n_17935;
wire n_16008;
wire n_20124;
wire n_1505;
wire n_6929;
wire n_21821;
wire n_14256;
wire n_21685;
wire n_11339;
wire n_651;
wire n_4636;
wire n_807;
wire n_4711;
wire n_12986;
wire n_13570;
wire n_10254;
wire n_3335;
wire n_20389;
wire n_3413;
wire n_15589;
wire n_8912;
wire n_2689;
wire n_18665;
wire n_4191;
wire n_16548;
wire n_4293;
wire n_8227;
wire n_21895;
wire n_21025;
wire n_3414;
wire n_14846;
wire n_17877;
wire n_7456;
wire n_13459;
wire n_21391;
wire n_10657;
wire n_13899;
wire n_9798;
wire n_17115;
wire n_18896;
wire n_16251;
wire n_15677;
wire n_15487;
wire n_1161;
wire n_19125;
wire n_11318;
wire n_3027;
wire n_3732;
wire n_21503;
wire n_4250;
wire n_5329;
wire n_8358;
wire n_9410;
wire n_880;
wire n_3297;
wire n_13594;
wire n_13991;
wire n_7909;
wire n_15133;
wire n_2683;
wire n_1360;
wire n_12278;
wire n_4854;
wire n_14428;
wire n_17028;
wire n_11850;
wire n_8396;
wire n_9838;
wire n_688;
wire n_7780;
wire n_17454;
wire n_3350;
wire n_17936;
wire n_2389;
wire n_7444;
wire n_11468;
wire n_4038;
wire n_5297;
wire n_915;
wire n_20378;
wire n_20088;
wire n_19242;
wire n_6816;
wire n_9752;
wire n_21874;
wire n_12540;
wire n_7049;
wire n_497;
wire n_13080;
wire n_16340;
wire n_6879;
wire n_17653;
wire n_1686;
wire n_947;
wire n_373;
wire n_21387;
wire n_6702;
wire n_16512;
wire n_14682;
wire n_4144;
wire n_15921;
wire n_5774;
wire n_929;
wire n_14527;
wire n_12619;
wire n_8792;
wire n_16953;
wire n_5131;
wire n_1576;
wire n_1182;
wire n_18232;
wire n_11870;
wire n_11186;
wire n_17720;
wire n_20064;
wire n_16519;
wire n_11233;
wire n_15193;
wire n_16264;
wire n_3258;
wire n_18233;
wire n_20382;
wire n_14726;
wire n_4989;
wire n_4622;
wire n_13511;
wire n_10786;
wire n_9598;
wire n_8382;
wire n_8971;
wire n_10602;
wire n_13699;
wire n_17657;
wire n_2983;
wire n_11878;
wire n_227;
wire n_19021;
wire n_2715;
wire n_6132;
wire n_6578;
wire n_1669;
wire n_16831;
wire n_12870;
wire n_5342;
wire n_19667;
wire n_2672;
wire n_12911;
wire n_19569;
wire n_19024;
wire n_6918;
wire n_1374;
wire n_4793;
wire n_9833;
wire n_11837;
wire n_6612;
wire n_4168;
wire n_12651;
wire n_7863;
wire n_5680;
wire n_1146;
wire n_8633;
wire n_5838;
wire n_897;
wire n_10969;
wire n_6375;
wire n_16680;
wire n_13825;
wire n_13798;
wire n_1872;
wire n_3389;
wire n_12304;
wire n_9698;
wire n_12270;
wire n_9124;
wire n_9695;
wire n_1070;
wire n_6447;
wire n_9497;
wire n_5206;
wire n_15983;
wire n_8479;
wire n_3222;
wire n_12210;
wire n_17442;
wire n_14525;
wire n_1801;
wire n_14058;
wire n_20694;
wire n_6130;
wire n_12858;
wire n_20251;
wire n_21431;
wire n_837;
wire n_15018;
wire n_2791;
wire n_3755;
wire n_8179;
wire n_15825;
wire n_5803;
wire n_14272;
wire n_16399;
wire n_21454;
wire n_7530;
wire n_2174;
wire n_2506;
wire n_4064;
wire n_16300;
wire n_10692;
wire n_1863;
wire n_20767;
wire n_8733;
wire n_11723;
wire n_2407;
wire n_16811;
wire n_9652;
wire n_5058;
wire n_12653;
wire n_19728;
wire n_18534;
wire n_6119;
wire n_11949;
wire n_1322;
wire n_15004;
wire n_889;
wire n_2358;
wire n_5192;
wire n_21728;
wire n_5141;
wire n_14743;
wire n_11880;
wire n_3252;
wire n_10385;
wire n_3544;
wire n_11377;
wire n_11302;
wire n_6338;
wire n_1523;
wire n_12425;
wire n_14922;
wire n_15181;
wire n_18423;
wire n_15211;
wire n_8425;
wire n_10809;
wire n_9349;
wire n_4908;
wire n_8241;
wire n_736;
wire n_16851;
wire n_18085;
wire n_19973;
wire n_7932;
wire n_11626;
wire n_14957;
wire n_5730;
wire n_11694;
wire n_13811;
wire n_1278;
wire n_19663;
wire n_16109;
wire n_18625;
wire n_16359;
wire n_2784;
wire n_7541;
wire n_4862;
wire n_17628;
wire n_2557;
wire n_1248;
wire n_10973;
wire n_18183;
wire n_12015;
wire n_289;
wire n_6625;
wire n_3781;
wire n_12135;
wire n_17284;
wire n_6302;
wire n_21449;
wire n_5748;
wire n_2942;
wire n_5525;
wire n_8152;
wire n_10526;
wire n_21182;
wire n_7636;
wire n_17086;
wire n_4224;
wire n_6483;
wire n_8829;
wire n_20103;
wire n_17698;
wire n_12869;
wire n_15764;
wire n_17268;
wire n_13841;
wire n_857;
wire n_18110;
wire n_14344;
wire n_19525;
wire n_16181;
wire n_20505;
wire n_12059;
wire n_20312;
wire n_20250;
wire n_20114;
wire n_1951;
wire n_1883;
wire n_13043;
wire n_13960;
wire n_10221;
wire n_4702;
wire n_14069;
wire n_17364;
wire n_10109;
wire n_18469;
wire n_15875;
wire n_10928;
wire n_971;
wire n_19620;
wire n_9024;
wire n_9523;
wire n_404;
wire n_16074;
wire n_21782;
wire n_20999;
wire n_5139;
wire n_13260;
wire n_6922;
wire n_14474;
wire n_9679;
wire n_9000;
wire n_9742;
wire n_20024;
wire n_2679;
wire n_21963;
wire n_19789;
wire n_6651;
wire n_7296;
wire n_14704;
wire n_7273;
wire n_18608;
wire n_266;
wire n_2930;
wire n_2777;
wire n_2434;
wire n_2660;
wire n_14675;
wire n_10600;
wire n_17533;
wire n_11056;
wire n_21896;
wire n_17726;
wire n_11774;
wire n_8627;
wire n_2698;
wire n_5043;
wire n_1481;
wire n_18043;
wire n_13910;
wire n_13369;
wire n_12099;
wire n_868;
wire n_2454;
wire n_15077;
wire n_4371;
wire n_4268;
wire n_12191;
wire n_19777;
wire n_3895;
wire n_17836;
wire n_17993;
wire n_5585;
wire n_6397;
wire n_19426;
wire n_4427;
wire n_14221;
wire n_6121;
wire n_16010;
wire n_4142;
wire n_1189;
wire n_9858;
wire n_4260;
wire n_20421;
wire n_18903;
wire n_11157;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_14932;
wire n_20565;
wire n_6954;
wire n_3279;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_523;
wire n_1537;
wire n_13417;
wire n_14350;
wire n_4262;
wire n_8362;
wire n_1798;
wire n_10344;
wire n_7131;
wire n_7769;
wire n_10882;
wire n_9303;
wire n_525;
wire n_15971;
wire n_11220;
wire n_14220;
wire n_21848;
wire n_14451;
wire n_8491;
wire n_9058;
wire n_6941;
wire n_17778;
wire n_17212;
wire n_2073;
wire n_5515;
wire n_8324;
wire n_14510;
wire n_17506;
wire n_7418;
wire n_20705;
wire n_5250;
wire n_3144;
wire n_18899;
wire n_21976;
wire n_10518;
wire n_21250;
wire n_20824;
wire n_1615;
wire n_19681;
wire n_2005;
wire n_526;
wire n_1916;
wire n_20823;
wire n_15447;
wire n_11481;
wire n_11712;
wire n_8625;
wire n_20304;
wire n_7204;
wire n_8180;
wire n_689;
wire n_1624;
wire n_4970;
wire n_640;
wire n_9062;
wire n_14606;
wire n_1279;
wire n_19718;
wire n_4108;
wire n_15510;
wire n_1090;
wire n_16086;
wire n_10486;
wire n_19934;
wire n_21175;
wire n_758;
wire n_16967;
wire n_16047;
wire n_20061;
wire n_19364;
wire n_13797;
wire n_7925;
wire n_1068;
wire n_2580;
wire n_15351;
wire n_9065;
wire n_11650;
wire n_5163;
wire n_17881;
wire n_18754;
wire n_21936;
wire n_5768;
wire n_3753;
wire n_7640;
wire n_8187;
wire n_3579;
wire n_18975;
wire n_7422;
wire n_7920;
wire n_9431;
wire n_10167;
wire n_9160;
wire n_20287;
wire n_17671;
wire n_152;
wire n_10442;
wire n_12829;
wire n_17026;
wire n_18242;
wire n_9808;
wire n_19419;
wire n_10534;
wire n_19093;
wire n_21703;
wire n_10406;
wire n_8316;
wire n_19662;
wire n_12783;
wire n_1017;
wire n_9184;
wire n_16813;
wire n_2116;
wire n_1054;
wire n_12631;
wire n_10965;
wire n_1828;
wire n_2320;
wire n_7175;
wire n_2137;
wire n_4973;
wire n_18370;
wire n_16748;
wire n_19862;
wire n_13964;
wire n_2583;
wire n_17183;
wire n_9207;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_18330;
wire n_19358;
wire n_5216;
wire n_18499;
wire n_17610;
wire n_20710;
wire n_16250;
wire n_9010;
wire n_4170;
wire n_14754;
wire n_11747;
wire n_3719;
wire n_7855;
wire n_10371;
wire n_3681;
wire n_12675;
wire n_2737;
wire n_12174;
wire n_4308;
wire n_2812;
wire n_17560;
wire n_15747;
wire n_12113;
wire n_15516;
wire n_1426;
wire n_19444;
wire n_8162;
wire n_2725;
wire n_21306;
wire n_6949;
wire n_14198;
wire n_21329;
wire n_7260;
wire n_13820;
wire n_12470;
wire n_14039;
wire n_8546;
wire n_9878;
wire n_18821;
wire n_208;
wire n_20598;
wire n_15323;
wire n_7263;
wire n_17992;
wire n_3149;
wire n_9674;
wire n_17121;
wire n_18143;
wire n_12799;
wire n_20315;
wire n_4200;
wire n_19509;
wire n_21828;
wire n_3466;
wire n_13976;
wire n_20188;
wire n_14862;
wire n_18745;
wire n_15833;
wire n_19260;
wire n_10960;
wire n_4271;
wire n_7509;
wire n_11620;
wire n_5171;
wire n_12617;
wire n_12919;
wire n_7240;
wire n_19614;
wire n_4071;
wire n_15933;
wire n_16591;
wire n_19812;
wire n_20255;
wire n_14005;
wire n_263;
wire n_10896;
wire n_8767;
wire n_16890;
wire n_13764;
wire n_2681;
wire n_17217;
wire n_11851;
wire n_16545;
wire n_4922;
wire n_7609;
wire n_19579;
wire n_14688;
wire n_8010;
wire n_7278;
wire n_12637;
wire n_1651;
wire n_17254;
wire n_12301;
wire n_8347;
wire n_14468;
wire n_2775;
wire n_19804;
wire n_6416;
wire n_4693;
wire n_5488;
wire n_21563;
wire n_18961;
wire n_17291;
wire n_16370;
wire n_8204;
wire n_14067;
wire n_3557;
wire n_7741;
wire n_20625;
wire n_4744;
wire n_7565;
wire n_11259;
wire n_20966;
wire n_11197;
wire n_15635;
wire n_174;
wire n_15403;
wire n_17171;
wire n_12977;
wire n_441;
wire n_7097;
wire n_13227;
wire n_2204;
wire n_6421;
wire n_7414;
wire n_10660;
wire n_20239;
wire n_20487;
wire n_13166;
wire n_365;
wire n_8312;
wire n_18449;
wire n_14242;
wire n_11153;
wire n_729;
wire n_4964;
wire n_21743;
wire n_6192;
wire n_20424;
wire n_13266;
wire n_21332;
wire n_13319;
wire n_13623;
wire n_15062;
wire n_12436;
wire n_20343;
wire n_12528;
wire n_20462;
wire n_19246;
wire n_14586;
wire n_5437;
wire n_623;
wire n_15959;
wire n_5826;
wire n_7659;
wire n_3881;
wire n_14095;
wire n_4583;
wire n_233;
wire n_16354;
wire n_17984;
wire n_6662;
wire n_5245;
wire n_7189;
wire n_8688;
wire n_4666;
wire n_10740;
wire n_17172;
wire n_16108;
wire n_10558;
wire n_8116;
wire n_12144;
wire n_10297;
wire n_13981;
wire n_4540;
wire n_21260;
wire n_16216;
wire n_4891;
wire n_8519;
wire n_19685;
wire n_15620;
wire n_17725;
wire n_1023;
wire n_17883;
wire n_3559;
wire n_15717;
wire n_11647;
wire n_12392;
wire n_2661;
wire n_13205;
wire n_18578;
wire n_17037;
wire n_5716;
wire n_19360;
wire n_18545;
wire n_3588;
wire n_21965;
wire n_2308;
wire n_7492;
wire n_19657;
wire n_13730;
wire n_15087;
wire n_12665;
wire n_5231;
wire n_7809;
wire n_19252;
wire n_3860;
wire n_1029;
wire n_12067;
wire n_19373;
wire n_12546;
wire n_2191;
wire n_13489;
wire n_10007;
wire n_10904;
wire n_2428;
wire n_3847;
wire n_9961;
wire n_18673;
wire n_2158;
wire n_11325;
wire n_5390;
wire n_14612;
wire n_2824;
wire n_20169;
wire n_19105;
wire n_16190;
wire n_3665;
wire n_20771;
wire n_20109;
wire n_20899;
wire n_5833;
wire n_3800;
wire n_9593;
wire n_20780;
wire n_18149;
wire n_14765;
wire n_2792;
wire n_18346;
wire n_20203;
wire n_19300;
wire n_3991;
wire n_3134;
wire n_11025;
wire n_19392;
wire n_4172;
wire n_13117;
wire n_13510;
wire n_17977;
wire n_13665;
wire n_17190;
wire n_5149;
wire n_16441;
wire n_4611;
wire n_14835;
wire n_2294;
wire n_19067;
wire n_455;
wire n_5135;
wire n_16092;
wire n_2948;
wire n_2309;
wire n_15025;
wire n_20599;
wire n_5494;
wire n_19090;
wire n_21446;
wire n_6200;
wire n_2123;
wire n_11437;
wire n_2685;
wire n_17022;
wire n_4422;
wire n_10902;
wire n_18661;
wire n_18453;
wire n_20186;
wire n_12487;
wire n_13861;
wire n_15471;
wire n_16977;
wire n_9320;
wire n_4555;
wire n_5136;
wire n_15451;
wire n_14580;
wire n_153;
wire n_14654;
wire n_3956;
wire n_13081;
wire n_4280;
wire n_9526;
wire n_8107;
wire n_842;
wire n_7642;
wire n_15993;
wire n_2082;
wire n_7045;
wire n_12646;
wire n_11665;
wire n_15880;
wire n_17458;
wire n_13444;
wire n_9692;
wire n_13267;
wire n_15737;
wire n_16437;
wire n_9141;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_9787;
wire n_8674;
wire n_13362;
wire n_21817;
wire n_7931;
wire n_12061;
wire n_12380;
wire n_18768;
wire n_323;
wire n_3253;
wire n_21714;
wire n_8899;
wire n_11127;
wire n_2280;
wire n_9015;
wire n_21014;
wire n_6796;
wire n_3689;
wire n_11632;
wire n_20410;
wire n_21753;
wire n_11762;
wire n_11843;
wire n_17109;
wire n_9389;
wire n_1616;
wire n_12247;
wire n_16435;
wire n_10129;
wire n_3869;
wire n_5042;
wire n_10084;
wire n_20588;
wire n_21385;
wire n_2810;
wire n_21864;
wire n_10318;
wire n_13785;
wire n_14665;
wire n_18649;
wire n_8561;
wire n_10877;
wire n_2126;
wire n_19307;
wire n_17859;
wire n_6281;
wire n_21626;
wire n_9381;
wire n_4079;
wire n_4091;
wire n_13634;
wire n_1638;
wire n_9873;
wire n_15738;
wire n_16636;
wire n_21483;
wire n_9575;
wire n_11817;
wire n_15887;
wire n_6094;
wire n_2935;
wire n_16941;
wire n_5191;
wire n_10298;
wire n_18408;
wire n_6240;
wire n_5293;
wire n_1358;
wire n_10293;
wire n_4316;
wire n_15228;
wire n_20291;
wire n_10432;
wire n_2638;
wire n_15192;
wire n_7515;
wire n_4062;
wire n_13191;
wire n_4843;
wire n_10640;
wire n_11546;
wire n_19061;
wire n_7894;
wire n_20325;
wire n_1506;
wire n_15045;
wire n_9029;
wire n_16455;
wire n_567;
wire n_12262;
wire n_6721;
wire n_8178;
wire n_2608;
wire n_13452;
wire n_20774;
wire n_16733;
wire n_2392;
wire n_14138;
wire n_16040;
wire n_21281;
wire n_10130;
wire n_2835;
wire n_6260;
wire n_16515;
wire n_1968;
wire n_10214;
wire n_3269;
wire n_19826;
wire n_19770;
wire n_12658;
wire n_11389;
wire n_17766;
wire n_7566;
wire n_7937;
wire n_7055;
wire n_3605;
wire n_16401;
wire n_10491;
wire n_20149;
wire n_10712;
wire n_17287;
wire n_4115;
wire n_726;
wire n_21534;
wire n_21274;
wire n_11034;
wire n_2766;
wire n_18520;
wire n_2201;
wire n_14062;
wire n_16235;
wire n_20712;
wire n_1957;
wire n_7954;
wire n_3226;
wire n_6570;
wire n_10062;
wire n_14553;
wire n_17930;
wire n_937;
wire n_2779;
wire n_487;
wire n_19742;
wire n_10216;
wire n_14377;
wire n_8386;
wire n_2115;
wire n_18441;
wire n_20405;
wire n_5327;
wire n_10431;
wire n_6045;
wire n_21871;
wire n_19200;
wire n_1302;
wire n_18666;
wire n_14776;
wire n_9220;
wire n_17255;
wire n_9834;
wire n_2811;
wire n_19199;
wire n_14551;
wire n_15001;
wire n_6489;
wire n_14449;
wire n_14919;
wire n_20893;
wire n_1803;
wire n_15535;
wire n_9642;
wire n_14768;
wire n_9020;
wire n_1991;
wire n_2224;
wire n_20152;
wire n_6806;
wire n_11439;
wire n_14744;
wire n_11752;
wire n_14081;
wire n_4743;
wire n_16287;
wire n_17941;
wire n_148;
wire n_15861;
wire n_4859;
wire n_9940;
wire n_20788;
wire n_7058;
wire n_6284;
wire n_21322;
wire n_8503;
wire n_19760;
wire n_19189;
wire n_9198;
wire n_4733;
wire n_11729;
wire n_3871;
wire n_11699;
wire n_7735;
wire n_8265;
wire n_1689;
wire n_20885;
wire n_1855;
wire n_11902;
wire n_401;
wire n_15716;
wire n_10080;
wire n_2199;
wire n_17264;
wire n_12344;
wire n_8937;
wire n_12961;
wire n_8272;
wire n_3285;
wire n_9249;
wire n_15527;
wire n_294;
wire n_12193;
wire n_21839;
wire n_15748;
wire n_2228;
wire n_14033;
wire n_4551;
wire n_13393;
wire n_684;
wire n_20902;
wire n_18218;
wire n_2902;
wire n_2480;
wire n_6034;
wire n_16627;
wire n_15032;
wire n_7499;
wire n_17253;
wire n_17972;
wire n_20127;
wire n_17298;
wire n_11006;
wire n_6762;
wire n_20739;
wire n_7895;
wire n_13250;
wire n_17655;
wire n_18996;
wire n_7391;
wire n_3711;
wire n_10890;
wire n_12093;
wire n_5837;
wire n_4436;
wire n_17276;
wire n_18462;
wire n_12705;
wire n_719;
wire n_17342;
wire n_8728;
wire n_12241;
wire n_6005;
wire n_21953;
wire n_1530;
wire n_20205;
wire n_3131;
wire n_19232;
wire n_21525;
wire n_15402;
wire n_16124;
wire n_20392;
wire n_5793;
wire n_5591;
wire n_21625;
wire n_13237;
wire n_508;
wire n_986;
wire n_19927;
wire n_21704;
wire n_1317;
wire n_9784;
wire n_2102;
wire n_1063;
wire n_21934;
wire n_10217;
wire n_12231;
wire n_4853;
wire n_12745;
wire n_15474;
wire n_20809;
wire n_15768;
wire n_9101;
wire n_15955;
wire n_6213;
wire n_18966;
wire n_10393;
wire n_18537;
wire n_2239;
wire n_12527;
wire n_16584;
wire n_21554;
wire n_19661;
wire n_14386;
wire n_8897;
wire n_3852;
wire n_812;
wire n_4520;
wire n_13913;
wire n_12354;
wire n_16078;
wire n_5507;
wire n_18023;
wire n_7214;
wire n_12886;
wire n_13564;
wire n_7408;
wire n_9250;
wire n_6115;
wire n_20726;
wire n_9572;
wire n_10375;
wire n_17006;
wire n_9483;
wire n_9816;
wire n_9253;
wire n_15080;
wire n_16981;
wire n_9136;
wire n_2710;
wire n_8357;
wire n_10726;
wire n_1745;
wire n_20864;
wire n_14017;
wire n_4571;
wire n_13434;
wire n_18603;
wire n_6430;
wire n_16510;
wire n_15916;
wire n_3439;
wire n_13657;
wire n_10002;
wire n_6822;
wire n_14639;
wire n_2535;
wire n_4205;
wire n_7599;
wire n_570;
wire n_20880;
wire n_20769;
wire n_5277;
wire n_20102;
wire n_15258;
wire n_9767;
wire n_19230;
wire n_16085;
wire n_6797;
wire n_11367;
wire n_2799;
wire n_4454;
wire n_5952;
wire n_21928;
wire n_2376;
wire n_10251;
wire n_787;
wire n_11562;
wire n_17159;
wire n_18925;
wire n_17194;
wire n_12854;
wire n_21604;
wire n_20704;
wire n_9949;
wire n_18319;
wire n_18881;
wire n_4879;
wire n_9684;
wire n_15418;
wire n_6152;
wire n_13430;
wire n_8243;
wire n_4221;
wire n_11117;
wire n_11046;
wire n_17614;
wire n_14901;
wire n_386;
wire n_13327;
wire n_1550;
wire n_5777;
wire n_20662;
wire n_10475;
wire n_21947;
wire n_141;
wire n_14195;
wire n_3102;
wire n_1648;
wire n_19068;
wire n_10467;
wire n_5156;
wire n_5926;
wire n_19235;
wire n_9399;
wire n_3551;
wire n_17393;
wire n_17544;
wire n_17522;
wire n_12506;
wire n_140;
wire n_15104;
wire n_3859;
wire n_3722;
wire n_21124;
wire n_928;
wire n_13844;
wire n_14462;
wire n_1943;
wire n_15773;
wire n_11934;
wire n_15638;
wire n_9013;
wire n_9290;
wire n_3351;
wire n_13342;
wire n_7698;
wire n_12884;
wire n_13187;
wire n_7344;
wire n_1348;
wire n_2883;
wire n_9586;
wire n_10751;
wire n_4825;
wire n_4549;
wire n_12502;
wire n_9104;
wire n_10225;
wire n_15517;
wire n_10570;
wire n_9293;
wire n_16987;
wire n_13298;
wire n_16504;
wire n_5470;
wire n_16174;
wire n_4565;
wire n_7675;
wire n_4039;
wire n_3227;
wire n_16949;
wire n_4574;
wire n_17511;
wire n_6696;
wire n_5222;
wire n_9919;
wire n_8826;
wire n_20907;
wire n_8715;
wire n_12761;
wire n_595;
wire n_14522;
wire n_6117;
wire n_632;
wire n_4231;
wire n_8117;
wire n_3652;
wire n_12822;
wire n_14148;
wire n_18804;
wire n_6681;
wire n_13539;
wire n_161;
wire n_15892;
wire n_1937;
wire n_11420;
wire n_21046;
wire n_11470;
wire n_8497;
wire n_12082;
wire n_745;
wire n_12151;
wire n_7940;
wire n_14493;
wire n_11230;
wire n_15468;
wire n_17459;
wire n_7606;
wire n_4939;
wire n_14534;
wire n_6896;
wire n_12183;
wire n_11669;
wire n_10734;
wire n_17174;
wire n_8798;
wire n_20973;
wire n_21005;
wire n_16128;
wire n_2404;
wire n_19511;
wire n_7884;
wire n_17668;
wire n_8502;
wire n_13293;
wire n_1936;
wire n_16465;
wire n_14487;
wire n_10445;
wire n_15241;
wire n_19994;
wire n_5974;
wire n_9298;
wire n_6438;
wire n_20509;
wire n_1402;
wire n_13285;
wire n_6316;
wire n_18315;
wire n_16711;
wire n_1397;
wire n_21730;
wire n_4596;
wire n_5413;
wire n_12459;
wire n_9425;
wire n_7976;
wire n_12648;
wire n_5412;
wire n_17170;
wire n_9620;
wire n_3694;
wire n_2586;
wire n_1398;
wire n_15319;
wire n_14867;
wire n_18753;
wire n_11209;
wire n_2972;
wire n_3225;
wire n_334;
wire n_8199;
wire n_17168;
wire n_3799;
wire n_5201;
wire n_6299;
wire n_9280;
wire n_8016;
wire n_10156;
wire n_8669;
wire n_17605;
wire n_20881;
wire n_11234;
wire n_19776;
wire n_16101;
wire n_12021;
wire n_17804;
wire n_16102;
wire n_7655;
wire n_17209;
wire n_21861;
wire n_17334;
wire n_7737;
wire n_16470;
wire n_18416;
wire n_11000;
wire n_12447;
wire n_4366;
wire n_12667;
wire n_18960;
wire n_278;
wire n_7347;
wire n_9487;
wire n_16552;
wire n_12906;
wire n_7633;
wire n_6177;
wire n_5912;
wire n_611;
wire n_1126;
wire n_10492;
wire n_13023;
wire n_1677;
wire n_19188;
wire n_14753;
wire n_20895;
wire n_1292;
wire n_8888;
wire n_19445;
wire n_12319;
wire n_20761;
wire n_8041;
wire n_9868;
wire n_14442;
wire n_11049;
wire n_10460;
wire n_9292;
wire n_21972;
wire n_12669;
wire n_15492;
wire n_1451;
wire n_1022;
wire n_6917;
wire n_11109;
wire n_5859;
wire n_173;
wire n_859;
wire n_18541;
wire n_10968;
wire n_3571;
wire n_8760;
wire n_19034;
wire n_854;
wire n_2396;
wire n_17558;
wire n_674;
wire n_17076;
wire n_1939;
wire n_2486;
wire n_14276;
wire n_8917;
wire n_6163;
wire n_516;
wire n_10811;
wire n_1152;
wire n_1869;
wire n_13516;
wire n_606;
wire n_3039;
wire n_275;
wire n_2011;
wire n_11737;
wire n_12058;
wire n_11799;
wire n_11788;
wire n_17395;
wire n_18609;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_13143;
wire n_14226;
wire n_21443;
wire n_14106;
wire n_9815;
wire n_8409;
wire n_9110;
wire n_5268;
wire n_6318;
wire n_11453;
wire n_659;
wire n_2639;
wire n_7927;
wire n_6089;
wire n_3325;
wire n_4021;
wire n_11955;
wire n_14596;
wire n_6315;
wire n_938;
wire n_10592;
wire n_7970;
wire n_10476;
wire n_1154;
wire n_8407;
wire n_21065;
wire n_5462;
wire n_13040;
wire n_11488;
wire n_17622;
wire n_12369;
wire n_2761;
wire n_13015;
wire n_17100;
wire n_19937;
wire n_11946;
wire n_9191;
wire n_11918;
wire n_2537;
wire n_2144;
wire n_920;
wire n_18367;
wire n_21356;
wire n_6886;
wire n_13761;
wire n_20333;
wire n_2936;
wire n_18295;
wire n_8783;
wire n_5914;
wire n_14523;
wire n_10695;
wire n_8504;
wire n_8445;
wire n_11950;
wire n_21905;
wire n_4715;
wire n_5039;
wire n_9118;
wire n_13214;
wire n_11410;
wire n_17411;
wire n_20338;
wire n_5542;
wire n_1850;
wire n_163;
wire n_18341;
wire n_17095;
wire n_3669;
wire n_215;
wire n_16840;
wire n_2663;
wire n_21927;
wire n_9123;
wire n_17041;
wire n_5586;
wire n_20777;
wire n_3798;
wire n_6378;
wire n_21711;
wire n_926;
wire n_2249;
wire n_2180;
wire n_14055;
wire n_2632;
wire n_15488;
wire n_777;
wire n_6407;
wire n_21853;
wire n_18872;
wire n_8297;
wire n_6749;
wire n_13921;
wire n_10533;
wire n_13635;
wire n_20786;
wire n_15206;
wire n_4263;
wire n_10455;
wire n_2915;
wire n_2300;
wire n_6217;
wire n_6680;
wire n_12016;
wire n_15837;
wire n_6446;
wire n_8072;
wire n_12017;
wire n_13428;
wire n_11672;
wire n_16016;
wire n_5344;
wire n_15398;
wire n_14914;
wire n_10601;
wire n_12197;
wire n_464;
wire n_19924;
wire n_18667;
wire n_9315;
wire n_9296;
wire n_12660;
wire n_14393;
wire n_14526;
wire n_15278;
wire n_1986;
wire n_4752;
wire n_19071;
wire n_1459;
wire n_14795;
wire n_14691;
wire n_13137;
wire n_11202;
wire n_7656;
wire n_10760;
wire n_7105;
wire n_18264;
wire n_18394;
wire n_2644;
wire n_17313;
wire n_6829;
wire n_9977;
wire n_9887;
wire n_4067;
wire n_7570;
wire n_7262;
wire n_1202;
wire n_8057;
wire n_9333;
wire n_5626;
wire n_16131;
wire n_15947;
wire n_6114;
wire n_1463;
wire n_9590;
wire n_13515;
wire n_3651;
wire n_4333;
wire n_7364;
wire n_12286;
wire n_2706;
wire n_20398;
wire n_11923;
wire n_3676;
wire n_15103;
wire n_17966;
wire n_20267;
wire n_17627;
wire n_10728;
wire n_4815;
wire n_13175;
wire n_4246;
wire n_13759;
wire n_19977;
wire n_18361;
wire n_19915;
wire n_14158;
wire n_10748;
wire n_18409;
wire n_15294;
wire n_6970;
wire n_11842;
wire n_20658;
wire n_2674;
wire n_7778;
wire n_4357;
wire n_3371;
wire n_15563;
wire n_12532;
wire n_4472;
wire n_647;
wire n_7320;
wire n_6255;
wire n_7343;
wire n_18980;
wire n_11473;
wire n_13735;
wire n_7875;
wire n_16065;
wire n_21160;
wire n_16113;
wire n_13258;
wire n_21291;
wire n_15891;
wire n_4151;
wire n_13617;
wire n_17207;
wire n_3528;
wire n_19495;
wire n_12138;
wire n_21285;
wire n_15175;
wire n_13013;
wire n_2322;
wire n_9219;
wire n_13625;
wire n_6427;
wire n_13054;
wire n_7753;
wire n_11924;
wire n_15410;
wire n_4344;
wire n_1368;
wire n_2762;
wire n_8392;
wire n_21610;
wire n_12967;
wire n_15383;
wire n_17702;
wire n_1162;
wire n_16080;
wire n_6360;
wire n_13026;
wire n_9553;
wire n_3602;
wire n_2967;
wire n_887;
wire n_10616;
wire n_19164;
wire n_5477;
wire n_20853;
wire n_12695;
wire n_3923;
wire n_11526;
wire n_11742;
wire n_20086;
wire n_18363;
wire n_18067;
wire n_18854;
wire n_2801;
wire n_17535;
wire n_20385;
wire n_4011;
wire n_15088;
wire n_2825;
wire n_15384;
wire n_17841;
wire n_12105;
wire n_9793;
wire n_6691;
wire n_3748;
wire n_17571;
wire n_20525;
wire n_20958;
wire n_187;
wire n_12360;
wire n_3370;
wire n_5053;
wire n_7912;
wire n_1259;
wire n_4553;
wire n_14981;
wire n_18338;
wire n_15936;
wire n_18404;
wire n_19886;
wire n_2491;
wire n_20059;
wire n_10331;
wire n_6773;
wire n_17840;
wire n_1222;
wire n_21948;
wire n_21901;
wire n_19730;
wire n_8463;
wire n_14120;
wire n_7041;
wire n_7802;
wire n_15489;
wire n_18496;
wire n_13366;
wire n_10074;
wire n_1191;
wire n_16885;
wire n_2992;
wire n_14529;
wire n_18612;
wire n_4920;
wire n_12828;
wire n_6776;
wire n_18038;
wire n_13078;
wire n_5426;
wire n_19905;
wire n_17730;
wire n_20444;
wire n_13387;
wire n_2631;
wire n_13226;
wire n_11037;
wire n_1529;
wire n_10381;
wire n_15237;
wire n_8517;
wire n_5778;
wire n_6396;
wire n_3355;
wire n_2007;
wire n_10569;
wire n_12326;
wire n_15830;
wire n_5531;
wire n_16867;
wire n_739;
wire n_1406;
wire n_1839;
wire n_17404;
wire n_5248;
wire n_11042;
wire n_12141;
wire n_12622;
wire n_11226;
wire n_16126;
wire n_999;
wire n_9358;
wire n_20602;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_19769;
wire n_10127;
wire n_21667;
wire n_3988;
wire n_563;
wire n_6161;
wire n_21432;
wire n_18620;
wire n_19871;
wire n_7987;
wire n_10328;
wire n_1871;
wire n_3630;
wire n_12343;
wire n_5719;
wire n_4771;
wire n_17598;
wire n_7037;
wire n_14900;
wire n_14966;
wire n_19633;
wire n_1781;
wire n_15646;
wire n_3075;
wire n_18814;
wire n_16495;
wire n_3701;
wire n_15209;
wire n_15818;
wire n_13999;
wire n_1773;
wire n_6334;
wire n_2666;
wire n_8984;
wire n_21842;
wire n_14502;
wire n_4708;
wire n_2314;
wire n_9268;
wire n_8764;
wire n_6794;
wire n_16865;
wire n_2420;
wire n_3343;
wire n_10245;
wire n_19425;
wire n_12466;
wire n_18797;
wire n_5489;
wire n_19074;
wire n_3767;
wire n_442;
wire n_12560;
wire n_2873;
wire n_2540;
wire n_4589;
wire n_15909;
wire n_5057;
wire n_10280;
wire n_16066;
wire n_19635;
wire n_19751;
wire n_6705;
wire n_14559;
wire n_9636;
wire n_19790;
wire n_3221;
wire n_5907;
wire n_11120;
wire n_2168;
wire n_11391;
wire n_6044;
wire n_185;
wire n_5286;
wire n_3502;
wire n_8853;
wire n_11371;
wire n_6495;
wire n_18628;
wire n_6902;
wire n_11591;
wire n_9560;
wire n_8711;
wire n_10976;
wire n_8229;
wire n_17776;
wire n_15127;
wire n_3607;
wire n_14079;
wire n_7548;
wire n_15112;
wire n_20246;
wire n_11460;
wire n_8567;
wire n_17056;
wire n_4510;
wire n_2571;
wire n_9235;
wire n_2124;
wire n_5715;
wire n_9085;
wire n_8085;
wire n_11891;
wire n_6528;
wire n_16546;
wire n_7604;
wire n_14499;
wire n_3827;
wire n_20800;
wire n_10845;
wire n_4447;
wire n_15942;
wire n_6774;
wire n_20622;
wire n_5887;
wire n_4651;
wire n_20098;
wire n_6741;
wire n_7424;
wire n_11557;
wire n_573;
wire n_18305;
wire n_20555;
wire n_13228;
wire n_19370;
wire n_13244;
wire n_12134;
wire n_582;
wire n_16317;
wire n_4433;
wire n_18922;
wire n_11163;
wire n_2879;
wire n_19384;
wire n_16446;
wire n_19513;
wire n_6700;
wire n_8098;
wire n_13880;
wire n_3399;
wire n_14418;
wire n_13011;
wire n_20179;
wire n_19887;
wire n_10503;
wire n_20896;
wire n_14880;
wire n_11732;
wire n_6012;
wire n_16630;
wire n_13222;
wire n_20482;
wire n_21017;
wire n_3675;
wire n_18959;
wire n_14136;
wire n_19954;
wire n_15961;
wire n_1140;
wire n_3387;
wire n_12550;
wire n_15772;
wire n_19753;
wire n_21924;
wire n_18239;
wire n_20260;
wire n_18114;
wire n_11508;
wire n_12965;
wire n_5828;
wire n_11634;
wire n_4993;
wire n_13402;
wire n_6337;
wire n_18755;
wire n_8970;
wire n_1885;
wire n_10119;
wire n_20978;
wire n_20905;
wire n_6770;
wire n_13218;
wire n_5238;
wire n_13239;
wire n_8856;
wire n_16926;
wire n_4595;
wire n_21991;
wire n_11503;
wire n_16140;
wire n_7799;
wire n_16022;
wire n_21778;
wire n_2288;
wire n_6314;
wire n_17084;
wire n_13983;
wire n_346;
wire n_21246;
wire n_3592;
wire n_5694;
wire n_8774;
wire n_7274;
wire n_17808;
wire n_5326;
wire n_20879;
wire n_14199;
wire n_13949;
wire n_8779;
wire n_879;
wire n_3394;
wire n_17021;
wire n_13090;
wire n_19216;
wire n_18602;
wire n_405;
wire n_12558;
wire n_19204;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_11288;
wire n_18354;
wire n_5528;
wire n_11027;
wire n_16448;
wire n_7785;
wire n_5422;
wire n_18434;
wire n_12591;
wire n_20770;
wire n_16518;
wire n_3059;
wire n_10581;
wire n_3465;
wire n_9576;
wire n_14832;
wire n_10097;
wire n_952;
wire n_1229;
wire n_18773;
wire n_4799;
wire n_9651;
wire n_6257;
wire n_14240;
wire n_12690;
wire n_3449;
wire n_18894;
wire n_13076;
wire n_17592;
wire n_2989;
wire n_10813;
wire n_2789;
wire n_21780;
wire n_2216;
wire n_531;
wire n_19878;
wire n_12414;
wire n_1897;
wire n_764;
wire n_16743;
wire n_2933;
wire n_19965;
wire n_17175;
wire n_5354;
wire n_6274;
wire n_7372;
wire n_10943;
wire n_7685;
wire n_8750;
wire n_14649;
wire n_4845;
wire n_9364;
wire n_16334;
wire n_9512;
wire n_17274;
wire n_3893;
wire n_14661;
wire n_8593;
wire n_14047;
wire n_18258;
wire n_17548;
wire n_2465;
wire n_21814;
wire n_7730;
wire n_315;
wire n_13165;
wire n_9314;
wire n_9459;
wire n_3334;
wire n_9549;
wire n_1139;
wire n_18926;
wire n_13670;
wire n_15245;
wire n_15102;
wire n_10210;
wire n_5370;
wire n_11944;
wire n_7706;
wire n_5594;
wire n_14301;
wire n_9865;
wire n_18191;
wire n_6471;
wire n_16816;
wire n_11511;
wire n_12981;
wire n_10263;
wire n_21521;
wire n_7512;
wire n_1644;
wire n_5550;
wire n_20043;
wire n_15405;
wire n_9656;
wire n_15442;
wire n_3537;
wire n_3080;
wire n_13004;
wire n_3362;
wire n_5559;
wire n_12694;
wire n_19080;
wire n_6488;
wire n_1048;
wire n_13864;
wire n_9629;
wire n_21397;
wire n_16590;
wire n_2556;
wire n_16347;
wire n_6457;
wire n_20101;
wire n_4470;
wire n_18726;
wire n_19873;
wire n_13874;
wire n_21381;
wire n_820;
wire n_3616;
wire n_10494;
wire n_4058;
wire n_3664;
wire n_16772;
wire n_10743;
wire n_21951;
wire n_8583;
wire n_20772;
wire n_4034;
wire n_15524;
wire n_15989;
wire n_18965;
wire n_492;
wire n_3327;
wire n_20090;
wire n_21756;
wire n_13274;
wire n_13827;
wire n_10050;
wire n_341;
wire n_7311;
wire n_19458;
wire n_5989;
wire n_8964;
wire n_543;
wire n_18080;
wire n_11388;
wire n_13786;
wire n_8539;
wire n_8745;
wire n_6456;
wire n_1214;
wire n_15568;
wire n_9319;
wire n_8554;
wire n_11748;
wire n_5227;
wire n_20990;
wire n_13463;
wire n_21591;
wire n_14351;
wire n_9442;
wire n_18095;
wire n_20701;
wire n_14385;
wire n_7198;
wire n_8802;
wire n_9587;
wire n_19864;
wire n_618;
wire n_8955;
wire n_12510;
wire n_17608;
wire n_1373;
wire n_7249;
wire n_14186;
wire n_4539;
wire n_18829;
wire n_17082;
wire n_18073;
wire n_14853;
wire n_16400;
wire n_17563;
wire n_13193;
wire n_13739;
wire n_12628;
wire n_7142;
wire n_3230;
wire n_3342;
wire n_6054;
wire n_7089;
wire n_4682;
wire n_12445;
wire n_16920;
wire n_17463;
wire n_3729;
wire n_14023;
wire n_4978;
wire n_21831;
wire n_12281;
wire n_12355;
wire n_5458;
wire n_8778;
wire n_10415;
wire n_17907;
wire n_6523;
wire n_13127;
wire n_14581;
wire n_16282;
wire n_3957;
wire n_12004;
wire n_11893;
wire n_20652;
wire n_8194;
wire n_14125;
wire n_2600;
wire n_20775;
wire n_19999;
wire n_13414;
wire n_7181;
wire n_5384;
wire n_8582;
wire n_10378;
wire n_17063;
wire n_216;
wire n_6056;
wire n_17438;
wire n_21023;
wire n_13425;
wire n_3829;
wire n_8951;
wire n_7818;
wire n_5125;
wire n_12024;
wire n_2207;
wire n_2619;
wire n_13182;
wire n_18158;
wire n_1110;
wire n_16952;
wire n_14787;
wire n_16237;
wire n_19476;
wire n_21084;
wire n_6369;
wire n_5056;
wire n_17201;
wire n_14883;
wire n_3393;
wire n_22002;
wire n_5360;
wire n_5269;
wire n_249;
wire n_5866;
wire n_8568;
wire n_12857;
wire n_20406;
wire n_9916;
wire n_13682;
wire n_16702;
wire n_693;
wire n_8716;
wire n_1389;
wire n_7601;
wire n_1256;
wire n_11135;
wire n_1465;
wire n_6026;
wire n_15177;
wire n_21193;
wire n_19791;
wire n_14335;
wire n_10075;
wire n_3727;
wire n_10068;
wire n_11596;
wire n_16877;
wire n_18945;
wire n_12555;
wire n_21315;
wire n_19338;
wire n_6679;
wire n_13296;
wire n_18324;
wire n_1371;
wire n_4956;
wire n_2206;
wire n_12839;
wire n_10495;
wire n_20549;
wire n_6259;
wire n_16551;
wire n_12983;
wire n_16361;
wire n_12945;
wire n_3450;
wire n_20657;
wire n_4729;
wire n_17567;
wire n_19365;
wire n_12451;
wire n_12376;
wire n_9022;
wire n_1453;
wire n_6630;
wire n_15463;
wire n_1183;
wire n_16817;
wire n_16133;
wire n_18108;
wire n_13256;
wire n_3432;
wire n_1514;
wire n_9344;
wire n_557;
wire n_15979;
wire n_15618;
wire n_10603;
wire n_17156;
wire n_527;
wire n_1168;
wire n_9764;
wire n_17164;
wire n_11294;
wire n_13024;
wire n_8273;
wire n_19148;
wire n_11021;
wire n_177;
wire n_9242;
wire n_9498;
wire n_8442;
wire n_7106;
wire n_16582;
wire n_1356;
wire n_6057;
wire n_7529;
wire n_2634;
wire n_910;
wire n_13740;
wire n_16576;
wire n_3972;
wire n_17314;
wire n_13064;
wire n_11951;
wire n_12219;
wire n_17814;
wire n_20830;
wire n_18631;
wire n_1533;
wire n_18320;
wire n_20062;
wire n_5547;
wire n_19130;
wire n_12758;
wire n_13302;
wire n_1720;
wire n_10972;
wire n_6291;
wire n_159;
wire n_17865;
wire n_14167;
wire n_20316;
wire n_18221;
wire n_9510;
wire n_1480;
wire n_9413;
wire n_7648;
wire n_9888;
wire n_8393;
wire n_18347;
wire n_21715;
wire n_11484;
wire n_8821;
wire n_11760;
wire n_10881;
wire n_8160;
wire n_9014;
wire n_10204;
wire n_11909;
wire n_2965;
wire n_5022;
wire n_18736;
wire n_14783;
wire n_3046;
wire n_18811;
wire n_19326;
wire n_10717;
wire n_13931;
wire n_13541;
wire n_3211;
wire n_14710;
wire n_20584;
wire n_5703;
wire n_19754;
wire n_8240;
wire n_12450;
wire n_21800;
wire n_20244;
wire n_20178;
wire n_14643;
wire n_8579;
wire n_12444;
wire n_8258;
wire n_9854;
wire n_6540;
wire n_1822;
wire n_16375;
wire n_13936;
wire n_18738;
wire n_17591;
wire n_4126;
wire n_5087;
wire n_18289;
wire n_3802;
wire n_4506;
wire n_11792;
wire n_17868;
wire n_17519;
wire n_4896;
wire n_7063;
wire n_2107;
wire n_4943;
wire n_2187;
wire n_8012;
wire n_11445;
wire n_718;
wire n_18405;
wire n_14464;
wire n_19578;
wire n_12228;
wire n_11832;
wire n_15953;
wire n_21679;
wire n_19875;
wire n_6487;
wire n_9146;
wire n_18140;
wire n_17309;
wire n_10283;
wire n_13944;
wire n_5195;
wire n_15926;
wire n_1715;
wire n_12742;
wire n_4393;
wire n_10618;
wire n_3720;
wire n_8576;
wire n_21409;
wire n_4535;
wire n_733;
wire n_18764;
wire n_21094;
wire n_6656;
wire n_21996;
wire n_792;
wire n_18342;
wire n_8148;
wire n_19833;
wire n_7953;
wire n_8343;
wire n_2104;
wire n_15850;
wire n_16809;
wire n_5164;
wire n_15173;
wire n_6485;
wire n_14882;
wire n_5498;
wire n_20543;
wire n_5183;
wire n_21073;
wire n_20784;
wire n_17375;
wire n_6120;
wire n_16878;
wire n_19979;
wire n_3412;
wire n_1995;
wire n_2411;
wire n_3761;
wire n_7689;
wire n_2986;
wire n_13792;
wire n_7824;
wire n_20869;
wire n_15832;
wire n_8726;
wire n_7796;
wire n_20493;
wire n_2172;
wire n_9450;
wire n_13272;
wire n_18025;
wire n_16797;
wire n_14725;
wire n_8796;
wire n_18536;
wire n_11638;
wire n_4100;
wire n_15246;
wire n_961;
wire n_2250;
wire n_7084;
wire n_9617;
wire n_8883;
wire n_169;
wire n_16634;
wire n_8251;
wire n_5990;
wire n_15464;
wire n_7253;
wire n_5663;
wire n_20156;
wire n_994;
wire n_20997;
wire n_5973;
wire n_15184;
wire n_12849;
wire n_19725;
wire n_15822;
wire n_19710;
wire n_18480;
wire n_5304;
wire n_13863;
wire n_5130;
wire n_16985;
wire n_12329;
wire n_12032;
wire n_12159;
wire n_9490;
wire n_6809;
wire n_11213;
wire n_12987;
wire n_12504;
wire n_8165;
wire n_15163;
wire n_18810;
wire n_16645;
wire n_9002;
wire n_11100;
wire n_17752;
wire n_13695;
wire n_18791;
wire n_14030;
wire n_8330;
wire n_5757;
wire n_20974;
wire n_17389;
wire n_20229;
wire n_7918;
wire n_11440;
wire n_21220;
wire n_8467;
wire n_13216;
wire n_18986;
wire n_21731;
wire n_16692;
wire n_12482;
wire n_4116;
wire n_21877;
wire n_17994;
wire n_16105;
wire n_16443;
wire n_18406;
wire n_9867;
wire n_1086;
wire n_1469;
wire n_15501;
wire n_2397;
wire n_15580;
wire n_16249;
wire n_17514;
wire n_384;
wire n_2208;
wire n_20689;
wire n_3063;
wire n_15011;
wire n_15152;
wire n_15244;
wire n_15122;
wire n_11189;
wire n_3794;
wire n_14779;
wire n_4505;
wire n_16269;
wire n_10542;
wire n_9611;
wire n_15203;
wire n_15217;
wire n_2591;
wire n_852;
wire n_8186;
wire n_1864;
wire n_6067;
wire n_9774;
wire n_5070;
wire n_13793;
wire n_420;
wire n_1337;
wire n_699;
wire n_8738;
wire n_16084;
wire n_18979;
wire n_1627;
wire n_13186;
wire n_19976;
wire n_10645;
wire n_18107;
wire n_273;
wire n_17748;
wire n_5296;
wire n_17251;
wire n_15147;
wire n_18624;
wire n_11195;
wire n_21652;
wire n_17331;
wire n_12254;
wire n_13580;
wire n_14178;
wire n_16462;
wire n_4914;
wire n_10737;
wire n_5834;
wire n_1076;
wire n_5874;
wire n_16229;
wire n_7977;
wire n_14582;
wire n_16643;
wire n_18310;
wire n_730;
wire n_7508;
wire n_13831;
wire n_11345;
wire n_5956;
wire n_14670;
wire n_18844;
wire n_4345;
wire n_14349;
wire n_10243;
wire n_3307;
wire n_7000;
wire n_1694;
wire n_15627;
wire n_18599;
wire n_10038;
wire n_17482;
wire n_10410;
wire n_16364;
wire n_2366;
wire n_15070;
wire n_3997;
wire n_1604;
wire n_16355;
wire n_5465;
wire n_1764;
wire n_16605;
wire n_3582;
wire n_20801;
wire n_7517;
wire n_17905;
wire n_5853;
wire n_15504;
wire n_2826;
wire n_15994;
wire n_14497;
wire n_17009;
wire n_17677;
wire n_12359;
wire n_11577;
wire n_5467;
wire n_21455;
wire n_4928;
wire n_1507;
wire n_4378;
wire n_16779;
wire n_4216;
wire n_12688;
wire n_19593;
wire n_20285;
wire n_6942;
wire n_2019;
wire n_1340;
wire n_9577;
wire n_2166;
wire n_3594;
wire n_14338;
wire n_2026;
wire n_9513;
wire n_1234;
wire n_21632;
wire n_1990;
wire n_11759;
wire n_2614;
wire n_10710;
wire n_17044;
wire n_7997;
wire n_20115;
wire n_9130;
wire n_2242;
wire n_2894;
wire n_11829;
wire n_17304;
wire n_7047;
wire n_8144;
wire n_14077;
wire n_18976;
wire n_2524;
wire n_20238;
wire n_13055;
wire n_11308;
wire n_13115;
wire n_6643;
wire n_18022;
wire n_6122;
wire n_2417;
wire n_2756;
wire n_16520;
wire n_7981;
wire n_15472;
wire n_12407;
wire n_9325;
wire n_7164;
wire n_17478;
wire n_15306;
wire n_2327;
wire n_19363;
wire n_21508;
wire n_3619;
wire n_5978;
wire n_20778;
wire n_5512;
wire n_14764;
wire n_14635;
wire n_20099;
wire n_17997;
wire n_9044;
wire n_17360;
wire n_7206;
wire n_19047;
wire n_15682;
wire n_9408;
wire n_4508;
wire n_8363;
wire n_12975;
wire n_11802;
wire n_10885;
wire n_2843;
wire n_2487;
wire n_1695;
wire n_19103;
wire n_8551;
wire n_14264;
wire n_17586;
wire n_18900;
wire n_18776;
wire n_13386;
wire n_21351;
wire n_12071;
wire n_12738;
wire n_20318;
wire n_16752;
wire n_4128;
wire n_8976;
wire n_4145;
wire n_20732;
wire n_15940;
wire n_9846;
wire n_7024;
wire n_19288;
wire n_16301;
wire n_9204;
wire n_13493;
wire n_16208;
wire n_9610;
wire n_877;
wire n_21669;
wire n_1696;
wire n_13220;
wire n_4988;
wire n_1285;
wire n_12028;
wire n_12357;
wire n_21106;
wire n_19292;
wire n_4615;
wire n_1728;
wire n_6090;
wire n_12515;
wire n_7010;
wire n_5480;
wire n_13158;
wire n_21723;
wire n_7315;
wire n_7004;
wire n_2770;
wire n_171;
wire n_3188;
wire n_20612;
wire n_8574;
wire n_3403;
wire n_16846;
wire n_20921;
wire n_3624;
wire n_8864;
wire n_21642;
wire n_20200;
wire n_3461;
wire n_19564;
wire n_7641;
wire n_21771;
wire n_3796;
wire n_15567;
wire n_5154;
wire n_3283;
wire n_19996;
wire n_11800;
wire n_2323;
wire n_16313;
wire n_19971;
wire n_2597;
wire n_18993;
wire n_15377;
wire n_14537;
wire n_2052;
wire n_16655;
wire n_9738;
wire n_19120;
wire n_1314;
wire n_18752;
wire n_317;
wire n_13771;
wire n_21538;
wire n_6408;
wire n_3214;
wire n_17245;
wire n_1517;
wire n_14800;
wire n_8706;
wire n_3806;
wire n_4691;
wire n_13000;
wire n_11594;
wire n_6698;
wire n_4678;
wire n_2587;
wire n_8104;
wire n_5848;
wire n_16689;
wire n_3490;
wire n_600;
wire n_15753;
wire n_10360;
wire n_1948;
wire n_18774;
wire n_9420;
wire n_9557;
wire n_12604;
wire n_19918;
wire n_10781;
wire n_11507;
wire n_7562;
wire n_10193;
wire n_9388;
wire n_4468;
wire n_16192;
wire n_21384;
wire n_9772;
wire n_3702;
wire n_1040;
wire n_8147;
wire n_6586;
wire n_11111;
wire n_5008;
wire n_5398;
wire n_19048;
wire n_2276;
wire n_14170;
wire n_10175;
wire n_2089;
wire n_9311;
wire n_17297;
wire n_18546;
wire n_553;
wire n_20749;
wire n_1880;
wire n_16324;
wire n_13309;
wire n_18683;
wire n_2238;
wire n_1151;
wire n_1706;
wire n_17010;
wire n_20617;
wire n_20104;
wire n_18035;
wire n_13542;
wire n_10683;
wire n_14109;
wire n_2859;
wire n_1075;
wire n_7086;
wire n_7349;
wire n_8317;
wire n_13706;
wire n_7647;
wire n_12224;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_10252;
wire n_9780;
wire n_4421;
wire n_10438;
wire n_19371;
wire n_18071;
wire n_16487;
wire n_19788;
wire n_15481;
wire n_15106;
wire n_11659;
wire n_1377;
wire n_5184;
wire n_7956;
wire n_15823;
wire n_12824;
wire n_21859;
wire n_9489;
wire n_8604;
wire n_15932;
wire n_11365;
wire n_13755;
wire n_11836;
wire n_7683;
wire n_19902;
wire n_1002;
wire n_19386;
wire n_3487;
wire n_11003;
wire n_838;
wire n_3983;
wire n_1224;
wire n_22004;
wire n_1926;
wire n_19342;
wire n_8416;
wire n_17273;
wire n_13219;
wire n_4969;
wire n_13547;
wire n_7575;
wire n_2776;
wire n_8879;
wire n_10664;
wire n_19571;
wire n_9115;
wire n_9367;
wire n_4531;
wire n_6043;
wire n_16780;
wire n_13747;
wire n_12812;
wire n_6271;
wire n_7171;
wire n_13223;
wire n_5315;
wire n_345;
wire n_4130;
wire n_21824;
wire n_15290;
wire n_2175;
wire n_5055;
wire n_14973;
wire n_16025;
wire n_20214;
wire n_12777;
wire n_20659;
wire n_14886;
wire n_16883;
wire n_3975;
wire n_15503;
wire n_21866;
wire n_6021;
wire n_4983;
wire n_9213;
wire n_7814;
wire n_21249;
wire n_21471;
wire n_10778;
wire n_4916;
wire n_11121;
wire n_3649;
wire n_7589;
wire n_5862;
wire n_19951;
wire n_21940;
wire n_19960;
wire n_1027;
wire n_6782;
wire n_5516;
wire n_4051;
wire n_9554;
wire n_15281;
wire n_17261;
wire n_12412;
wire n_1276;
wire n_20526;
wire n_18956;
wire n_10935;
wire n_19428;
wire n_6126;
wire n_19185;
wire n_12612;
wire n_8795;
wire n_352;
wire n_1038;
wire n_520;
wire n_10401;
wire n_6598;
wire n_4647;
wire n_870;
wire n_16183;
wire n_12180;
wire n_6900;
wire n_14016;
wire n_13295;
wire n_19208;
wire n_965;
wire n_3790;
wire n_7264;
wire n_3491;
wire n_12608;
wire n_7457;
wire n_16556;
wire n_4649;
wire n_7617;
wire n_16940;
wire n_19876;
wire n_9197;
wire n_20055;
wire n_21338;
wire n_21170;
wire n_5615;
wire n_2226;
wire n_12057;
wire n_2891;
wire n_14098;
wire n_19750;
wire n_15913;
wire n_14143;
wire n_5479;
wire n_19168;
wire n_10964;
wire n_13234;
wire n_16020;
wire n_13896;
wire n_20933;
wire n_6013;
wire n_9564;
wire n_10864;
wire n_2297;
wire n_9739;
wire n_15687;
wire n_1759;
wire n_17642;
wire n_2227;
wire n_3346;
wire n_21110;
wire n_452;
wire n_1746;
wire n_17938;
wire n_21257;
wire n_9812;
wire n_1464;
wire n_14905;
wire n_649;
wire n_17978;
wire n_10553;
wire n_19478;
wire n_12393;
wire n_16914;
wire n_7076;
wire n_21369;
wire n_8780;
wire n_19759;
wire n_9928;
wire n_17410;
wire n_19772;
wire n_3038;
wire n_14238;
wire n_3068;
wire n_5943;
wire n_14641;
wire n_17491;
wire n_1680;
wire n_14713;
wire n_18019;
wire n_13167;
wire n_15185;
wire n_7848;
wire n_6727;
wire n_8218;
wire n_9267;
wire n_18775;
wire n_4391;
wire n_19805;
wire n_11865;
wire n_4157;
wire n_15605;
wire n_8368;
wire n_12163;
wire n_1468;
wire n_18963;
wire n_6097;
wire n_14116;
wire n_12516;
wire n_20247;
wire n_18045;
wire n_1994;
wire n_6677;
wire n_1195;
wire n_20906;
wire n_14740;
wire n_6624;
wire n_7121;
wire n_18215;
wire n_21551;
wire n_17546;
wire n_15285;
wire n_14830;
wire n_4156;
wire n_19687;
wire n_14975;
wire n_12198;
wire n_21491;
wire n_11201;
wire n_15404;
wire n_7781;
wire n_524;
wire n_14677;
wire n_5714;
wire n_5806;
wire n_13675;
wire n_741;
wire n_10653;
wire n_20142;
wire n_4898;
wire n_16741;
wire n_1163;
wire n_8063;
wire n_21010;
wire n_15229;
wire n_6185;
wire n_1207;
wire n_5010;
wire n_13097;
wire n_21151;
wire n_7762;
wire n_8731;
wire n_15744;
wire n_2846;
wire n_17718;
wire n_2925;
wire n_21191;
wire n_3918;
wire n_16075;
wire n_14955;
wire n_12802;
wire n_9011;
wire n_20243;
wire n_4528;
wire n_3932;
wire n_16697;
wire n_12570;
wire n_4673;
wire n_940;
wire n_7552;
wire n_8059;
wire n_19988;
wire n_3516;
wire n_20959;
wire n_2516;
wire n_3797;
wire n_2947;
wire n_16661;
wire n_18470;
wire n_14589;
wire n_1269;
wire n_18082;
wire n_2473;
wire n_19092;
wire n_11816;
wire n_7746;
wire n_14068;
wire n_11062;
wire n_18131;
wire n_6873;
wire n_14610;
wire n_8032;
wire n_12710;
wire n_10016;
wire n_1732;
wire n_10070;
wire n_19171;
wire n_17246;
wire n_4125;
wire n_374;
wire n_10190;
wire n_20962;
wire n_12128;
wire n_6594;
wire n_962;
wire n_10812;
wire n_20530;
wire n_9460;
wire n_17184;
wire n_9638;
wire n_19459;
wire n_19343;
wire n_17600;
wire n_6387;
wire n_1336;
wire n_10134;
wire n_11379;
wire n_13700;
wire n_20518;
wire n_18632;
wire n_9740;
wire n_17469;
wire n_12147;
wire n_9190;
wire n_19159;
wire n_19919;
wire n_4610;
wire n_12909;
wire n_18699;
wire n_4489;
wire n_3730;
wire n_18447;
wire n_16805;
wire n_6976;
wire n_4967;
wire n_15547;
wire n_5657;
wire n_16685;
wire n_6889;
wire n_17363;
wire n_3945;
wire n_18816;
wire n_9891;
wire n_6295;
wire n_9804;
wire n_16392;
wire n_18492;
wire n_8087;
wire n_12468;
wire n_18130;
wire n_4534;
wire n_15242;
wire n_6241;
wire n_14035;
wire n_8019;
wire n_15327;
wire n_20842;
wire n_13307;
wire n_14921;
wire n_11335;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_20833;
wire n_13509;
wire n_16349;
wire n_19018;
wire n_20664;
wire n_2231;
wire n_2017;
wire n_14949;
wire n_6994;
wire n_10987;
wire n_322;
wire n_15599;
wire n_13238;
wire n_21070;
wire n_14813;
wire n_6790;
wire n_12860;
wire n_20220;
wire n_15801;
wire n_10666;
wire n_19533;
wire n_20009;
wire n_6273;
wire n_14482;
wire n_19784;
wire n_15433;
wire n_16581;
wire n_10189;
wire n_9879;
wire n_17114;
wire n_8221;
wire n_1913;
wire n_8468;
wire n_18137;
wire n_3679;
wire n_13211;
wire n_15570;
wire n_3422;
wire n_7115;
wire n_18102;
wire n_13391;
wire n_5584;
wire n_14102;
wire n_3429;
wire n_21513;
wire n_3849;
wire n_3946;
wire n_5965;
wire n_19275;
wire n_13475;
wire n_10434;
wire n_9441;
wire n_11913;
wire n_15718;
wire n_19044;
wire n_5641;
wire n_6218;
wire n_8863;
wire n_19715;
wire n_8106;
wire n_21425;
wire n_20795;
wire n_2727;
wire n_10690;
wire n_20437;
wire n_14212;
wire n_560;
wire n_15639;
wire n_20949;
wire n_20358;
wire n_18188;
wire n_16857;
wire n_9200;
wire n_21223;
wire n_3683;
wire n_13787;
wire n_16187;
wire n_5980;
wire n_824;
wire n_18070;
wire n_18257;
wire n_14445;
wire n_3590;
wire n_12846;
wire n_8287;
wire n_15604;
wire n_13550;
wire n_7989;
wire n_3424;
wire n_12908;
wire n_1037;
wire n_21035;
wire n_15997;
wire n_12747;
wire n_21960;
wire n_12426;
wire n_2419;
wire n_5146;
wire n_589;
wire n_19926;
wire n_15621;
wire n_16600;
wire n_13067;
wire n_7192;
wire n_11324;
wire n_20890;
wire n_15803;
wire n_238;
wire n_11566;
wire n_7580;
wire n_9880;
wire n_10072;
wire n_11869;
wire n_3462;
wire n_14326;
wire n_222;
wire n_20715;
wire n_8559;
wire n_15938;
wire n_10838;
wire n_14075;
wire n_634;
wire n_6967;
wire n_6433;
wire n_12178;
wire n_9128;
wire n_20887;
wire n_1519;
wire n_950;
wire n_19628;
wire n_5461;
wire n_13192;
wire n_16333;
wire n_1811;
wire n_7632;
wire n_16608;
wire n_4575;
wire n_12554;
wire n_8771;
wire n_380;
wire n_9528;
wire n_18028;
wire n_12912;
wire n_20946;
wire n_19319;
wire n_11529;
wire n_9507;
wire n_22008;
wire n_17301;
wire n_16389;
wire n_19688;
wire n_13557;
wire n_9533;
wire n_5362;
wire n_15924;
wire n_16901;
wire n_16023;
wire n_15941;
wire n_19696;
wire n_20160;
wire n_14379;
wire n_14991;
wire n_721;
wire n_12171;
wire n_1157;
wire n_12815;
wire n_12472;
wire n_19723;
wire n_16815;
wire n_8090;
wire n_10504;
wire n_15715;
wire n_2265;
wire n_4104;
wire n_3554;
wire n_4377;
wire n_17024;
wire n_5266;
wire n_13418;
wire n_873;
wire n_16434;
wire n_17540;
wire n_2334;
wire n_18163;
wire n_690;
wire n_8260;
wire n_15261;
wire n_583;
wire n_6811;
wire n_3051;
wire n_6209;
wire n_13799;
wire n_15369;
wire n_17755;
wire n_3632;
wire n_14685;
wire n_18749;
wire n_20980;
wire n_11076;
wire n_1288;
wire n_212;
wire n_14877;
wire n_2415;
wire n_5551;
wire n_3715;
wire n_7803;
wire n_7747;
wire n_15648;
wire n_6073;
wire n_19352;
wire n_8401;
wire n_3040;
wire n_20593;
wire n_1938;
wire n_10199;
wire n_13020;
wire n_19703;
wire n_14310;
wire n_5475;
wire n_3737;
wire n_14608;
wire n_1185;
wire n_8510;
wire n_1967;
wire n_576;
wire n_13163;
wire n_4856;
wire n_7726;
wire n_11623;
wire n_12825;
wire n_5921;
wire n_8024;
wire n_21907;
wire n_13119;
wire n_6477;
wire n_3734;
wire n_14469;
wire n_19222;
wire n_4778;
wire n_21079;
wire n_6159;
wire n_19589;
wire n_9647;
wire n_6283;
wire n_21661;
wire n_14237;
wire n_16617;
wire n_16884;
wire n_11698;
wire n_856;
wire n_17365;
wire n_10485;
wire n_16879;
wire n_6943;
wire n_9329;
wire n_4761;
wire n_10652;
wire n_6173;
wire n_4095;
wire n_8543;
wire n_14803;
wire n_18867;
wire n_13994;
wire n_5371;
wire n_12334;
wire n_2291;
wire n_20872;
wire n_15044;
wire n_11196;
wire n_12847;
wire n_16037;
wire n_7770;
wire n_18000;
wire n_1865;
wire n_16939;
wire n_19081;
wire n_7664;
wire n_19078;
wire n_13969;
wire n_15005;
wire n_225;
wire n_20226;
wire n_21045;
wire n_13209;
wire n_2751;
wire n_11609;
wire n_16853;
wire n_13712;
wire n_14864;
wire n_4406;
wire n_2758;
wire n_13263;
wire n_18839;
wire n_2618;
wire n_7428;
wire n_763;
wire n_17797;
wire n_9766;
wire n_16213;
wire n_2840;
wire n_2822;
wire n_287;
wire n_20451;
wire n_12409;
wire n_11307;
wire n_19854;
wire n_4117;
wire n_15477;
wire n_10703;
wire n_16048;
wire n_19583;
wire n_11973;
wire n_21289;
wire n_4487;
wire n_19819;
wire n_5001;
wire n_9622;
wire n_19853;
wire n_16387;
wire n_21553;
wire n_11252;
wire n_20785;
wire n_4817;
wire n_19033;
wire n_3380;
wire n_21794;
wire n_13865;
wire n_12454;
wire n_19669;
wire n_10103;
wire n_19490;
wire n_16793;
wire n_2068;
wire n_21595;
wire n_2641;
wire n_20273;
wire n_20682;
wire n_10995;
wire n_17443;
wire n_20286;
wire n_9794;
wire n_11858;
wire n_4728;
wire n_13963;
wire n_7117;
wire n_14845;
wire n_20671;
wire n_789;
wire n_9354;
wire n_4933;
wire n_21472;
wire n_13448;
wire n_15931;
wire n_21097;
wire n_1105;
wire n_17226;
wire n_11478;
wire n_16228;
wire n_12955;
wire n_21772;
wire n_18266;
wire n_3872;
wire n_10856;
wire n_13626;
wire n_4336;
wire n_17792;
wire n_20802;
wire n_2496;
wire n_20261;
wire n_16132;
wire n_11283;
wire n_20003;
wire n_13616;
wire n_20060;
wire n_16729;
wire n_21707;
wire n_3877;
wire n_2494;
wire n_3977;
wire n_13233;
wire n_10677;
wire n_7596;
wire n_20319;
wire n_14211;
wire n_4398;
wire n_8553;
wire n_6490;
wire n_15003;
wire n_10610;
wire n_19318;
wire n_19939;
wire n_20545;
wire n_14572;
wire n_15626;
wire n_5333;
wire n_15724;
wire n_1303;
wire n_14851;
wire n_21414;
wire n_8518;
wire n_6802;
wire n_7527;
wire n_5570;
wire n_3736;
wire n_9514;
wire n_19936;
wire n_18991;
wire n_9402;
wire n_12634;
wire n_20502;
wire n_8364;
wire n_253;
wire n_9005;
wire n_1661;
wire n_8621;
wire n_6167;
wire n_15231;
wire n_8993;
wire n_4701;
wire n_14545;
wire n_19863;
wire n_7101;
wire n_12398;
wire n_6948;
wire n_16861;
wire n_9921;
wire n_20547;
wire n_8910;
wire n_18502;
wire n_15364;
wire n_19512;
wire n_11855;
wire n_14930;
wire n_11667;
wire n_6765;
wire n_7577;
wire n_18485;
wire n_13738;
wire n_19178;
wire n_18840;
wire n_3533;
wire n_17259;
wire n_19032;
wire n_2148;
wire n_393;
wire n_12292;
wire n_18892;
wire n_421;
wire n_15536;
wire n_13346;
wire n_9982;
wire n_12056;
wire n_13149;
wire n_8508;
wire n_20944;
wire n_14179;
wire n_15262;
wire n_12811;
wire n_19597;
wire n_13100;
wire n_14821;
wire n_5886;
wire n_7080;
wire n_7744;
wire n_12897;
wire n_8034;
wire n_17179;
wire n_17447;
wire n_10970;
wire n_14401;
wire n_708;
wire n_14363;
wire n_6960;
wire n_19283;
wire n_13840;
wire n_11983;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_193;
wire n_13389;
wire n_5785;
wire n_4538;
wire n_11680;
wire n_20128;
wire n_6010;
wire n_11446;
wire n_9225;
wire n_18593;
wire n_1742;
wire n_11972;
wire n_14247;
wire n_5376;
wire n_13862;
wire n_16674;
wire n_21437;
wire n_7292;
wire n_15987;
wire n_13486;
wire n_21897;
wire n_1155;
wire n_16936;
wire n_8507;
wire n_2917;
wire n_14323;
wire n_4150;
wire n_827;
wire n_14667;
wire n_21684;
wire n_6265;
wire n_1650;
wire n_8661;
wire n_4985;
wire n_6373;
wire n_20668;
wire n_8573;
wire n_3922;
wire n_3846;
wire n_7692;
wire n_6887;
wire n_11343;
wire n_13277;
wire n_2498;
wire n_19487;
wire n_14366;
wire n_2630;
wire n_16750;
wire n_8136;
wire n_2430;
wire n_14650;
wire n_14657;
wire n_5508;
wire n_12424;
wire n_7440;
wire n_840;
wire n_4852;
wire n_7758;
wire n_11639;
wire n_13528;
wire n_13419;
wire n_17621;
wire n_14087;
wire n_10832;
wire n_12490;
wire n_15053;
wire n_3139;
wire n_14656;
wire n_14757;
wire n_8075;
wire n_20660;
wire n_1890;
wire n_9675;
wire n_8071;
wire n_17929;
wire n_15766;
wire n_16064;
wire n_17266;
wire n_21926;
wire n_13347;
wire n_4515;
wire n_4351;
wire n_14547;
wire n_11795;
wire n_9537;
wire n_10833;
wire n_7413;
wire n_15381;
wire n_1663;
wire n_19970;
wire n_8630;
wire n_7622;
wire n_11266;
wire n_11151;
wire n_7353;
wire n_10071;
wire n_21276;
wire n_15654;
wire n_14992;
wire n_19502;
wire n_15811;
wire n_21535;
wire n_21766;
wire n_6965;
wire n_21248;
wire n_1489;
wire n_8314;
wire n_16279;
wire n_6032;
wire n_21254;
wire n_15729;
wire n_13094;
wire n_7174;
wire n_6402;
wire n_19858;
wire n_7166;
wire n_15495;
wire n_8209;
wire n_2448;
wire n_9654;
wire n_8560;
wire n_17039;
wire n_7591;
wire n_15500;
wire n_5775;
wire n_14139;
wire n_2748;
wire n_3272;
wire n_2717;
wire n_16453;
wire n_21732;
wire n_3691;
wire n_3628;
wire n_19543;
wire n_4235;
wire n_16288;
wire n_21893;
wire n_10183;
wire n_14674;
wire n_18224;
wire n_12704;
wire n_11237;
wire n_11741;
wire n_14130;
wire n_14402;
wire n_15839;
wire n_17924;
wire n_20875;
wire n_8457;
wire n_10549;
wire n_8248;
wire n_7966;
wire n_7070;
wire n_15775;
wire n_19749;
wire n_11721;
wire n_17828;
wire n_17711;
wire n_12245;
wire n_21142;
wire n_751;
wire n_6084;
wire n_10301;
wire n_15888;
wire n_9496;
wire n_21336;
wire n_18384;
wire n_7157;
wire n_6472;
wire n_11097;
wire n_10394;
wire n_17158;
wire n_11105;
wire n_12647;
wire n_12377;
wire n_9251;
wire n_15906;
wire n_2691;
wire n_16398;
wire n_12316;
wire n_6567;
wire n_19554;
wire n_6771;
wire n_2526;
wire n_10182;
wire n_15037;
wire n_12399;
wire n_18641;
wire n_15189;
wire n_17495;
wire n_6910;
wire n_16725;
wire n_5541;
wire n_2709;
wire n_15868;
wire n_19005;
wire n_21082;
wire n_21502;
wire n_5935;
wire n_4865;
wire n_11219;
wire n_1344;
wire n_18672;
wire n_18493;
wire n_1339;
wire n_17960;
wire n_3518;
wire n_3733;
wire n_16886;
wire n_19134;
wire n_17925;
wire n_16593;
wire n_12379;
wire n_12257;
wire n_3738;
wire n_17089;
wire n_5995;
wire n_12246;
wire n_18285;
wire n_21640;
wire n_14099;
wire n_6331;
wire n_6006;
wire n_8421;
wire n_4417;
wire n_14855;
wire n_402;
wire n_6872;
wire n_20311;
wire n_1502;
wire n_15858;
wire n_21144;
wire n_1012;
wire n_7754;
wire n_17332;
wire n_12272;
wire n_6990;
wire n_14885;
wire n_277;
wire n_21608;
wire n_18092;
wire n_6830;
wire n_12662;
wire n_20198;
wire n_7939;
wire n_8675;
wire n_14889;
wire n_1193;
wire n_9375;
wire n_3118;
wire n_8858;
wire n_1226;
wire n_3443;
wire n_20147;
wire n_10296;
wire n_17831;
wire n_3644;
wire n_5076;
wire n_17739;
wire n_3562;
wire n_21216;
wire n_4750;
wire n_20633;
wire n_18168;
wire n_1515;
wire n_17688;
wire n_21031;
wire n_12031;
wire n_11743;
wire n_14274;
wire n_2918;
wire n_10512;
wire n_13658;
wire n_2112;
wire n_2958;
wire n_4981;
wire n_9985;
wire n_17473;
wire n_2394;
wire n_17344;
wire n_3612;
wire n_2954;
wire n_4430;
wire n_6439;
wire n_10026;
wire n_9355;
wire n_17286;
wire n_10041;
wire n_1103;
wire n_16210;
wire n_8102;
wire n_312;
wire n_17939;
wire n_18588;
wire n_4894;
wire n_5780;
wire n_8460;
wire n_3238;
wire n_21959;
wire n_3210;
wire n_16088;
wire n_14234;
wire n_3267;
wire n_13752;
wire n_4995;
wire n_15093;
wire n_14360;
wire n_17910;
wire n_9875;
wire n_10593;
wire n_5524;
wire n_14827;
wire n_229;
wire n_20793;
wire n_10597;
wire n_9963;
wire n_437;
wire n_9582;
wire n_12172;
wire n_10817;
wire n_6465;
wire n_20268;
wire n_16459;
wire n_19619;
wire n_12049;
wire n_13973;
wire n_13229;
wire n_2525;
wire n_11687;
wire n_9732;
wire n_13070;
wire n_14440;
wire n_8699;
wire n_2820;
wire n_14946;
wire n_269;
wire n_13878;
wire n_19640;
wire n_9992;
wire n_2719;
wire n_4057;
wire n_15899;
wire n_16488;
wire n_19572;
wire n_3809;
wire n_7545;
wire n_1448;
wire n_8438;
wire n_14831;
wire n_6194;
wire n_20934;
wire n_3939;
wire n_5401;
wire n_21054;
wire n_8095;
wire n_7537;
wire n_3212;
wire n_13690;
wire n_1433;
wire n_10746;
wire n_10339;
wire n_15572;
wire n_18121;
wire n_319;
wire n_11559;
wire n_14629;
wire n_18474;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_8112;
wire n_12835;
wire n_14727;
wire n_20848;
wire n_5883;
wire n_18734;
wire n_20375;
wire n_1018;
wire n_13432;
wire n_15800;
wire n_21308;
wire n_16161;
wire n_713;
wire n_9090;
wire n_166;
wire n_10684;
wire n_3159;
wire n_17440;
wire n_9226;
wire n_9018;
wire n_12336;
wire n_10949;
wire n_21121;
wire n_12044;
wire n_11727;
wire n_12905;
wire n_8878;
wire n_4604;
wire n_5223;
wire n_14018;
wire n_6620;
wire n_3179;
wire n_17633;
wire n_15348;
wire n_11725;
wire n_15565;
wire n_10279;
wire n_667;
wire n_18460;
wire n_15138;
wire n_7060;
wire n_15643;
wire n_1007;
wire n_6885;
wire n_2369;
wire n_12495;
wire n_2927;
wire n_19961;
wire n_17083;
wire n_18147;
wire n_5364;
wire n_19631;
wire n_16207;
wire n_3064;
wire n_21234;
wire n_13506;
wire n_4639;
wire n_3663;
wire n_12654;
wire n_18939;
wire n_15017;
wire n_6423;
wire n_1535;
wire n_7233;
wire n_10228;
wire n_18786;
wire n_6558;
wire n_8522;
wire n_18857;
wire n_7352;
wire n_951;
wire n_21836;
wire n_18834;
wire n_2069;
wire n_7246;
wire n_19574;
wire n_11807;
wire n_14907;
wire n_15678;
wire n_1563;
wire n_11998;
wire n_4227;
wire n_15562;
wire n_18763;
wire n_10643;
wire n_7056;
wire n_8727;
wire n_15333;
wire n_2482;
wire n_10389;
wire n_10423;
wire n_16573;
wire n_14042;
wire n_11080;
wire n_7729;
wire n_20838;
wire n_5987;
wire n_7740;
wire n_6180;
wire n_6925;
wire n_5919;
wire n_579;
wire n_1698;
wire n_2329;
wire n_8206;
wire n_18539;
wire n_2142;
wire n_11940;
wire n_6176;
wire n_13727;
wire n_16009;
wire n_13986;
wire n_15520;
wire n_10250;
wire n_19802;
wire n_20856;
wire n_12176;
wire n_19362;
wire n_2058;
wire n_2458;
wire n_17826;
wire n_15105;
wire n_3786;
wire n_16123;
wire n_15644;
wire n_371;
wire n_5742;
wire n_8649;
wire n_17416;
wire n_8684;
wire n_21932;
wire n_18093;
wire n_10828;
wire n_17745;
wire n_11139;
wire n_21545;
wire n_2669;
wire n_1778;
wire n_9139;
wire n_2306;
wire n_6614;
wire n_15059;
wire n_16148;
wire n_7839;
wire n_10996;
wire n_12795;
wire n_21973;
wire n_2566;
wire n_12045;
wire n_10636;
wire n_7301;
wire n_9041;
wire n_9643;
wire n_8904;
wire n_20434;
wire n_3060;
wire n_7794;
wire n_11479;
wire n_7366;
wire n_8184;
wire n_5605;
wire n_1984;
wire n_21316;
wire n_2408;
wire n_7025;
wire n_5320;
wire n_1877;
wire n_6947;
wire n_20916;
wire n_9648;
wire n_4485;
wire n_9376;
wire n_183;
wire n_7309;
wire n_9288;
wire n_15507;
wire n_7860;
wire n_6735;
wire n_2659;
wire n_12500;
wire n_7911;
wire n_578;
wire n_15455;
wire n_8530;
wire n_9278;
wire n_344;
wire n_11227;
wire n_9456;
wire n_3089;
wire n_15532;
wire n_19526;
wire n_14925;
wire n_13206;
wire n_16869;
wire n_14123;
wire n_12922;
wire n_496;
wire n_21852;
wire n_20396;
wire n_20866;
wire n_7610;
wire n_663;
wire n_11813;
wire n_5903;
wire n_2682;
wire n_6371;
wire n_18978;
wire n_16973;
wire n_20797;
wire n_8643;
wire n_4569;
wire n_6468;
wire n_11134;
wire n_3436;
wire n_11716;
wire n_8825;
wire n_14548;
wire n_1064;
wire n_16652;
wire n_18169;
wire n_12208;
wire n_20698;
wire n_17873;
wire n_18446;
wire n_19674;
wire n_2868;
wire n_9237;
wire n_20515;
wire n_6850;
wire n_18012;
wire n_19547;
wire n_16612;
wire n_7119;
wire n_13728;
wire n_10714;
wire n_15358;
wire n_19094;
wire n_461;
wire n_5328;
wire n_20813;
wire n_14634;
wire n_4503;
wire n_3507;
wire n_6959;
wire n_19270;
wire n_6909;
wire n_16329;
wire n_1211;
wire n_14613;
wire n_13567;
wire n_15912;
wire n_7006;
wire n_12351;
wire n_907;
wire n_15659;
wire n_17885;
wire n_20616;
wire n_2356;
wire n_488;
wire n_7068;
wire n_14573;
wire n_4556;
wire n_11084;
wire n_6322;
wire n_8668;
wire n_13301;
wire n_16327;
wire n_13492;
wire n_14376;
wire n_16924;
wire n_2620;
wire n_10326;
wire n_14728;
wire n_7526;
wire n_7376;
wire n_7268;
wire n_16198;
wire n_7044;
wire n_12452;
wire n_4327;
wire n_230;
wire n_16357;
wire n_953;
wire n_16335;
wire n_2150;
wire n_10047;
wire n_16319;
wire n_1052;
wire n_12633;
wire n_5573;
wire n_11253;
wire n_18528;
wire n_12936;
wire n_12035;
wire n_13928;
wire n_20717;
wire n_9196;
wire n_13947;
wire n_17594;
wire n_534;
wire n_20757;
wire n_21724;
wire n_15462;
wire n_12915;
wire n_4990;
wire n_21804;
wire n_17582;
wire n_12275;
wire n_10784;
wire n_12947;
wire n_18525;
wire n_9589;
wire n_5800;
wire n_17599;
wire n_16344;
wire n_19082;
wire n_12308;
wire n_1387;
wire n_18510;
wire n_21273;
wire n_1156;
wire n_20352;
wire n_7431;
wire n_21212;
wire n_7654;
wire n_2798;
wire n_16330;
wire n_21633;
wire n_847;
wire n_13379;
wire n_17724;
wire n_10313;
wire n_14983;
wire n_6290;
wire n_9983;
wire n_3655;
wire n_12700;
wire n_8182;
wire n_2548;
wire n_15540;
wire n_13672;
wire n_11204;
wire n_3640;
wire n_20700;
wire n_12985;
wire n_4206;
wire n_16911;
wire n_18343;
wire n_7441;
wire n_13470;
wire n_12788;
wire n_16597;
wire n_11485;
wire n_9962;
wire n_18473;
wire n_17559;
wire n_8007;
wire n_3944;
wire n_12752;
wire n_7394;
wire n_18660;
wire n_8311;
wire n_12194;
wire n_20474;
wire n_4837;
wire n_7022;
wire n_3042;
wire n_21952;
wire n_16306;
wire n_1942;
wire n_9829;
wire n_2510;
wire n_4219;
wire n_21846;
wire n_3659;
wire n_2120;
wire n_411;
wire n_10121;
wire n_1876;
wire n_20027;
wire n_14417;
wire n_14652;
wire n_14002;
wire n_13099;
wire n_7879;
wire n_4438;
wire n_16242;
wire n_2222;
wire n_3510;
wire n_7985;
wire n_16221;
wire n_17338;
wire n_9045;
wire n_9466;
wire n_6515;
wire n_21691;
wire n_16650;
wire n_7935;
wire n_15783;
wire n_13595;
wire n_14358;
wire n_15140;
wire n_21954;
wire n_6984;
wire n_19046;
wire n_1733;
wire n_15167;
wire n_13212;
wire n_851;
wire n_16138;
wire n_10018;
wire n_8987;
wire n_4133;
wire n_3775;
wire n_7256;
wire n_12391;
wire n_17147;
wire n_7595;
wire n_18439;
wire n_9239;
wire n_6183;
wire n_13341;
wire n_16034;
wire n_10051;
wire n_547;
wire n_4030;
wire n_14796;
wire n_16906;
wire n_7380;
wire n_19348;
wire n_12356;
wire n_1710;
wire n_2928;
wire n_8960;
wire n_1734;
wire n_4820;
wire n_14133;
wire n_17712;
wire n_5094;
wire n_18350;
wire n_11107;
wire n_4938;
wire n_16505;
wire n_3469;
wire n_9693;
wire n_15378;
wire n_372;
wire n_677;
wire n_9477;
wire n_15761;
wire n_314;
wire n_4641;
wire n_5548;
wire n_21335;
wire n_10822;
wire n_8895;
wire n_1008;
wire n_15927;
wire n_3158;
wire n_2623;
wire n_11173;
wire n_4078;
wire n_11922;
wire n_16115;
wire n_568;
wire n_18187;
wire n_8867;
wire n_20836;
wire n_1832;
wire n_9599;
wire n_18639;
wire n_3666;
wire n_16382;
wire n_3288;
wire n_13075;
wire n_20876;
wire n_4404;
wire n_5091;
wire n_10903;
wire n_13562;
wire n_1987;
wire n_11868;
wire n_5486;
wire n_21177;
wire n_6611;
wire n_10543;
wire n_18778;
wire n_9449;
wire n_15098;
wire n_20512;
wire n_2545;
wire n_11260;
wire n_18930;
wire n_21378;
wire n_906;
wire n_919;
wire n_20884;
wire n_19741;
wire n_4356;
wire n_12252;
wire n_18984;
wire n_11981;
wire n_15831;
wire n_4432;
wire n_21277;
wire n_13534;
wire n_13750;
wire n_13275;
wire n_13331;
wire n_20297;
wire n_16425;
wire n_535;
wire n_13536;
wire n_20623;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_21214;
wire n_6310;
wire n_7840;
wire n_17796;
wire n_20501;
wire n_14607;
wire n_1692;
wire n_11797;
wire n_7429;
wire n_8948;
wire n_2507;
wire n_9754;
wire n_16898;
wire n_17888;
wire n_457;
wire n_7017;
wire n_4637;
wire n_13249;
wire n_6365;
wire n_21057;
wire n_14225;
wire n_19266;
wire n_20471;
wire n_20729;
wire n_5608;
wire n_3741;
wire n_12455;
wire n_18629;
wire n_10136;
wire n_14759;
wire n_21894;
wire n_11758;
wire n_2029;
wire n_19109;
wire n_21011;
wire n_19568;
wire n_17355;
wire n_1609;
wire n_11162;
wire n_7887;
wire n_1887;
wire n_12559;
wire n_9177;
wire n_6777;
wire n_12614;
wire n_19489;
wire n_12797;
wire n_14396;
wire n_8722;
wire n_12429;
wire n_19756;
wire n_6945;
wire n_9350;
wire n_1721;
wire n_5726;
wire n_7637;
wire n_10454;
wire n_3672;
wire n_13105;
wire n_3109;
wire n_11374;
wire n_12146;
wire n_7321;
wire n_10501;
wire n_15796;
wire n_10766;
wire n_13533;
wire n_11999;
wire n_6583;
wire n_18841;
wire n_6936;
wire n_16742;
wire n_3897;
wire n_8742;
wire n_12921;
wire n_16006;
wire n_6882;
wire n_16893;
wire n_21622;
wire n_19584;
wire n_10288;
wire n_7362;
wire n_19605;
wire n_9960;
wire n_5589;
wire n_13060;
wire n_2179;
wire n_10776;
wire n_11611;
wire n_9785;
wire n_17765;
wire n_16818;
wire n_17700;
wire n_5712;
wire n_1420;
wire n_1132;
wire n_3330;
wire n_4774;
wire n_18849;
wire n_18076;
wire n_2477;
wire n_13563;
wire n_22000;
wire n_7542;
wire n_4093;
wire n_17723;
wire n_7147;
wire n_14653;
wire n_20988;
wire n_15601;
wire n_16440;
wire n_652;
wire n_17181;
wire n_1365;
wire n_6980;
wire n_19592;
wire n_9457;
wire n_15071;
wire n_288;
wire n_18972;
wire n_7889;
wire n_3929;
wire n_19537;
wire n_20805;
wire n_893;
wire n_6341;
wire n_10012;
wire n_1941;
wire n_8444;
wire n_8654;
wire n_10035;
wire n_16579;
wire n_20982;
wire n_504;
wire n_6697;
wire n_5652;
wire n_15577;
wire n_4110;
wire n_3189;
wire n_15752;
wire n_6449;
wire n_17405;
wire n_3154;
wire n_1551;
wire n_19898;
wire n_21760;
wire n_19309;
wire n_10099;
wire n_8449;
wire n_1217;
wire n_2220;
wire n_10985;
wire n_628;
wire n_9224;
wire n_2410;
wire n_12671;
wire n_970;
wire n_10377;
wire n_6036;
wire n_21749;
wire n_18303;
wire n_21568;
wire n_21822;
wire n_10801;
wire n_8443;
wire n_9756;
wire n_7222;
wire n_6071;
wire n_13435;
wire n_3525;
wire n_8271;
wire n_9594;
wire n_3995;
wire n_9277;
wire n_4036;
wire n_20867;
wire n_21657;
wire n_20589;
wire n_921;
wire n_1795;
wire n_19417;
wire n_7400;
wire n_16290;
wire n_19891;
wire n_10000;
wire n_16670;
wire n_14738;
wire n_3478;
wire n_13816;
wire n_21618;
wire n_12323;
wire n_14767;
wire n_21215;
wire n_5616;
wire n_1708;
wire n_16761;
wire n_19618;
wire n_17832;
wire n_7859;
wire n_8900;
wire n_17987;
wire n_6522;
wire n_14057;
wire n_20629;
wire n_6732;
wire n_18240;
wire n_13806;
wire n_21310;
wire n_6562;
wire n_21238;
wire n_17659;
wire n_20196;
wire n_21410;
wire n_1757;
wire n_21060;
wire n_890;
wire n_960;
wire n_15656;
wire n_20535;
wire n_1290;
wire n_20548;
wire n_8344;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_1252;
wire n_8822;
wire n_3784;
wire n_3195;
wire n_9758;
wire n_7212;
wire n_3678;
wire n_7908;
wire n_15160;
wire n_20635;
wire n_17074;
wire n_3456;
wire n_10479;
wire n_18111;
wire n_9876;
wire n_5628;
wire n_18875;
wire n_10277;
wire n_18570;
wire n_4428;
wire n_146;
wire n_18943;
wire n_6689;
wire n_14858;
wire n_13724;
wire n_6143;
wire n_3166;
wire n_21350;
wire n_18863;
wire n_16791;
wire n_3979;
wire n_4582;
wire n_5981;
wire n_12896;
wire n_6095;
wire n_10429;
wire n_22009;
wire n_16966;
wire n_6247;
wire n_21709;
wire n_9257;
wire n_15141;
wire n_9270;
wire n_21584;
wire n_6880;
wire n_10901;
wire n_3749;
wire n_10101;
wire n_14000;
wire n_13422;
wire n_13633;
wire n_17958;
wire n_17585;
wire n_14741;
wire n_14972;
wire n_20798;
wire n_4096;
wire n_12030;
wire n_14679;
wire n_2881;
wire n_8400;
wire n_21143;
wire n_1763;
wire n_13989;
wire n_1966;
wire n_14859;
wire n_321;
wire n_18964;
wire n_6946;
wire n_11593;
wire n_15904;
wire n_11773;
wire n_14074;
wire n_5759;
wire n_15056;
wire n_7484;
wire n_11896;
wire n_20607;
wire n_7231;
wire n_13707;
wire n_20411;
wire n_7272;
wire n_4106;
wire n_17523;
wire n_21541;
wire n_3052;
wire n_7324;
wire n_6693;
wire n_10931;
wire n_8541;
wire n_3743;
wire n_20357;
wire n_12000;
wire n_18104;
wire n_19659;
wire n_11159;
wire n_1932;
wire n_21225;
wire n_17445;
wire n_13001;
wire n_7635;
wire n_13842;
wire n_16568;
wire n_4029;
wire n_19393;
wire n_900;
wire n_21312;
wire n_3870;
wire n_11083;
wire n_10382;
wire n_13664;
wire n_1977;
wire n_2153;
wire n_6235;
wire n_9870;
wire n_4338;
wire n_6504;
wire n_13900;
wire n_3952;
wire n_8638;
wire n_2860;
wire n_7184;
wire n_11090;
wire n_19474;
wire n_1470;
wire n_2318;
wire n_19422;
wire n_14784;
wire n_7491;
wire n_15866;
wire n_2974;
wire n_1940;
wire n_10488;
wire n_13084;
wire n_1114;
wire n_7479;
wire n_13203;
wire n_1176;
wire n_5940;
wire n_8170;
wire n_20350;
wire n_16379;
wire n_17696;
wire n_21884;
wire n_7807;
wire n_8589;
wire n_4107;
wire n_17348;
wire n_11094;
wire n_18353;
wire n_5555;
wire n_6914;
wire n_7978;
wire n_20595;
wire n_15379;
wire n_15441;
wire n_12195;
wire n_15115;
wire n_17695;
wire n_5576;
wire n_6840;
wire n_3898;
wire n_6871;
wire n_11590;
wire n_17618;
wire n_11845;
wire n_9126;
wire n_19089;
wire n_19328;
wire n_5308;
wire n_18410;
wire n_4274;
wire n_16749;
wire n_18918;
wire n_20929;
wire n_14490;
wire n_17882;
wire n_3684;
wire n_11136;
wire n_3137;
wire n_7048;
wire n_11142;
wire n_16843;
wire n_13569;
wire n_18247;
wire n_19374;
wire n_20326;
wire n_5578;
wire n_1173;
wire n_13010;
wire n_14375;
wire n_1401;
wire n_18977;
wire n_20332;
wire n_20449;
wire n_10805;
wire n_1998;
wire n_19124;
wire n_4686;
wire n_21736;
wire n_11414;
wire n_20187;
wire n_21981;
wire n_3759;
wire n_14322;
wire n_18223;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_10528;
wire n_5741;
wire n_8570;
wire n_5991;
wire n_13815;
wire n_3933;
wire n_3206;
wire n_7928;
wire n_12201;
wire n_17894;
wire n_5243;
wire n_5449;
wire n_16415;
wire n_13924;
wire n_1122;
wire n_10625;
wire n_9545;
wire n_4233;
wire n_7099;
wire n_10557;
wire n_19206;
wire n_4709;
wire n_16125;
wire n_13002;
wire n_14732;
wire n_19984;
wire n_6657;
wire n_8129;
wire n_2542;
wire n_15521;
wire n_1174;
wire n_4625;
wire n_18675;
wire n_21663;
wire n_17953;
wire n_11883;
wire n_17479;
wire n_8259;
wire n_2063;
wire n_3803;
wire n_2252;
wire n_9056;
wire n_8094;
wire n_10357;
wire n_8572;
wire n_2576;
wire n_21302;
wire n_7588;
wire n_17578;
wire n_3746;
wire n_11241;
wire n_9172;
wire n_12441;
wire n_9145;
wire n_210;
wire n_8099;
wire n_774;
wire n_2493;
wire n_8770;
wire n_5078;
wire n_16039;
wire n_2885;
wire n_14250;
wire n_20323;
wire n_12827;
wire n_9920;
wire n_3485;
wire n_18376;
wire n_7378;
wire n_15689;
wire n_11152;
wire n_2845;
wire n_6144;
wire n_17059;
wire n_20313;
wire n_10147;
wire n_4616;
wire n_13765;
wire n_15962;
wire n_21272;
wire n_17133;
wire n_11990;
wire n_14554;
wire n_17899;
wire n_10889;
wire n_12363;
wire n_15788;
wire n_14699;
wire n_1930;
wire n_1955;
wire n_10816;
wire n_16428;
wire n_13385;
wire n_10032;
wire n_17756;
wire n_10898;
wire n_5856;
wire n_20084;
wire n_19550;
wire n_4895;
wire n_9735;
wire n_21122;
wire n_21337;
wire n_15569;
wire n_15078;
wire n_1482;
wire n_6413;
wire n_7679;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_13608;
wire n_10680;
wire n_7783;
wire n_5684;
wire n_21333;
wire n_21174;
wire n_4789;
wire n_19897;
wire n_10675;
wire n_19291;
wire n_3217;
wire n_3425;
wire n_16117;
wire n_13829;
wire n_5890;
wire n_16409;
wire n_7820;
wire n_7833;
wire n_8820;
wire n_21911;
wire n_14750;
wire n_15454;
wire n_21171;
wire n_7643;
wire n_12460;
wire n_13586;
wire n_12821;
wire n_9922;
wire n_6712;
wire n_8781;
wire n_19462;
wire n_8000;
wire n_10961;
wire n_19624;
wire n_5839;
wire n_4418;
wire n_2549;
wire n_21166;
wire n_20975;
wire n_12361;
wire n_1318;
wire n_8575;
wire n_17369;
wire n_12593;
wire n_6474;
wire n_1454;
wire n_3723;
wire n_8670;
wire n_20716;
wire n_6573;
wire n_13151;
wire n_6053;
wire n_14380;
wire n_7234;
wire n_21114;
wire n_1388;
wire n_20215;
wire n_7930;
wire n_1625;
wire n_19301;
wire n_5167;
wire n_8934;
wire n_4913;
wire n_19622;
wire n_15928;
wire n_21504;
wire n_15485;
wire n_6685;
wire n_19234;
wire n_18079;
wire n_2850;
wire n_11964;
wire n_1817;
wire n_19049;
wire n_2654;
wire n_4621;
wire n_10158;
wire n_3176;
wire n_11933;
wire n_10043;
wire n_18001;
wire n_6253;
wire n_17753;
wire n_19894;
wire n_15575;
wire n_3581;
wire n_4077;
wire n_10930;
wire n_16408;
wire n_2221;
wire n_1024;
wire n_16406;
wire n_1564;
wire n_18160;
wire n_5214;
wire n_13551;
wire n_19050;
wire n_12461;
wire n_3879;
wire n_12893;
wire n_17876;
wire n_8790;
wire n_11624;
wire n_18010;
wire n_20480;
wire n_13791;
wire n_7190;
wire n_13807;
wire n_13142;
wire n_11560;
wire n_1772;
wire n_13678;
wire n_1476;
wire n_13433;
wire n_20488;
wire n_3646;
wire n_18554;
wire n_4546;
wire n_17572;
wire n_862;
wire n_6356;
wire n_18309;
wire n_19575;
wire n_16703;
wire n_11616;
wire n_18723;
wire n_14746;
wire n_21365;
wire n_19196;
wire n_6514;
wire n_7369;
wire n_21269;
wire n_1554;
wire n_10159;
wire n_9210;
wire n_21961;
wire n_7359;
wire n_20492;
wire n_15443;
wire n_10462;
wire n_8756;
wire n_19798;
wire n_16351;
wire n_2345;
wire n_17208;
wire n_3062;
wire n_16316;
wire n_21207;
wire n_16151;
wire n_1142;
wire n_10350;
wire n_16431;
wire n_9351;
wire n_11179;
wire n_6923;
wire n_11708;
wire n_17027;
wire n_9950;
wire n_10418;
wire n_10336;
wire n_138;
wire n_20953;
wire n_8021;
wire n_12092;
wire n_11240;
wire n_20603;
wire n_13155;
wire n_21910;
wire n_3364;
wire n_21152;
wire n_14565;
wire n_15277;
wire n_3201;
wire n_20917;
wire n_18952;
wire n_20860;
wire n_17379;
wire n_10609;
wire n_17785;
wire n_20339;
wire n_21197;
wire n_6151;
wire n_19968;
wire n_18036;
wire n_20119;
wire n_2874;
wire n_5179;
wire n_6469;
wire n_21294;
wire n_3543;
wire n_15530;
wire n_18432;
wire n_9688;
wire n_12330;
wire n_13597;
wire n_18950;
wire n_19901;
wire n_313;
wire n_12717;
wire n_20254;
wire n_1478;
wire n_8280;
wire n_15119;
wire n_9530;
wire n_2742;
wire n_3314;
wire n_2360;
wire n_19553;
wire n_20630;
wire n_8598;
wire n_20519;
wire n_11178;
wire n_5740;
wire n_17705;
wire n_2834;
wire n_17001;
wire n_517;
wire n_11840;
wire n_5015;
wire n_20091;
wire n_20582;
wire n_5729;
wire n_19551;
wire n_12084;
wire n_2030;
wire n_18517;
wire n_17228;
wire n_1404;
wire n_11472;
wire n_16948;
wire n_4804;
wire n_17651;
wire n_9285;
wire n_12997;
wire n_11295;
wire n_8847;
wire n_11171;
wire n_7051;
wire n_11030;
wire n_13394;
wire n_20063;
wire n_2321;
wire n_6297;
wire n_6975;
wire n_8979;
wire n_12080;
wire n_15514;
wire n_18668;
wire n_5688;
wire n_2612;
wire n_20696;
wire n_10894;
wire n_979;
wire n_19840;
wire n_9393;
wire n_2505;
wire n_4061;
wire n_20533;
wire n_2070;
wire n_270;
wire n_6521;
wire n_2904;
wire n_8355;
wire n_9736;
wire n_13691;
wire n_3004;
wire n_5986;
wire n_3112;
wire n_19431;
wire n_6581;
wire n_14372;
wire n_3874;
wire n_10241;
wire n_7064;
wire n_19411;
wire n_10180;
wire n_19755;
wire n_21988;
wire n_8784;
wire n_14666;
wire n_12335;
wire n_6545;
wire n_19448;
wire n_16974;
wire n_13669;
wire n_575;
wire n_14371;
wire n_8171;
wire n_3266;
wire n_13731;
wire n_7899;
wire n_10370;
wire n_15263;
wire n_9728;
wire n_6065;
wire n_13845;
wire n_1130;
wire n_15475;
wire n_21903;
wire n_9659;
wire n_6987;
wire n_14328;
wire n_4725;
wire n_6190;
wire n_5331;
wire n_14311;
wire n_21408;
wire n_14847;
wire n_11149;
wire n_6623;
wire n_12055;
wire n_15922;
wire n_11707;
wire n_18004;
wire n_12413;
wire n_11086;
wire n_657;
wire n_5814;
wire n_12803;
wire n_16792;
wire n_491;
wire n_15026;
wire n_16709;
wire n_14034;
wire n_566;
wire n_7015;
wire n_5263;
wire n_11772;
wire n_14618;
wire n_19904;
wire n_3444;
wire n_1181;
wire n_11764;
wire n_13904;
wire n_11225;
wire n_5622;
wire n_13648;
wire n_14844;
wire n_11112;
wire n_9723;
wire n_20256;
wire n_21712;
wire n_1969;
wire n_1138;
wire n_5546;
wire n_927;
wire n_14491;
wire n_7143;
wire n_5224;
wire n_14267;
wire n_3688;
wire n_15116;
wire n_21966;
wire n_19347;
wire n_2599;
wire n_15774;
wire n_3338;
wire n_10866;
wire n_10348;
wire n_12991;
wire n_4671;
wire n_20429;
wire n_1271;
wire n_5966;
wire n_11359;
wire n_16318;
wire n_17656;
wire n_7420;
wire n_9681;
wire n_9414;
wire n_1166;
wire n_8607;
wire n_20839;
wire n_21887;
wire n_1508;
wire n_18514;
wire n_3261;
wire n_19280;
wire n_19958;
wire n_3863;
wire n_11830;
wire n_15428;
wire n_17123;
wire n_1150;
wire n_9379;
wire n_17869;
wire n_20725;
wire n_1780;
wire n_17879;
wire n_6605;
wire n_19128;
wire n_21109;
wire n_18482;
wire n_4699;
wire n_16983;
wire n_18009;
wire n_4127;
wire n_544;
wire n_15408;
wire n_17576;
wire n_14751;
wire n_9151;
wire n_3641;
wire n_4577;
wire n_11863;
wire n_18228;
wire n_16651;
wire n_7168;
wire n_7736;
wire n_5000;
wire n_10322;
wire n_1323;
wire n_13952;
wire n_14478;
wire n_2880;
wire n_9701;
wire n_20654;
wire n_8223;
wire n_864;
wire n_7030;
wire n_5420;
wire n_16027;
wire n_1264;
wire n_6311;
wire n_11192;
wire n_11569;
wire n_20861;
wire n_447;
wire n_3407;
wire n_6424;
wire n_6220;
wire n_12769;
wire n_5234;
wire n_16744;
wire n_5835;
wire n_2244;
wire n_16533;
wire n_2257;
wire n_6029;
wire n_18175;
wire n_1607;
wire n_17626;
wire n_15807;
wire n_20355;
wire n_21346;
wire n_3163;
wire n_5440;
wire n_5679;
wire n_5938;
wire n_3710;
wire n_4155;
wire n_2031;
wire n_3891;
wire n_5724;
wire n_17229;
wire n_8793;
wire n_20965;
wire n_11679;
wire n_1124;
wire n_7280;
wire n_2127;
wire n_8489;
wire n_6915;
wire n_18868;
wire n_1104;
wire n_7511;
wire n_6856;
wire n_7941;
wire n_9385;
wire n_19179;
wire n_3834;
wire n_8454;
wire n_10536;
wire n_17032;
wire n_12268;
wire n_7345;
wire n_12656;
wire n_20221;
wire n_21775;
wire n_18293;
wire n_19117;
wire n_20082;
wire n_12678;
wire n_14521;
wire n_1016;
wire n_12876;
wire n_2047;
wire n_13107;
wire n_15667;
wire n_240;
wire n_13523;
wire n_2478;
wire n_19408;
wire n_1483;
wire n_6363;
wire n_18610;
wire n_10620;
wire n_16049;
wire n_13420;
wire n_10079;
wire n_10188;
wire n_8721;
wire n_9391;
wire n_17132;
wire n_6406;
wire n_17619;
wire n_2085;
wire n_13603;
wire n_370;
wire n_15429;
wire n_2782;
wire n_1670;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_20138;
wire n_16296;
wire n_15588;
wire n_10107;
wire n_8664;
wire n_5677;
wire n_5511;
wire n_9719;
wire n_21857;
wire n_17531;
wire n_14507;
wire n_5280;
wire n_6479;
wire n_19636;
wire n_16482;
wire n_12563;
wire n_16845;
wire n_3836;
wire n_12331;
wire n_17648;
wire n_14599;
wire n_15049;
wire n_4187;
wire n_6263;
wire n_1030;
wire n_17871;
wire n_21112;
wire n_1267;
wire n_5419;
wire n_2970;
wire n_12382;
wire n_2235;
wire n_673;
wire n_3980;
wire n_1473;
wire n_11148;
wire n_13286;
wire n_6014;
wire n_20568;
wire n_11396;
wire n_20143;
wire n_17216;
wire n_9775;
wire n_17636;
wire n_14980;
wire n_19062;
wire n_184;
wire n_16164;
wire n_14427;
wire n_3841;
wire n_12107;
wire n_8809;
wire n_20000;
wire n_19412;
wire n_20458;
wire n_17943;
wire n_11009;
wire n_17942;
wire n_6158;
wire n_9709;
wire n_3262;
wire n_8447;
wire n_14202;
wire n_1450;
wire n_4006;
wire n_4861;
wire n_9324;
wire n_13311;
wire n_18769;
wire n_11957;
wire n_11538;
wire n_17923;
wire n_19471;
wire n_11264;
wire n_12774;
wire n_477;
wire n_3191;
wire n_3837;
wire n_17060;
wire n_7145;
wire n_2855;
wire n_17077;
wire n_9657;
wire n_14319;
wire n_9352;
wire n_15917;
wire n_12807;
wire n_3025;
wire n_4674;
wire n_21492;
wire n_15268;
wire n_10113;
wire n_16485;
wire n_11267;
wire n_10990;
wire n_3899;
wire n_14014;
wire n_4159;
wire n_3714;
wire n_11618;
wire n_9969;
wire n_4069;
wire n_19828;
wire n_20409;
wire n_12715;
wire n_14945;
wire n_13814;
wire n_17956;
wire n_12968;
wire n_9618;
wire n_20637;
wire n_10732;
wire n_14257;
wire n_7464;
wire n_2590;
wire n_20146;
wire n_15239;
wire n_2330;
wire n_6759;
wire n_3106;
wire n_3328;
wire n_944;
wire n_3889;
wire n_6139;
wire n_7434;
wire n_13832;
wire n_21837;
wire n_3508;
wire n_9205;
wire n_14630;
wire n_17234;
wire n_5650;
wire n_2636;
wire n_14104;
wire n_19677;
wire n_15482;
wire n_11098;
wire n_2759;
wire n_5552;
wire n_7299;
wire n_15086;
wire n_13281;
wire n_8515;
wire n_17005;
wire n_13556;
wire n_8648;
wire n_9377;
wire n_16395;
wire n_10839;
wire n_11875;
wire n_6800;
wire n_21076;
wire n_2319;
wire n_596;
wire n_9016;
wire n_7503;
wire n_13979;
wire n_18563;
wire n_12514;
wire n_10091;
wire n_7091;
wire n_1838;
wire n_9690;
wire n_1660;
wire n_13400;
wire n_21275;
wire n_14268;
wire n_4090;
wire n_9451;
wire n_10849;
wire n_15456;
wire n_11108;
wire n_9760;
wire n_7555;
wire n_10947;
wire n_16439;
wire n_10272;
wire n_9035;
wire n_12806;
wire n_21292;
wire n_6422;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_14965;
wire n_5521;
wire n_7578;
wire n_5028;
wire n_2350;
wire n_17632;
wire n_4194;
wire n_9070;
wire n_20808;
wire n_14012;
wire n_1571;
wire n_3119;
wire n_7531;
wire n_3479;
wire n_9981;
wire n_19250;
wire n_12235;
wire n_21891;
wire n_6981;
wire n_15647;
wire n_18058;
wire n_4372;
wire n_20506;
wire n_11733;
wire n_13632;
wire n_12471;
wire n_8428;
wire n_9021;
wire n_21933;
wire n_13130;
wire n_21078;
wire n_12083;
wire n_15251;
wire n_19783;
wire n_15156;
wire n_12065;
wire n_9495;
wire n_21747;
wire n_1647;
wire n_12167;
wire n_20351;
wire n_4685;
wire n_5968;
wire n_20132;
wire n_2387;
wire n_21340;
wire n_20553;
wire n_12087;
wire n_17703;
wire n_12243;
wire n_18575;
wire n_4757;
wire n_2913;
wire n_20510;
wire n_20034;
wire n_19226;
wire n_11899;
wire n_1233;
wire n_15842;
wire n_21105;
wire n_15688;
wire n_10583;
wire n_16420;
wire n_293;
wire n_4648;
wire n_14308;
wire n_8269;
wire n_19658;
wire n_21002;
wire n_6081;
wire n_8458;
wire n_13857;
wire n_3823;
wire n_19353;
wire n_4173;
wire n_8499;
wire n_738;
wire n_13315;
wire n_13180;
wire n_16666;
wire n_5404;
wire n_8306;
wire n_610;
wire n_16929;
wire n_12375;
wire n_8167;
wire n_5438;
wire n_19423;
wire n_439;
wire n_4627;
wire n_8613;
wire n_11790;
wire n_19764;
wire n_7354;
wire n_17012;
wire n_13474;
wire n_13224;
wire n_12684;
wire n_9099;
wire n_3369;
wire n_3783;
wire n_20206;
wire n_20403;
wire n_21405;
wire n_15957;
wire n_10952;
wire n_1639;
wire n_12566;
wire n_21364;
wire n_7571;
wire n_13919;
wire n_19224;
wire n_14466;
wire n_16547;
wire n_331;
wire n_2039;
wire n_11518;
wire n_16982;
wire n_19515;
wire n_14061;
wire n_15365;
wire n_21077;
wire n_15615;
wire n_18847;
wire n_11663;
wire n_10991;
wire n_18358;
wire n_9837;
wire n_4855;
wire n_12681;
wire n_3969;
wire n_19982;
wire n_17118;
wire n_17979;
wire n_2459;
wire n_9433;
wire n_6588;
wire n_20706;
wire n_13593;
wire n_14912;
wire n_16976;
wire n_5685;
wire n_11726;
wire n_1923;
wire n_13188;
wire n_10465;
wire n_20280;
wire n_12149;
wire n_8397;
wire n_5374;
wire n_17373;
wire n_19310;
wire n_6621;
wire n_18099;
wire n_18606;
wire n_18826;
wire n_21579;
wire n_10517;
wire n_6323;
wire n_1033;
wire n_18762;
wire n_18789;
wire n_13485;
wire n_16727;
wire n_13355;
wire n_13368;
wire n_13160;
wire n_13676;
wire n_1009;
wire n_21559;
wire n_454;
wire n_3818;
wire n_8294;
wire n_11856;
wire n_16774;
wire n_4387;
wire n_7878;
wire n_15176;
wire n_15972;
wire n_14904;
wire n_8915;
wire n_13006;
wire n_1959;
wire n_9841;
wire n_1574;
wire n_2355;
wire n_12831;
wire n_10582;
wire n_9132;
wire n_18982;
wire n_8855;
wire n_18790;
wire n_1355;
wire n_2565;
wire n_17976;
wire n_12154;
wire n_16653;
wire n_743;
wire n_5948;
wire n_18646;
wire n_10662;
wire n_16586;
wire n_6911;
wire n_3268;
wire n_11512;
wire n_19520;
wire n_18530;
wire n_15555;
wire n_19060;
wire n_13114;
wire n_3614;
wire n_3301;
wire n_8869;
wire n_5900;
wire n_15860;
wire n_16804;
wire n_15731;
wire n_13200;
wire n_2595;
wire n_9063;
wire n_8998;
wire n_18377;
wire n_15652;
wire n_3411;
wire n_7209;
wire n_3586;
wire n_5554;
wire n_17260;
wire n_9926;
wire n_14620;
wire n_17414;
wire n_11907;
wire n_14291;
wire n_14092;
wire n_12796;
wire n_5427;
wire n_15876;
wire n_5639;
wire n_21464;
wire n_10585;
wire n_5417;
wire n_8772;
wire n_12008;
wire n_12279;
wire n_8307;
wire n_224;
wire n_15273;
wire n_3103;
wire n_18884;
wire n_765;
wire n_2424;
wire n_20008;
wire n_16294;
wire n_19545;
wire n_1015;
wire n_15878;
wire n_9263;
wire n_7630;
wire n_11831;
wire n_14766;
wire n_9632;
wire n_19341;
wire n_1106;
wire n_2230;
wire n_9282;
wire n_2490;
wire n_10933;
wire n_12192;
wire n_7410;
wire n_4213;
wire n_2849;
wire n_10546;
wire n_12864;
wire n_9503;
wire n_20963;
wire n_15486;
wire n_13348;
wire n_19896;
wire n_19177;
wire n_18853;
wire n_7495;
wire n_9782;
wire n_9855;
wire n_4929;
wire n_15400;
wire n_8040;
wire n_9347;
wire n_20057;
wire n_10923;
wire n_6079;
wire n_10836;
wire n_6458;
wire n_1354;
wire n_15698;
wire n_1044;
wire n_19382;
wire n_8132;
wire n_2508;
wire n_21609;
wire n_18467;
wire n_13544;
wire n_12792;
wire n_15556;
wire n_16719;
wire n_2416;
wire n_21210;
wire n_9148;
wire n_16757;
wire n_17130;
wire n_13530;
wire n_2461;
wire n_19084;
wire n_14289;
wire n_16588;
wire n_6287;
wire n_572;
wire n_12923;
wire n_9585;
wire n_17249;
wire n_4210;
wire n_16891;
wire n_2555;
wire n_2662;
wire n_16450;
wire n_6851;
wire n_12716;
wire n_2890;
wire n_8356;
wire n_20007;
wire n_21676;
wire n_18505;
wire n_14614;
wire n_3698;
wire n_1840;
wire n_716;
wire n_12463;
wire n_17728;
wire n_21241;
wire n_14484;
wire n_15399;
wire n_6619;
wire n_11456;
wire n_8193;
wire n_17396;
wire n_14536;
wire n_18614;
wire n_6804;
wire n_803;
wire n_9370;
wire n_19746;
wire n_13421;
wire n_2572;
wire n_17734;
wire n_18054;
wire n_7490;
wire n_10578;
wire n_4590;
wire n_13349;
wire n_8329;
wire n_9626;
wire n_14501;
wire n_16073;
wire n_8154;
wire n_16812;
wire n_5456;
wire n_21802;
wire n_18589;
wire n_14825;
wire n_15125;
wire n_15479;
wire n_13488;
wire n_15542;
wire n_5727;
wire n_3290;
wire n_7114;
wire n_19153;
wire n_248;
wire n_2440;
wire n_4883;
wire n_17457;
wire n_12963;
wire n_3264;
wire n_9536;
wire n_14316;
wire n_12620;
wire n_8746;
wire n_20849;
wire n_11411;
wire n_14506;
wire n_21524;
wire n_1085;
wire n_2403;
wire n_18297;
wire n_20443;
wire n_15613;
wire n_9017;
wire n_5407;
wire n_16874;
wire n_4608;
wire n_5232;
wire n_20164;
wire n_7271;
wire n_21682;
wire n_1112;
wire n_18125;
wire n_12213;
wire n_6739;
wire n_10450;
wire n_12397;
wire n_2463;
wire n_9565;
wire n_6666;
wire n_15284;
wire n_18364;
wire n_2993;
wire n_13993;
wire n_385;
wire n_15701;
wire n_7419;
wire n_20563;
wire n_18348;
wire n_1560;
wire n_9337;
wire n_21434;
wire n_15602;
wire n_2037;
wire n_11436;
wire n_7784;
wire n_8714;
wire n_10607;
wire n_6934;
wire n_11463;
wire n_14152;
wire n_1363;
wire n_3482;
wire n_18580;
wire n_10668;
wire n_2233;
wire n_1312;
wire n_10713;
wire n_17233;
wire n_19083;
wire n_21879;
wire n_7864;
wire n_7129;
wire n_5323;
wire n_3572;
wire n_19437;
wire n_992;
wire n_6952;
wire n_7062;
wire n_16166;
wire n_14300;
wire n_9077;
wire n_5941;
wire n_1643;
wire n_5879;
wire n_15340;
wire n_11277;
wire n_15195;
wire n_13777;
wire n_11061;
wire n_18697;
wire n_3423;
wire n_7238;
wire n_12733;
wire n_16560;
wire n_7126;
wire n_9745;
wire n_3854;
wire n_12944;
wire n_2468;
wire n_10309;
wire n_1610;
wire n_1422;
wire n_13190;
wire n_3078;
wire n_18765;
wire n_8482;
wire n_11462;
wire n_17199;
wire n_10024;
wire n_9892;
wire n_16227;
wire n_7405;
wire n_7739;
wire n_19612;
wire n_19616;
wire n_13790;
wire n_8761;
wire n_16418;
wire n_4027;
wire n_7934;
wire n_831;
wire n_14283;
wire n_4599;
wire n_21363;
wire n_21558;
wire n_14492;
wire n_20259;
wire n_15457;
wire n_4628;
wire n_9435;
wire n_5668;
wire n_988;
wire n_4873;
wire n_21382;
wire n_14470;
wire n_16479;
wire n_11403;
wire n_15794;
wire n_6870;
wire n_10520;
wire n_13666;
wire n_2298;
wire n_18671;
wire n_4307;
wire n_635;
wire n_15966;
wire n_2303;
wire n_16193;
wire n_10519;
wire n_7776;
wire n_12966;
wire n_2747;
wire n_20924;
wire n_7059;
wire n_21838;
wire n_7035;
wire n_1848;
wire n_5571;
wire n_11854;
wire n_8029;
wire n_21562;
wire n_5289;
wire n_6713;
wire n_6747;
wire n_13588;
wire n_10289;
wire n_18967;
wire n_14496;
wire n_13261;
wire n_11925;
wire n_20342;
wire n_15855;
wire n_7317;
wire n_14043;
wire n_3712;
wire n_20479;
wire n_11961;
wire n_830;
wire n_21735;
wire n_12433;
wire n_21211;
wire n_10940;
wire n_6262;
wire n_12765;
wire n_1655;
wire n_9023;
wire n_12097;
wire n_10723;
wire n_6412;
wire n_2574;
wire n_7782;
wire n_7220;
wire n_717;
wire n_11824;
wire n_3697;
wire n_19086;
wire n_1232;
wire n_734;
wire n_10161;
wire n_11532;
wire n_4044;
wire n_12728;
wire n_16751;
wire n_16447;
wire n_6684;
wire n_13766;
wire n_13784;
wire n_7065;
wire n_10271;
wire n_1338;
wire n_5510;
wire n_6046;
wire n_1522;
wire n_9733;
wire n_5363;
wire n_5200;
wire n_9502;
wire n_338;
wire n_5659;
wire n_5618;
wire n_6325;
wire n_13374;
wire n_20446;
wire n_10163;
wire n_13824;
wire n_5356;
wire n_16289;
wire n_5258;
wire n_12708;
wire n_5255;
wire n_15202;
wire n_18129;
wire n_19460;
wire n_10576;
wire n_9623;
wire n_10424;
wire n_21795;
wire n_711;
wire n_3517;
wire n_2522;
wire n_16163;
wire n_1834;
wire n_17708;
wire n_19517;
wire n_20388;
wire n_21482;
wire n_7501;
wire n_18783;
wire n_5080;
wire n_1516;
wire n_6665;
wire n_3506;
wire n_19651;
wire n_12372;
wire n_8053;
wire n_13141;
wire n_17434;
wire n_11015;
wire n_5817;
wire n_6690;
wire n_20227;
wire n_10192;
wire n_17959;
wire n_4998;
wire n_19271;
wire n_19767;
wire n_1731;
wire n_8735;
wire n_21445;
wire n_818;
wire n_18908;
wire n_15541;
wire n_10219;
wire n_15722;
wire n_5627;
wire n_16524;
wire n_21748;
wire n_7242;
wire n_3835;
wire n_6461;
wire n_8830;
wire n_2205;
wire n_1777;
wire n_17420;
wire n_3967;
wire n_1912;
wire n_18327;
wire n_6212;
wire n_1410;
wire n_707;
wire n_9532;
wire n_8415;
wire n_19557;
wire n_16873;
wire n_9561;
wire n_16478;
wire n_8547;
wire n_10788;
wire n_6074;
wire n_10910;
wire n_7561;
wire n_1584;
wire n_2164;
wire n_8426;
wire n_9326;
wire n_8672;
wire n_18418;
wire n_20495;
wire n_7994;
wire n_8540;
wire n_15421;
wire n_18542;
wire n_15767;
wire n_5137;
wire n_13705;
wire n_16097;
wire n_3348;
wire n_179;
wire n_7415;
wire n_410;
wire n_20815;
wire n_7793;
wire n_5796;
wire n_6320;
wire n_6068;
wire n_14290;
wire n_3358;
wire n_5791;
wire n_9458;
wire n_10608;
wire n_5098;
wire n_1543;
wire n_9910;
wire n_11014;
wire n_9100;
wire n_11119;
wire n_8816;
wire n_7957;
wire n_8712;
wire n_6831;
wire n_16172;
wire n_3657;
wire n_4924;
wire n_12255;
wire n_13881;
wire n_8663;
wire n_7217;
wire n_2692;
wire n_18501;
wire n_799;
wire n_18106;
wire n_6785;
wire n_8959;
wire n_21200;
wire n_9117;
wire n_6930;
wire n_16623;
wire n_4272;
wire n_1753;
wire n_3278;
wire n_8049;
wire n_6838;
wire n_869;
wire n_12212;
wire n_12126;
wire n_21201;
wire n_12686;
wire n_6443;
wire n_13328;
wire n_6105;
wire n_16236;
wire n_7558;
wire n_14142;
wire n_137;
wire n_18281;
wire n_11628;
wire n_10594;
wire n_3968;
wire n_9398;
wire n_5099;
wire n_11606;
wire n_12749;
wire n_4957;
wire n_15821;
wire n_235;
wire n_19535;
wire n_16405;
wire n_643;
wire n_4072;
wire n_5579;
wire n_19315;
wire n_1115;
wire n_8381;
wire n_16423;
wire n_12079;
wire n_21236;
wire n_4781;
wire n_19405;
wire n_10879;
wire n_2550;
wire n_15090;
wire n_7341;
wire n_467;
wire n_13602;
wire n_4424;
wire n_823;
wire n_17188;
wire n_10792;
wire n_725;
wire n_21093;
wire n_16616;
wire n_20811;
wire n_18770;
wire n_14539;
wire n_3292;
wire n_21059;
wire n_21222;
wire n_3878;
wire n_7646;
wire n_9889;
wire n_3553;
wire n_6169;
wire n_4746;
wire n_13975;
wire n_16391;
wire n_3850;
wire n_13833;
wire n_4459;
wire n_11757;
wire n_13169;
wire n_8614;
wire n_21759;
wire n_17716;
wire n_1320;
wire n_9081;
wire n_7496;
wire n_12446;
wire n_19558;
wire n_13354;
wire n_12856;
wire n_16106;
wire n_10544;
wire n_19824;
wire n_20810;
wire n_5681;
wire n_20465;
wire n_12841;
wire n_8656;
wire n_587;
wire n_19446;
wire n_18193;
wire n_7605;
wire n_11400;
wire n_9696;
wire n_7342;
wire n_19786;
wire n_21678;
wire n_16535;
wire n_14926;
wire n_13297;
wire n_10945;
wire n_14601;
wire n_16679;
wire n_11791;
wire n_10541;
wire n_12196;
wire n_11910;
wire n_1330;
wire n_3072;
wire n_21219;
wire n_9426;
wire n_18568;
wire n_18171;
wire n_8143;
wire n_14027;
wire n_18886;
wire n_6462;
wire n_21912;
wire n_9896;
wire n_9650;
wire n_16541;
wire n_20020;
wire n_20511;
wire n_18213;
wire n_16218;
wire n_11974;
wire n_20052;
wire n_20231;
wire n_14730;
wire n_1083;
wire n_15207;
wire n_20768;
wire n_5483;
wire n_17488;
wire n_9055;
wire n_13585;
wire n_6916;
wire n_20217;
wire n_17951;
wire n_3904;
wire n_5150;
wire n_16899;
wire n_17706;
wire n_5075;
wire n_16907;
wire n_18331;
wire n_18259;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_8236;
wire n_11547;
wire n_21620;
wire n_18478;
wire n_12676;
wire n_19349;
wire n_21844;
wire n_18351;
wire n_7949;
wire n_1498;
wire n_21360;
wire n_19975;
wire n_4225;
wire n_17361;
wire n_16760;
wire n_10020;
wire n_2567;
wire n_19429;
wire n_5142;
wire n_21462;
wire n_18072;
wire n_9839;
wire n_15816;
wire n_4300;
wire n_20741;
wire n_432;
wire n_1769;
wire n_4783;
wire n_14254;
wire n_14044;
wire n_7579;
wire n_21198;
wire n_2673;
wire n_15393;
wire n_4267;
wire n_8139;
wire n_7917;
wire n_5951;
wire n_10907;
wire n_2442;
wire n_21577;
wire n_11256;
wire n_19486;
wire n_9658;
wire n_12124;
wire n_19794;
wire n_17872;
wire n_14004;
wire n_8156;
wire n_15446;
wire n_14913;
wire n_12189;
wire n_7886;
wire n_6154;
wire n_6020;
wire n_12310;
wire n_2912;
wire n_16728;
wire n_13821;
wire n_21872;
wire n_1315;
wire n_18142;
wire n_10706;
wire n_10774;
wire n_16467;
wire n_1910;
wire n_3955;
wire n_11963;
wire n_10744;
wire n_8645;
wire n_7774;
wire n_8189;
wire n_4839;
wire n_13810;
wire n_17736;
wire n_6210;
wire n_17225;
wire n_3435;
wire n_19229;
wire n_20157;
wire n_14399;
wire n_10083;
wire n_15561;
wire n_12918;
wire n_11825;
wire n_18724;
wire n_7670;
wire n_4923;
wire n_14126;
wire n_20270;
wire n_5971;
wire n_4083;
wire n_13532;
wire n_12223;
wire n_8018;
wire n_6640;
wire n_20025;
wire n_3916;
wire n_13335;
wire n_2569;
wire n_18621;
wire n_3556;
wire n_2196;
wire n_7721;
wire n_16965;
wire n_18050;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_19736;
wire n_5169;
wire n_4389;
wire n_17110;
wire n_20672;
wire n_12143;
wire n_19332;
wire n_20439;
wire n_11493;
wire n_2083;
wire n_10281;
wire n_6718;
wire n_9685;
wire n_20436;
wire n_6542;
wire n_10126;
wire n_10759;
wire n_11786;
wire n_21126;
wire n_5568;
wire n_403;
wire n_11722;
wire n_16667;
wire n_21592;
wire n_10092;
wire n_8635;
wire n_6763;
wire n_9567;
wire n_3194;
wire n_2414;
wire n_13614;
wire n_20045;
wire n_9059;
wire n_17352;
wire n_4319;
wire n_5474;
wire n_18463;
wire n_8872;
wire n_644;
wire n_21923;
wire n_8752;
wire n_18214;
wire n_2004;
wire n_6069;
wire n_10963;
wire n_10191;
wire n_13330;
wire n_16127;
wire n_4751;
wire n_13412;
wire n_1196;
wire n_12638;
wire n_19015;
wire n_13561;
wire n_13306;
wire n_16961;
wire n_4298;
wire n_16122;
wire n_9517;
wire n_1089;
wire n_6386;
wire n_9192;
wire n_14089;
wire n_10025;
wire n_5957;
wire n_15603;
wire n_12066;
wire n_3383;
wire n_14822;
wire n_5490;
wire n_8291;
wire n_2704;
wire n_15337;
wire n_10179;
wire n_14076;
wire n_7433;
wire n_16856;
wire n_11702;
wire n_533;
wire n_10466;
wire n_1251;
wire n_18888;
wire n_15782;
wire n_8145;
wire n_10268;
wire n_13560;
wire n_15392;
wire n_10679;
wire n_19860;
wire n_7798;
wire n_4871;
wire n_12416;
wire n_16284;
wire n_17699;
wire n_2617;
wire n_13436;
wire n_6033;
wire n_1859;
wire n_18161;
wire n_5557;
wire n_7397;
wire n_16860;
wire n_13920;
wire n_20368;
wire n_8069;
wire n_14571;
wire n_5711;
wire n_4138;
wire n_19065;
wire n_21875;
wire n_5396;
wire n_1528;
wire n_2520;
wire n_17503;
wire n_956;
wire n_14908;
wire n_15522;
wire n_15534;
wire n_8797;
wire n_2134;
wire n_4236;
wire n_18325;
wire n_15225;
wire n_15386;
wire n_20994;
wire n_18743;
wire n_18953;
wire n_4238;
wire n_15508;
wire n_11491;
wire n_6142;
wire n_7510;
wire n_1545;
wire n_21050;
wire n_1799;
wire n_10729;
wire n_17680;
wire n_20666;
wire n_4013;
wire n_9884;
wire n_12127;
wire n_9857;
wire n_11637;
wire n_7257;
wire n_20536;
wire n_4242;
wire n_13537;
wire n_16521;
wire n_13808;
wire n_150;
wire n_3036;
wire n_12868;
wire n_12642;
wire n_17073;
wire n_10110;
wire n_14531;
wire n_8215;
wire n_11184;
wire n_191;
wire n_19042;
wire n_4561;
wire n_20314;
wire n_19962;
wire n_8629;
wire n_18548;
wire n_14887;
wire n_14172;
wire n_15518;
wire n_5556;
wire n_16100;
wire n_3696;
wire n_14593;
wire n_13507;
wire n_18280;
wire n_21578;
wire n_12300;
wire n_257;
wire n_14934;
wire n_709;
wire n_18664;
wire n_14988;
wire n_17538;
wire n_9004;
wire n_12832;
wire n_13839;
wire n_7865;
wire n_2652;
wire n_19909;
wire n_2635;
wire n_19846;
wire n_15746;
wire n_19921;
wire n_12290;
wire n_976;
wire n_20194;
wire n_20779;
wire n_6912;
wire n_10496;
wire n_11464;
wire n_14763;
wire n_11648;
wire n_8250;
wire n_18283;
wire n_10994;
wire n_11576;
wire n_1328;
wire n_2141;
wire n_13950;
wire n_6061;
wire n_4369;
wire n_14025;
wire n_12969;
wire n_8408;
wire n_10120;
wire n_15499;
wire n_11251;
wire n_1598;
wire n_16159;
wire n_3101;
wire n_6009;
wire n_12264;
wire n_11641;
wire n_5278;
wire n_8818;
wire n_17372;
wire n_7518;
wire n_12352;
wire n_580;
wire n_2693;
wire n_19238;
wire n_13619;
wire n_5675;
wire n_4135;
wire n_8275;
wire n_1218;
wire n_9327;
wire n_5771;
wire n_1547;
wire n_11555;
wire n_1755;
wire n_19345;
wire n_415;
wire n_485;
wire n_10611;
wire n_21480;
wire n_12368;
wire n_14038;
wire n_7705;
wire n_15259;
wire n_8590;
wire n_3291;
wire n_12538;
wire n_21203;
wire n_16537;
wire n_3405;
wire n_4745;
wire n_6155;
wire n_6738;
wire n_7854;
wire n_7707;
wire n_20636;
wire n_4629;
wire n_213;
wire n_8151;
wire n_6350;
wire n_18494;
wire n_9802;
wire n_8599;
wire n_4226;
wire n_4741;
wire n_1471;
wire n_11567;
wire n_1750;
wire n_19483;
wire n_4376;
wire n_5705;
wire n_12350;
wire n_10798;
wire n_20235;
wire n_571;
wire n_4552;
wire n_12891;
wire n_2713;
wire n_5196;
wire n_16298;
wire n_19007;
wire n_16057;
wire n_11779;
wire n_10166;
wire n_2951;
wire n_11684;
wire n_15843;
wire n_5126;
wire n_2214;
wire n_9842;
wire n_3427;
wire n_2055;
wire n_14893;
wire n_4042;
wire n_9524;
wire n_11129;
wire n_4385;
wire n_20177;
wire n_15079;
wire n_10848;
wire n_9122;
wire n_8743;
wire n_6603;
wire n_16136;
wire n_17590;
wire n_3359;
wire n_8473;
wire n_21221;
wire n_10342;
wire n_6245;
wire n_2865;
wire n_10439;
wire n_14284;
wire n_6703;
wire n_4717;
wire n_5604;
wire n_9676;
wire n_3789;
wire n_3598;
wire n_7714;
wire n_12759;
wire n_8535;
wire n_18832;
wire n_7011;
wire n_2139;
wire n_18555;
wire n_7621;
wire n_8068;
wire n_10565;
wire n_12935;
wire n_11058;
wire n_17270;
wire n_16955;
wire n_5114;
wire n_21514;
wire n_7028;
wire n_3433;
wire n_14437;
wire n_1072;
wire n_2305;
wire n_5699;
wire n_7525;
wire n_2450;
wire n_20023;
wire n_3447;
wire n_5810;
wire n_18635;
wire n_18852;
wire n_16077;
wire n_17715;
wire n_20740;
wire n_16672;
wire n_5762;
wire n_16705;
wire n_13713;
wire n_18715;
wire n_10686;
wire n_15975;
wire n_2271;
wire n_8327;
wire n_18969;
wire n_20191;
wire n_5408;
wire n_15810;
wire n_12374;
wire n_16099;
wire n_14266;
wire n_18784;
wire n_15440;
wire n_5366;
wire n_10132;
wire n_9872;
wire n_1847;
wire n_15354;
wire n_2767;
wire n_3116;
wire n_18020;
wire n_1884;
wire n_409;
wire n_18248;
wire n_11585;
wire n_9150;
wire n_2553;
wire n_17674;
wire n_3706;
wire n_16717;
wire n_21123;
wire n_18344;
wire n_300;
wire n_9984;
wire n_5451;
wire n_2626;
wire n_3441;
wire n_13855;
wire n_12179;
wire n_21342;
wire n_5086;
wire n_9814;
wire n_15513;
wire n_14689;
wire n_21739;
wire n_19930;
wire n_10211;
wire n_15335;
wire n_21088;
wire n_9461;
wire n_1997;
wire n_8997;
wire n_1477;
wire n_3142;
wire n_4623;
wire n_20029;
wire n_15838;
wire n_2690;
wire n_4410;
wire n_12952;
wire n_18968;
wire n_6803;
wire n_10446;
wire n_11735;
wire n_784;
wire n_6340;
wire n_8109;
wire n_1244;
wire n_17505;
wire n_19443;
wire n_7995;
wire n_11405;
wire n_6048;
wire n_1788;
wire n_14733;
wire n_16994;
wire n_12103;
wire n_9403;
wire n_5632;
wire n_865;
wire n_16268;
wire n_776;
wire n_2022;
wire n_3814;
wire n_19317;
wire n_4911;
wire n_14243;
wire n_4340;
wire n_9731;
wire n_5660;
wire n_21662;
wire n_13677;
wire n_4645;
wire n_7557;
wire n_21536;
wire n_20222;
wire n_18300;
wire n_6463;
wire n_20175;
wire n_16836;
wire n_21476;
wire n_1767;
wire n_9699;
wire n_6372;
wire n_9305;
wire n_12003;
wire n_19613;
wire n_20711;
wire n_11556;
wire n_13480;
wire n_17541;
wire n_18582;
wire n_3765;
wire n_15449;
wire n_18203;
wire n_9534;
wire n_18021;
wire n_1010;
wire n_1231;
wire n_5818;
wire n_6394;
wire n_9546;
wire n_3471;
wire n_7590;
wire n_15804;
wire n_2046;
wire n_11328;
wire n_16756;
wire n_21133;
wire n_21417;
wire n_3564;
wire n_14214;
wire n_16472;
wire n_11525;
wire n_9066;
wire n_10800;
wire n_3457;
wire n_9185;
wire n_1678;
wire n_17768;
wire n_9318;
wire n_4821;
wire n_8631;
wire n_18407;
wire n_5445;
wire n_16550;
wire n_21650;
wire n_15396;
wire n_15422;
wire n_7225;
wire n_11820;
wire n_14863;
wire n_10314;
wire n_3648;
wire n_12296;
wire n_9339;
wire n_5332;
wire n_13038;
wire n_456;
wire n_10006;
wire n_3031;
wire n_18196;
wire n_11441;
wire n_7432;
wire n_11242;
wire n_12804;
wire n_11471;
wire n_3385;
wire n_10346;
wire n_18917;
wire n_10539;
wire n_6321;
wire n_2768;
wire n_17948;
wire n_4826;
wire n_14479;
wire n_20306;
wire n_21733;
wire n_514;
wire n_1079;
wire n_7761;
wire n_7197;
wire n_20702;
wire n_16585;
wire n_15560;
wire n_12106;
wire n_1593;
wire n_17192;
wire n_21426;
wire n_9097;
wire n_12895;
wire n_11432;
wire n_4578;
wire n_19959;
wire n_14676;
wire n_7619;
wire n_12125;
wire n_2847;
wire n_1148;
wire n_750;
wire n_2790;
wire n_17113;
wire n_11164;
wire n_11527;
wire n_18277;
wire n_2359;
wire n_3674;
wire n_8083;
wire n_18662;
wire n_3098;
wire n_18292;
wire n_7403;
wire n_19056;
wire n_10145;
wire n_5569;
wire n_15631;
wire n_19101;
wire n_21705;
wire n_5439;
wire n_21939;
wire n_4147;
wire n_20500;
wire n_6481;
wire n_9810;
wire n_21125;
wire n_1309;
wire n_12047;
wire n_6534;
wire n_13289;
wire n_4974;
wire n_18561;
wire n_14224;
wire n_1800;
wire n_14015;
wire n_4932;
wire n_1421;
wire n_6181;
wire n_1177;
wire n_11642;
wire n_17176;
wire n_14566;
wire n_16796;
wire n_13549;
wire n_5119;
wire n_14874;
wire n_9264;
wire n_21379;
wire n_17050;
wire n_829;
wire n_3354;
wire n_2724;
wire n_14155;
wire n_16226;
wire n_16909;
wire n_17047;
wire n_4285;
wire n_20195;
wire n_9550;
wire n_6282;
wire n_21674;
wire n_9929;
wire n_274;
wire n_15877;
wire n_21494;
wire n_20760;
wire n_11092;
wire n_1332;
wire n_18392;
wire n_2090;
wire n_16195;
wire n_20416;
wire n_3153;
wire n_15362;
wire n_12770;
wire n_5932;
wire n_6234;
wire n_15226;
wire n_2400;
wire n_4633;
wire n_14518;
wire n_3838;
wire n_10857;
wire n_15279;
wire n_15750;
wire n_5092;
wire n_10708;
wire n_21313;
wire n_20618;
wire n_11045;
wire n_19510;
wire n_8619;
wire n_9559;
wire n_11993;
wire n_15448;
wire n_9806;
wire n_4662;
wire n_18823;
wire n_4882;
wire n_15031;
wire n_7582;
wire n_13997;
wire n_987;
wire n_4868;
wire n_8923;
wire n_14302;
wire n_21115;
wire n_11408;
wire n_2452;
wire n_17223;
wire n_14829;
wire n_8876;
wire n_3925;
wire n_11670;
wire n_10067;
wire n_19516;
wire n_19484;
wire n_4059;
wire n_18653;
wire n_11604;
wire n_16575;
wire n_14433;
wire n_19099;
wire n_6682;
wire n_5054;
wire n_2467;
wire n_6539;
wire n_17844;
wire n_18294;
wire n_7179;
wire n_5399;
wire n_10222;
wire n_11293;
wire n_4650;
wire n_12072;
wire n_21430;
wire n_1435;
wire n_19059;
wire n_13941;
wire n_4339;
wire n_6595;
wire n_1645;
wire n_14986;
wire n_7738;
wire n_9223;
wire n_2658;
wire n_10647;
wire n_9499;
wire n_21974;
wire n_16788;
wire n_13036;
wire n_5391;
wire n_20527;
wire n_8073;
wire n_4541;
wire n_13225;
wire n_6385;
wire n_3388;
wire n_13587;
wire n_5523;
wire n_16205;
wire n_21668;
wire n_21851;
wire n_4796;
wire n_18519;
wire n_9120;
wire n_14917;
wire n_10405;
wire n_20331;
wire n_12726;
wire n_12833;
wire n_14206;
wire n_2694;
wire n_15787;
wire n_9386;
wire n_16087;
wire n_6346;
wire n_4775;
wire n_9779;
wire n_18891;
wire n_7587;
wire n_4381;
wire n_3886;
wire n_16882;
wire n_4455;
wire n_14381;
wire n_2328;
wire n_19322;
wire n_7760;
wire n_10588;
wire n_15699;
wire n_9444;
wire n_19282;
wire n_20597;
wire n_7057;
wire n_15840;
wire n_8031;
wire n_14193;
wire n_4554;
wire n_5595;
wire n_6815;
wire n_1299;
wire n_9317;
wire n_14968;
wire n_20737;
wire n_17529;
wire n_21118;
wire n_14262;
wire n_14723;
wire n_8509;
wire n_16773;
wire n_13659;
wire n_21726;
wire n_11564;
wire n_10641;
wire n_11719;
wire n_19678;
wire n_15795;
wire n_9275;
wire n_19356;
wire n_21071;
wire n_13248;
wire n_5372;
wire n_17359;
wire n_2402;
wire n_4301;
wire n_11754;
wire n_1050;
wire n_14369;
wire n_17991;
wire n_17066;
wire n_11075;
wire n_17370;
wire n_3777;
wire n_10722;
wire n_14422;
wire n_13005;
wire n_20882;
wire n_8429;
wire n_21992;
wire n_15033;
wire n_2701;
wire n_5929;
wire n_1631;
wire n_3105;
wire n_13972;
wire n_7388;
wire n_16225;
wire n_7694;
wire n_4286;
wire n_21395;
wire n_16532;
wire n_5102;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_21539;
wire n_2816;
wire n_16571;
wire n_7982;
wire n_11384;
wire n_18527;
wire n_19907;
wire n_10763;
wire n_21636;
wire n_18595;
wire n_8773;
wire n_18296;
wire n_8225;
wire n_18047;
wire n_6867;
wire n_17646;
wire n_9556;
wire n_1143;
wire n_6230;
wire n_12810;
wire n_9259;
wire n_9995;
wire n_12820;
wire n_8080;
wire n_14927;
wire n_18372;
wire n_19434;
wire n_14236;
wire n_17315;
wire n_15606;
wire n_15051;
wire n_21024;
wire n_17075;
wire n_1992;
wire n_4402;
wire n_15660;
wire n_4239;
wire n_6854;
wire n_21630;
wire n_17282;
wire n_2169;
wire n_17240;
wire n_19240;
wire n_18938;
wire n_6784;
wire n_6168;
wire n_16781;
wire n_8431;
wire n_8453;
wire n_3316;
wire n_18495;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_8634;
wire n_3603;
wire n_2192;
wire n_3633;
wire n_9713;
wire n_16111;
wire n_10104;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_6799;
wire n_10115;
wire n_13654;
wire n_19643;
wire n_8015;
wire n_10397;
wire n_10398;
wire n_17480;
wire n_18733;
wire n_21047;
wire n_21264;
wire n_6149;
wire n_1671;
wire n_19729;
wire n_10065;
wire n_11156;
wire n_11598;
wire n_13977;
wire n_5808;
wire n_21400;
wire n_1062;
wire n_11176;
wire n_12687;
wire n_12260;
wire n_19217;
wire n_5353;
wire n_3708;
wire n_8074;
wire n_4437;
wire n_16819;
wire n_3861;
wire n_7042;
wire n_8039;
wire n_5382;
wire n_1188;
wire n_18547;
wire n_17428;
wire n_12474;
wire n_9241;
wire n_21165;
wire n_10422;
wire n_10736;
wire n_19587;
wire n_6134;
wire n_8537;
wire n_4513;
wire n_3233;
wire n_20423;
wire n_9600;
wire n_11095;
wire n_2352;
wire n_4040;
wire n_9927;
wire n_17145;
wire n_10046;
wire n_15157;
wire n_20724;
wire n_16525;
wire n_19656;
wire n_3123;
wire n_18157;
wire n_20950;
wire n_8437;
wire n_7447;
wire n_13956;
wire n_21282;
wire n_14617;
wire n_5233;
wire n_13819;
wire n_3520;
wire n_11602;
wire n_2492;
wire n_21856;
wire n_12934;
wire n_6493;
wire n_14843;
wire n_13566;
wire n_14315;
wire n_18167;
wire n_4904;
wire n_8980;
wire n_1419;
wire n_7629;
wire n_18880;
wire n_7104;
wire n_9844;
wire n_15376;
wire n_15467;
wire n_21406;
wire n_12457;
wire n_12743;
wire n_20182;
wire n_4290;
wire n_5247;
wire n_8030;
wire n_9663;
wire n_10168;
wire n_18267;
wire n_306;
wire n_6544;
wire n_20095;
wire n_14424;
wire n_13077;
wire n_21815;
wire n_1597;
wire n_9628;
wire n_1659;
wire n_20524;
wire n_14560;
wire n_14273;
wire n_13891;
wire n_14090;
wire n_5380;
wire n_18382;
wire n_5924;
wire n_3182;
wire n_2564;
wire n_876;
wire n_19413;
wire n_11246;
wire n_17545;
wire n_21418;
wire n_16830;
wire n_4656;
wire n_12766;
wire n_3896;
wire n_3958;
wire n_6390;
wire n_21444;
wire n_11970;
wire n_13466;
wire n_20513;
wire n_1116;
wire n_7971;
wire n_3174;
wire n_982;
wire n_18033;
wire n_10927;
wire n_10704;
wire n_3398;
wire n_5388;
wire n_2640;
wire n_13231;
wire n_6279;
wire n_14461;
wire n_21001;
wire n_8751;
wire n_18729;
wire n_679;
wire n_12875;
wire n_11085;
wire n_12808;
wire n_14897;
wire n_1427;
wire n_14041;
wire n_14817;
wire n_15675;
wire n_21427;
wire n_10011;
wire n_6675;
wire n_4323;
wire n_2212;
wire n_6476;
wire n_14397;
wire n_19615;
wire n_10982;
wire n_5539;
wire n_6268;
wire n_21979;
wire n_17660;
wire n_6878;
wire n_6286;
wire n_9088;
wire n_3308;
wire n_5036;
wire n_18703;
wire n_12910;
wire n_4772;
wire n_19505;
wire n_20573;
wire n_5893;
wire n_17794;
wire n_20425;
wire n_5273;
wire n_10262;
wire n_8360;
wire n_8036;
wire n_16121;
wire n_11423;
wire n_17616;
wire n_7853;
wire n_17818;
wire n_3757;
wire n_11370;
wire n_1782;
wire n_2245;
wire n_12394;
wire n_9411;
wire n_1524;
wire n_1485;
wire n_9543;
wire n_416;
wire n_3635;
wire n_17742;
wire n_5005;
wire n_13174;
wire n_21484;
wire n_1570;
wire n_3882;
wire n_16640;
wire n_1170;
wire n_305;
wire n_2213;
wire n_6425;
wire n_14201;
wire n_12253;
wire n_2095;
wire n_3121;
wire n_18429;
wire n_20585;
wire n_14296;
wire n_17134;
wire n_13579;
wire n_2527;
wire n_9404;
wire n_16331;
wire n_5534;
wire n_1461;
wire n_9678;
wire n_21919;
wire n_15414;
wire n_11071;
wire n_11979;
wire n_18895;
wire n_8626;
wire n_6955;
wire n_9481;
wire n_5174;
wire n_4952;
wire n_15872;
wire n_19450;
wire n_17897;
wire n_3005;
wire n_1235;
wire n_9672;
wire n_14009;
wire n_3129;
wire n_7237;
wire n_1783;
wire n_8935;
wire n_20213;
wire n_12590;
wire n_2375;
wire n_6388;
wire n_17472;
wire n_10240;
wire n_5904;
wire n_13465;
wire n_14026;
wire n_8009;
wire n_11329;
wire n_2344;
wire n_20472;
wire n_5620;
wire n_12034;
wire n_1295;
wire n_5750;
wire n_21167;
wire n_3219;
wire n_9042;
wire n_9506;
wire n_1762;
wire n_15655;
wire n_8008;
wire n_19795;
wire n_3023;
wire n_6664;
wire n_15695;
wire n_5815;
wire n_17195;
wire n_18842;
wire n_13926;
wire n_14163;
wire n_612;
wire n_4737;
wire n_6729;
wire n_17016;
wire n_9862;
wire n_15407;
wire n_5949;
wire n_16302;
wire n_10469;
wire n_7483;
wire n_20001;
wire n_6608;
wire n_14145;
wire n_19221;
wire n_9619;
wire n_1952;
wire n_13902;
wire n_11088;
wire n_9508;
wire n_7668;
wire n_17839;
wire n_16567;
wire n_2560;
wire n_4522;
wire n_13504;
wire n_5955;
wire n_7476;
wire n_19925;
wire n_21321;
wire n_18809;
wire n_13491;
wire n_14135;
wire n_6843;
wire n_3140;
wire n_16322;
wire n_3724;
wire n_8118;
wire n_14182;
wire n_298;
wire n_21180;
wire n_12882;
wire n_11449;
wire n_16445;
wire n_4675;
wire n_5340;
wire n_7100;
wire n_19424;
wire n_5783;
wire n_11123;
wire n_3084;
wire n_1727;
wire n_17322;
wire n_5549;
wire n_9935;
wire n_20940;
wire n_16410;
wire n_8376;
wire n_9827;
wire n_4889;
wire n_5442;
wire n_5739;
wire n_20181;
wire n_13161;
wire n_3184;
wire n_16167;
wire n_5385;
wire n_8799;
wire n_4558;
wire n_15607;
wire n_15232;
wire n_15512;
wire n_6086;
wire n_17645;
wire n_6650;
wire n_158;
wire n_4768;
wire n_12941;
wire n_21758;
wire n_14476;
wire n_10088;
wire n_14208;
wire n_5845;
wire n_20296;
wire n_20681;
wire n_10247;
wire n_18526;
wire n_9236;
wire n_400;
wire n_6060;
wire n_12537;
wire n_2194;
wire n_848;
wire n_17421;
wire n_16633;
wire n_5537;
wire n_2680;
wire n_13835;
wire n_6059;
wire n_17220;
wire n_7520;
wire n_3122;
wire n_4808;
wire n_16686;
wire n_6103;
wire n_3265;
wire n_15328;
wire n_10986;
wire n_19378;
wire n_2957;
wire n_9127;
wire n_12521;
wire n_18935;
wire n_20202;
wire n_5855;
wire n_10069;
wire n_15300;
wire n_19719;
wire n_12866;
wire n_1250;
wire n_3309;
wire n_12170;
wire n_19330;
wire n_8886;
wire n_10844;
wire n_772;
wire n_16613;
wire n_3357;
wire n_10330;
wire n_15571;
wire n_7163;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_18623;
wire n_11765;
wire n_3754;
wire n_16372;
wire n_14648;
wire n_12440;
wire n_21600;
wire n_4287;
wire n_10584;
wire n_16188;
wire n_21034;
wire n_16118;
wire n_4516;
wire n_18617;
wire n_12834;
wire n_14791;
wire n_2809;
wire n_2050;
wire n_8720;
wire n_1676;
wire n_1113;
wire n_21490;
wire n_18146;
wire n_11278;
wire n_5172;
wire n_4449;
wire n_13497;
wire n_8219;
wire n_502;
wire n_14941;
wire n_16986;
wire n_15725;
wire n_6377;
wire n_466;
wire n_19611;
wire n_21886;
wire n_20615;
wire n_5414;
wire n_1245;
wire n_20993;
wire n_11713;
wire n_1321;
wire n_15691;
wire n_12214;
wire n_13282;
wire n_6348;
wire n_7713;
wire n_15545;
wire n_20028;
wire n_2135;
wire n_17167;
wire n_3493;
wire n_10124;
wire n_18053;
wire n_14816;
wire n_12320;
wire n_2734;
wire n_9792;
wire n_6136;
wire n_19257;
wire n_8066;
wire n_14459;
wire n_14970;
wire n_21099;
wire n_14063;
wire n_14976;
wire n_20898;
wire n_13527;
wire n_9712;
wire n_7021;
wire n_16147;
wire n_1606;
wire n_17684;
wire n_17431;
wire n_2485;
wire n_15905;
wire n_17579;
wire n_10144;
wire n_8402;
wire n_7130;
wire n_20154;
wire n_11714;
wire n_4032;
wire n_21530;
wire n_13794;
wire n_14948;
wire n_1583;
wire n_16436;
wire n_20258;
wire n_11300;
wire n_1493;
wire n_11338;
wire n_6642;
wire n_5522;
wire n_11930;
wire n_10525;
wire n_2708;
wire n_18944;
wire n_20721;
wire n_11334;
wire n_2225;
wire n_18744;
wire n_17494;
wire n_7546;
wire n_5934;
wire n_8418;
wire n_18291;
wire n_20447;
wire n_18278;
wire n_2938;
wire n_9111;
wire n_12677;
wire n_11482;
wire n_17639;
wire n_6001;
wire n_6007;
wire n_6606;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_14327;
wire n_13901;
wire n_7078;
wire n_3463;
wire n_18937;
wire n_7107;
wire n_16360;
wire n_20301;
wire n_21878;
wire n_16758;
wire n_10325;
wire n_2728;
wire n_14786;

INVx2_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_39),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_114),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_84),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_14),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_20),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_45),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_74),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_124),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_41),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_19),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_80),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_78),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_6),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_112),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_52),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_72),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_0),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_75),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_118),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_54),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_70),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_15),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_85),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_119),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_89),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_90),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_71),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_13),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_53),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_27),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_28),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_40),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_63),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_64),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_4),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_103),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_37),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_60),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_129),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_1),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_105),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_69),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_32),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_1),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_76),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_35),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_108),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_16),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_3),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_111),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_62),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_127),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_25),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_23),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_30),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_51),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_68),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_95),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_61),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_122),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_56),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_38),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_48),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_21),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_130),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_98),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_26),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_46),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_115),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_9),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_47),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_5),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_12),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_96),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_91),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_43),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_94),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_106),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_82),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_83),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_49),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_81),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_44),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_8),
.Y(n_247)
);

BUFx10_ASAP7_75t_L g248 ( 
.A(n_79),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_17),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_31),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_113),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_33),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_117),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_58),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_24),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_7),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_92),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_99),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_22),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_134),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_10),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_0),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_110),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_67),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_34),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_29),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_36),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_57),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_202),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_140),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_141),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_202),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_144),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_169),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_197),
.B(n_11),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_137),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_143),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_145),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_148),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_146),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_150),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_151),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_152),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_155),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_165),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_157),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_167),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_174),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_158),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_159),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_175),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_257),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_179),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_181),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_185),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_189),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g304 ( 
.A(n_194),
.B(n_42),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_195),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_160),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_201),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_231),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_206),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_171),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_271),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_274),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_275),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_297),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

BUFx6f_ASAP7_75t_SL g323 ( 
.A(n_273),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_309),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_282),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_310),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_298),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_307),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_276),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_311),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_283),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_304),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_291),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_294),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_295),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_296),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_306),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_286),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_270),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_312),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_186),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g363 ( 
.A1(n_349),
.A2(n_223),
.B(n_253),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

BUFx12f_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

AND2x2_ASAP7_75t_SL g370 ( 
.A(n_344),
.B(n_136),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

NOR2x1_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_147),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g373 ( 
.A(n_313),
.B(n_138),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

AOI22x1_ASAP7_75t_SL g376 ( 
.A1(n_360),
.A2(n_230),
.B1(n_269),
.B2(n_184),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_341),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_327),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

AOI22x1_ASAP7_75t_SL g382 ( 
.A1(n_314),
.A2(n_163),
.B1(n_154),
.B2(n_164),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_329),
.B(n_180),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_237),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_317),
.A2(n_217),
.B1(n_211),
.B2(n_221),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_139),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_334),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_335),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_338),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_339),
.B(n_153),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_315),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_356),
.A2(n_210),
.B1(n_226),
.B2(n_261),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_357),
.B(n_248),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_340),
.B(n_173),
.Y(n_397)
);

BUFx12f_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_161),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_345),
.B(n_259),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_343),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_354),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_353),
.A2(n_256),
.B(n_255),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_162),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_320),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_320),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_333),
.B(n_207),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_320),
.Y(n_416)
);

INVx6_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_320),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_320),
.Y(n_420)
);

INVx6_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_344),
.B(n_248),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_313),
.Y(n_423)
);

CKINVDCx11_ASAP7_75t_R g424 ( 
.A(n_360),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_R g425 ( 
.A1(n_344),
.A2(n_218),
.B1(n_265),
.B2(n_212),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_349),
.B(n_166),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_349),
.B(n_268),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_341),
.A2(n_267),
.B1(n_266),
.B2(n_258),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_320),
.Y(n_429)
);

AND2x4_ASAP7_75t_SL g430 ( 
.A(n_344),
.B(n_264),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_333),
.B(n_215),
.Y(n_431)
);

BUFx12f_ASAP7_75t_L g432 ( 
.A(n_342),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_349),
.B(n_213),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_320),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_320),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_322),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_333),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_320),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_320),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_341),
.A2(n_208),
.B1(n_241),
.B2(n_235),
.Y(n_440)
);

CKINVDCx11_ASAP7_75t_R g441 ( 
.A(n_360),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_333),
.B(n_216),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_320),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_349),
.B(n_209),
.Y(n_444)
);

OA21x2_ASAP7_75t_L g445 ( 
.A1(n_349),
.A2(n_191),
.B(n_214),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_320),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_342),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_320),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_320),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_322),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_333),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_320),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_320),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_320),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_320),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_349),
.A2(n_177),
.B(n_156),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_320),
.Y(n_458)
);

BUFx8_ASAP7_75t_L g459 ( 
.A(n_323),
.Y(n_459)
);

INVxp33_ASAP7_75t_SL g460 ( 
.A(n_344),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_350),
.A2(n_222),
.B1(n_251),
.B2(n_250),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_320),
.Y(n_462)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_313),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_322),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_322),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_320),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_333),
.B(n_247),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_344),
.Y(n_468)
);

CKINVDCx6p67_ASAP7_75t_R g469 ( 
.A(n_323),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_320),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_320),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_320),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_349),
.B(n_204),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_349),
.B(n_205),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_320),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_333),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_333),
.B(n_246),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_320),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_344),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_344),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_322),
.Y(n_481)
);

AND3x1_ASAP7_75t_L g482 ( 
.A(n_347),
.B(n_244),
.C(n_260),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_344),
.B(n_264),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_320),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_342),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_320),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_333),
.B(n_240),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_320),
.Y(n_488)
);

NOR2x1_ASAP7_75t_L g489 ( 
.A(n_350),
.B(n_142),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_322),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_320),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_349),
.B(n_203),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_322),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_409),
.A2(n_149),
.B(n_238),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_404),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_361),
.B(n_242),
.Y(n_496)
);

AND2x2_ASAP7_75t_SL g497 ( 
.A(n_370),
.B(n_245),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_367),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_363),
.A2(n_227),
.B(n_236),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_369),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_480),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_381),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_412),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_412),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_389),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_365),
.B(n_196),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_390),
.Y(n_508)
);

NAND2x1_ASAP7_75t_L g509 ( 
.A(n_401),
.B(n_262),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_391),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_392),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_437),
.B(n_198),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_422),
.B(n_193),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_413),
.B(n_199),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_436),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_418),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_394),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_418),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_414),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_402),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_403),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_451),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_464),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_465),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_481),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_490),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_493),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_372),
.B(n_262),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_434),
.Y(n_531)
);

AND2x2_ASAP7_75t_SL g532 ( 
.A(n_396),
.B(n_262),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_446),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_399),
.B(n_192),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_452),
.B(n_190),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g536 ( 
.A1(n_457),
.A2(n_254),
.B(n_252),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_449),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_383),
.B(n_188),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_435),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_476),
.B(n_187),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_479),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_453),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_375),
.B(n_380),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_483),
.B(n_234),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_489),
.A2(n_232),
.B(n_219),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_410),
.B(n_426),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_462),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_375),
.B(n_183),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_364),
.B(n_233),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_435),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_471),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_470),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_416),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_472),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_475),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_377),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_486),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_368),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_374),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_419),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_380),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_SL g567 ( 
.A(n_385),
.B(n_395),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_386),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_362),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_429),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_373),
.A2(n_182),
.B1(n_229),
.B2(n_168),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_427),
.B(n_176),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_466),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_478),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_386),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_379),
.A2(n_178),
.B1(n_228),
.B2(n_170),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_484),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_491),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_371),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_433),
.B(n_220),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_444),
.B(n_172),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_473),
.B(n_224),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_400),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_471),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_439),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_387),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_428),
.B(n_225),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_406),
.B(n_219),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_443),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_447),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_458),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_488),
.Y(n_593)
);

OA21x2_ASAP7_75t_L g594 ( 
.A1(n_474),
.A2(n_232),
.B(n_59),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_445),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_407),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_388),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_440),
.B(n_232),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_393),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_407),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_492),
.B(n_232),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_397),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_423),
.B(n_93),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_415),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_417),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_431),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_421),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_384),
.B(n_232),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_442),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_467),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_477),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_430),
.B(n_405),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_R g613 ( 
.A(n_448),
.B(n_485),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_378),
.B(n_487),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_482),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_425),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_461),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_423),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_408),
.B(n_463),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_463),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_424),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_366),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_398),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_469),
.B(n_432),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_376),
.Y(n_625)
);

OA21x2_ASAP7_75t_L g626 ( 
.A1(n_382),
.A2(n_441),
.B(n_459),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_404),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_437),
.B(n_452),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_367),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_367),
.Y(n_630)
);

AND2x6_ASAP7_75t_L g631 ( 
.A(n_372),
.B(n_489),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_361),
.B(n_365),
.Y(n_632)
);

BUFx8_ASAP7_75t_L g633 ( 
.A(n_468),
.Y(n_633)
);

CKINVDCx8_ASAP7_75t_R g634 ( 
.A(n_423),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_367),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_468),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_361),
.B(n_312),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_468),
.B(n_344),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_404),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_404),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_468),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_414),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_412),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_404),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_367),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_414),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_404),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_372),
.B(n_489),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_367),
.Y(n_649)
);

OA21x2_ASAP7_75t_L g650 ( 
.A1(n_409),
.A2(n_457),
.B(n_363),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_468),
.B(n_344),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_367),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_468),
.B(n_344),
.Y(n_653)
);

OA21x2_ASAP7_75t_L g654 ( 
.A1(n_409),
.A2(n_457),
.B(n_363),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_404),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_448),
.B(n_360),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_437),
.B(n_452),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_367),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_468),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_367),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_361),
.B(n_312),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_367),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_367),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_468),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_367),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_367),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_424),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_404),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_367),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_468),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_367),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_367),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_367),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_367),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_370),
.B(n_361),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_437),
.B(n_452),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_367),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_412),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_367),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_404),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_412),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_404),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_367),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_417),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_SL g685 ( 
.A1(n_395),
.A2(n_385),
.B1(n_460),
.B2(n_370),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_367),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_367),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_367),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_414),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_367),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_468),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_367),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_414),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_468),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_404),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_404),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_404),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_367),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_412),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_412),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_404),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_404),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_361),
.B(n_365),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_414),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_404),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_367),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_404),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_412),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_367),
.Y(n_709)
);

OA21x2_ASAP7_75t_L g710 ( 
.A1(n_409),
.A2(n_457),
.B(n_363),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_367),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_361),
.B(n_365),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_367),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_437),
.B(n_452),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_468),
.B(n_344),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_448),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_367),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_363),
.A2(n_457),
.B(n_409),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_367),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_404),
.Y(n_720)
);

NAND2x1p5_ASAP7_75t_L g721 ( 
.A(n_364),
.B(n_407),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_370),
.A2(n_361),
.B1(n_372),
.B2(n_379),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_404),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_367),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_367),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_361),
.B(n_312),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_367),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_404),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_367),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_437),
.B(n_452),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_468),
.B(n_344),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_367),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_367),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_361),
.B(n_365),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_437),
.B(n_452),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_468),
.B(n_344),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_367),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_468),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_404),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_367),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_361),
.B(n_365),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_468),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_367),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_468),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_367),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_468),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_370),
.B(n_361),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_361),
.B(n_365),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_367),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_370),
.B(n_361),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_370),
.B(n_361),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_437),
.B(n_452),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_367),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_404),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_404),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_412),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_367),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_404),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_448),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_367),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_404),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_361),
.B(n_312),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_395),
.A2(n_385),
.B1(n_460),
.B2(n_370),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_367),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_367),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_437),
.B(n_452),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_404),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_367),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_404),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_363),
.A2(n_457),
.B(n_409),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_404),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_404),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_404),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_370),
.B(n_361),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_367),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_367),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_414),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_367),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_367),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_417),
.Y(n_780)
);

AND3x1_ASAP7_75t_L g781 ( 
.A(n_396),
.B(n_483),
.C(n_422),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_414),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_370),
.B(n_361),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_468),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_367),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_367),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_367),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_404),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_370),
.B(n_361),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_412),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_414),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_404),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_468),
.B(n_344),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_414),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_361),
.B(n_365),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_372),
.B(n_489),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_370),
.B(n_361),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_367),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_412),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_367),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_367),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_404),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_361),
.B(n_365),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_367),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_404),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_468),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_367),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_367),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_367),
.Y(n_809)
);

BUFx6f_ASAP7_75t_L g810 ( 
.A(n_412),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_372),
.B(n_489),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_523),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_527),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_637),
.B(n_726),
.C(n_661),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_497),
.B(n_722),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_684),
.B(n_780),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_632),
.B(n_703),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_712),
.B(n_734),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_741),
.B(n_748),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_499),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_501),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_503),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_795),
.B(n_803),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_675),
.B(n_747),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_506),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_750),
.B(n_751),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_641),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_774),
.A2(n_783),
.B1(n_797),
.B2(n_789),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_508),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_510),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_596),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_550),
.B(n_597),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_511),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_513),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_516),
.Y(n_835)
);

BUFx10_ASAP7_75t_L g836 ( 
.A(n_618),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_762),
.B(n_715),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_599),
.B(n_602),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_607),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_496),
.B(n_573),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_524),
.Y(n_841)
);

NOR2x1p5_ASAP7_75t_L g842 ( 
.A(n_596),
.B(n_600),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_525),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_607),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_664),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_532),
.B(n_638),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_SL g847 ( 
.A(n_716),
.B(n_759),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_600),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_526),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_631),
.B(n_648),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_504),
.Y(n_851)
);

AND2x6_ASAP7_75t_L g852 ( 
.A(n_617),
.B(n_615),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_534),
.B(n_528),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_629),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_605),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_630),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_567),
.B(n_616),
.C(n_651),
.Y(n_857)
);

NAND2xp33_ASAP7_75t_SL g858 ( 
.A(n_613),
.B(n_685),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_635),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_504),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_645),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_731),
.B(n_653),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_649),
.B(n_652),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_658),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_660),
.B(n_662),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_663),
.B(n_665),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_736),
.B(n_793),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_666),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_631),
.B(n_648),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_669),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_738),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_671),
.B(n_672),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_673),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_542),
.B(n_636),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_744),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_674),
.B(n_677),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_659),
.Y(n_877)
);

BUFx6f_ASAP7_75t_SL g878 ( 
.A(n_618),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_561),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_679),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_505),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_683),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_686),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_620),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_687),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_688),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_690),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_781),
.B(n_514),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_692),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_698),
.B(n_706),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_601),
.A2(n_538),
.B(n_595),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_709),
.Y(n_892)
);

NAND3xp33_ASAP7_75t_L g893 ( 
.A(n_670),
.B(n_742),
.C(n_694),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_505),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_711),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_713),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_620),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_717),
.B(n_719),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_724),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_517),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_498),
.B(n_502),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_725),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_598),
.A2(n_729),
.B1(n_732),
.B2(n_727),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_733),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_737),
.Y(n_905)
);

OAI22xp33_ASAP7_75t_L g906 ( 
.A1(n_740),
.A2(n_745),
.B1(n_778),
.B2(n_743),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_749),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_517),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_519),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_753),
.B(n_757),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_547),
.B(n_614),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_760),
.B(n_764),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_765),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_768),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_775),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_691),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_746),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_519),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_776),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_779),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_603),
.B(n_612),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_785),
.Y(n_922)
);

OAI22xp33_ASAP7_75t_L g923 ( 
.A1(n_786),
.A2(n_798),
.B1(n_804),
.B2(n_787),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_SL g924 ( 
.A(n_763),
.B(n_572),
.C(n_625),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_800),
.B(n_801),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_807),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_784),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_808),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_628),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_809),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_796),
.A2(n_811),
.B1(n_648),
.B2(n_631),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_539),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_539),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_L g934 ( 
.A(n_577),
.B(n_806),
.C(n_555),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_554),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_SL g936 ( 
.A1(n_608),
.A2(n_546),
.B(n_515),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_721),
.B(n_566),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_530),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_606),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_531),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_533),
.Y(n_941)
);

BUFx8_ASAP7_75t_SL g942 ( 
.A(n_667),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_657),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_554),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_586),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_495),
.B(n_627),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_540),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_544),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_537),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_676),
.B(n_714),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_568),
.B(n_576),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_545),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_549),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_730),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_639),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_543),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_581),
.B(n_582),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_640),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_551),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_556),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_735),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_556),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_604),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_553),
.B(n_512),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_644),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_583),
.B(n_643),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_647),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_557),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_655),
.B(n_668),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_559),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_680),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_643),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_682),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_560),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_695),
.B(n_696),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_697),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_562),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_609),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_701),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_702),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_705),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_811),
.B(n_529),
.Y(n_982)
);

INVxp33_ASAP7_75t_L g983 ( 
.A(n_656),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_707),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_610),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_811),
.A2(n_529),
.B1(n_773),
.B2(n_767),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_720),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_529),
.B(n_723),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_728),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_739),
.B(n_754),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_755),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_678),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_758),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_611),
.Y(n_994)
);

AND2x2_ASAP7_75t_SL g995 ( 
.A(n_626),
.B(n_621),
.Y(n_995)
);

AND3x2_ASAP7_75t_L g996 ( 
.A(n_624),
.B(n_622),
.C(n_623),
.Y(n_996)
);

NAND2xp33_ASAP7_75t_L g997 ( 
.A(n_678),
.B(n_681),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_761),
.B(n_769),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_L g999 ( 
.A(n_681),
.B(n_699),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_771),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_772),
.B(n_788),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_699),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_792),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_802),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_805),
.Y(n_1005)
);

OAI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_518),
.A2(n_522),
.B1(n_521),
.B2(n_563),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_564),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_700),
.B(n_799),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_588),
.B(n_766),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_700),
.B(n_708),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_708),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_569),
.Y(n_1012)
);

NAND3xp33_ASAP7_75t_L g1013 ( 
.A(n_584),
.B(n_507),
.C(n_541),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_585),
.B(n_810),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_756),
.B(n_810),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_752),
.B(n_565),
.Y(n_1016)
);

NAND2xp33_ASAP7_75t_L g1017 ( 
.A(n_756),
.B(n_799),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_535),
.B(n_580),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_790),
.B(n_575),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_790),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_520),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_571),
.B(n_578),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_558),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_570),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_621),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_574),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_591),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_642),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_579),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_646),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_587),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_634),
.B(n_552),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_619),
.B(n_794),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_590),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_592),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_689),
.B(n_791),
.Y(n_1036)
);

NAND2xp33_ASAP7_75t_L g1037 ( 
.A(n_589),
.B(n_593),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_693),
.B(n_782),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_704),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_589),
.B(n_777),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_633),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_548),
.B(n_770),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_509),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_594),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_589),
.B(n_494),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_500),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_650),
.B(n_654),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_718),
.B(n_536),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_710),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_497),
.B(n_370),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_607),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_499),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_632),
.B(n_703),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_499),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_499),
.Y(n_1055)
);

OAI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_496),
.A2(n_722),
.B1(n_617),
.B2(n_550),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_632),
.B(n_703),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_497),
.B(n_370),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_607),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_498),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_499),
.Y(n_1061)
);

INVx5_ASAP7_75t_L g1062 ( 
.A(n_618),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_499),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_523),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_523),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_607),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_636),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_499),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_523),
.Y(n_1069)
);

HAxp5_ASAP7_75t_SL g1070 ( 
.A(n_616),
.B(n_722),
.CON(n_1070),
.SN(n_1070)
);

BUFx10_ASAP7_75t_L g1071 ( 
.A(n_618),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_523),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_638),
.B(n_344),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_684),
.B(n_780),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_638),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_596),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_632),
.B(n_703),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_632),
.B(n_703),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_497),
.B(n_370),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_499),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_637),
.B(n_726),
.C(n_661),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_523),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_523),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_499),
.Y(n_1084)
);

INVx4_ASAP7_75t_L g1085 ( 
.A(n_596),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_636),
.Y(n_1086)
);

INVxp67_ASAP7_75t_SL g1087 ( 
.A(n_504),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_499),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_523),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_499),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_523),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_L g1092 ( 
.A(n_631),
.B(n_811),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_523),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_523),
.Y(n_1094)
);

OR2x6_ASAP7_75t_L g1095 ( 
.A(n_596),
.B(n_600),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_607),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_499),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_523),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_497),
.B(n_370),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_504),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_607),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_523),
.Y(n_1102)
);

AND3x1_ASAP7_75t_L g1103 ( 
.A(n_616),
.B(n_396),
.C(n_615),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_523),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_632),
.B(n_703),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_632),
.B(n_703),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_607),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_497),
.B(n_370),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_715),
.B(n_731),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_499),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_632),
.B(n_703),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_523),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_499),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_SL g1114 ( 
.A(n_618),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_607),
.Y(n_1115)
);

AND2x6_ASAP7_75t_L g1116 ( 
.A(n_617),
.B(n_550),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_607),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_523),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_596),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_499),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_523),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_632),
.B(n_703),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_607),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_618),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_499),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_497),
.A2(n_617),
.B1(n_496),
.B2(n_598),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_523),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_496),
.A2(n_550),
.B(n_661),
.C(n_637),
.Y(n_1128)
);

INVx8_ASAP7_75t_L g1129 ( 
.A(n_596),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_596),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_638),
.Y(n_1131)
);

OAI22x1_ASAP7_75t_L g1132 ( 
.A1(n_616),
.A2(n_344),
.B1(n_480),
.B2(n_468),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_499),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_499),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_499),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_523),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_632),
.B(n_703),
.Y(n_1137)
);

INVx6_ASAP7_75t_L g1138 ( 
.A(n_596),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_632),
.B(n_703),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_499),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_596),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_499),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_499),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_596),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_523),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_636),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_607),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_523),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_497),
.B(n_370),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_607),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_523),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_499),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_523),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_632),
.B(n_703),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_632),
.B(n_703),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_499),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_523),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_499),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_499),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_499),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_632),
.B(n_703),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_618),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_L g1163 ( 
.A(n_618),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_497),
.B(n_370),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_596),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_638),
.B(n_344),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_499),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_497),
.B(n_370),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_499),
.Y(n_1169)
);

NOR3xp33_ASAP7_75t_L g1170 ( 
.A(n_685),
.B(n_313),
.C(n_385),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_613),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_523),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_607),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_636),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_523),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_632),
.B(n_703),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_523),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_499),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_523),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_499),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_596),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_596),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_497),
.B(n_370),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_499),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_675),
.A2(n_747),
.B1(n_751),
.B2(n_750),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_523),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_499),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_499),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_523),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_L g1190 ( 
.A(n_631),
.B(n_811),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_499),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_499),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_607),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_596),
.Y(n_1194)
);

OR2x6_ASAP7_75t_L g1195 ( 
.A(n_596),
.B(n_600),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_497),
.A2(n_370),
.B1(n_532),
.B2(n_685),
.Y(n_1196)
);

INVxp67_ASAP7_75t_SL g1197 ( 
.A(n_504),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_523),
.Y(n_1198)
);

NAND2xp33_ASAP7_75t_R g1199 ( 
.A(n_641),
.B(n_460),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_641),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_499),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_638),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_499),
.Y(n_1203)
);

NAND2xp33_ASAP7_75t_R g1204 ( 
.A(n_641),
.B(n_460),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_715),
.B(n_731),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_499),
.Y(n_1206)
);

NAND2xp33_ASAP7_75t_SL g1207 ( 
.A(n_613),
.B(n_596),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_499),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_499),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_523),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_523),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_499),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_638),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_638),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_499),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_638),
.B(n_344),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_499),
.Y(n_1217)
);

AND2x6_ASAP7_75t_L g1218 ( 
.A(n_617),
.B(n_550),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_596),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_675),
.B(n_460),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_632),
.B(n_703),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_601),
.A2(n_550),
.B(n_538),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_523),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_523),
.Y(n_1224)
);

NOR2x1p5_ASAP7_75t_L g1225 ( 
.A(n_596),
.B(n_469),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_523),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_523),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_499),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_632),
.B(n_703),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_523),
.Y(n_1230)
);

NAND2xp33_ASAP7_75t_SL g1231 ( 
.A(n_613),
.B(n_596),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_675),
.B(n_460),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_499),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_497),
.B(n_370),
.Y(n_1234)
);

AO21x2_ASAP7_75t_L g1235 ( 
.A1(n_550),
.A2(n_770),
.B(n_718),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_523),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_499),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_499),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_499),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_497),
.B(n_370),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_499),
.Y(n_1241)
);

AND3x2_ASAP7_75t_L g1242 ( 
.A(n_555),
.B(n_344),
.C(n_396),
.Y(n_1242)
);

NAND2xp33_ASAP7_75t_L g1243 ( 
.A(n_631),
.B(n_811),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_715),
.B(n_731),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_499),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_499),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_499),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_632),
.B(n_703),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_638),
.B(n_344),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_632),
.B(n_703),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_499),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_607),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_497),
.B(n_370),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_596),
.B(n_600),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_632),
.B(n_703),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_523),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_523),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_496),
.A2(n_722),
.B1(n_617),
.B2(n_550),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_607),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_596),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_632),
.B(n_703),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_498),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_523),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_607),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_499),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_499),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_523),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_499),
.Y(n_1268)
);

AND3x2_ASAP7_75t_L g1269 ( 
.A(n_555),
.B(n_344),
.C(n_396),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_632),
.B(n_703),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_607),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_523),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_632),
.B(n_703),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_632),
.B(n_703),
.Y(n_1274)
);

AND2x2_ASAP7_75t_SL g1275 ( 
.A(n_532),
.B(n_497),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_837),
.B(n_814),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_821),
.Y(n_1277)
);

NAND2xp33_ASAP7_75t_R g1278 ( 
.A(n_924),
.B(n_827),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_877),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_822),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_825),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_829),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_856),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1216),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_859),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_861),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_864),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_868),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1249),
.B(n_867),
.Y(n_1290)
);

OR2x6_ASAP7_75t_L g1291 ( 
.A(n_1129),
.B(n_1095),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_901),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_R g1293 ( 
.A(n_845),
.B(n_875),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_873),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_862),
.B(n_911),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_882),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1081),
.B(n_832),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_883),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_895),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1109),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1129),
.Y(n_1301)
);

XOR2xp5_ASAP7_75t_L g1302 ( 
.A(n_983),
.B(n_1171),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1047),
.A2(n_840),
.B(n_957),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_896),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_899),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_820),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_902),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_904),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1220),
.B(n_1232),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_907),
.Y(n_1310)
);

INVxp33_ASAP7_75t_SL g1311 ( 
.A(n_847),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1275),
.B(n_1056),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1205),
.B(n_1244),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_818),
.B(n_819),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1085),
.B(n_1144),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_913),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1202),
.B(n_1075),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_842),
.B(n_964),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1258),
.B(n_828),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1138),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1067),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_853),
.A2(n_1049),
.B(n_1235),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_914),
.Y(n_1323)
);

INVxp33_ASAP7_75t_L g1324 ( 
.A(n_1060),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_942),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1185),
.B(n_1196),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_830),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_920),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_922),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_926),
.Y(n_1330)
);

XNOR2x2_ASAP7_75t_L g1331 ( 
.A(n_1050),
.B(n_1058),
.Y(n_1331)
);

CKINVDCx16_ASAP7_75t_R g1332 ( 
.A(n_1199),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1052),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1054),
.Y(n_1334)
);

AOI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1042),
.A2(n_891),
.B(n_1222),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_833),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1055),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1131),
.B(n_1213),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1061),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_834),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_835),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1063),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1200),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1068),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1080),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1084),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1088),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1090),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1086),
.B(n_1146),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1214),
.B(n_1174),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1204),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1097),
.Y(n_1352)
);

NAND2xp33_ASAP7_75t_SL g1353 ( 
.A(n_831),
.B(n_1076),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1110),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1207),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_841),
.Y(n_1356)
);

INVxp67_ASAP7_75t_SL g1357 ( 
.A(n_831),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_843),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1113),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_878),
.Y(n_1360)
);

OR2x6_ASAP7_75t_L g1361 ( 
.A(n_1095),
.B(n_1195),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_849),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1120),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1053),
.B(n_1057),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1114),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1125),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1077),
.B(n_1078),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1105),
.B(n_1106),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1128),
.B(n_1079),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1133),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_879),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1138),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1134),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1135),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1140),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1099),
.B(n_1108),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1142),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1143),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1152),
.Y(n_1379)
);

XOR2xp5_ASAP7_75t_L g1380 ( 
.A(n_1070),
.B(n_1013),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_854),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1111),
.B(n_1122),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1156),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1195),
.B(n_1254),
.Y(n_1384)
);

NAND2xp33_ASAP7_75t_R g1385 ( 
.A(n_917),
.B(n_1242),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1158),
.Y(n_1386)
);

XOR2xp5_ASAP7_75t_L g1387 ( 
.A(n_934),
.B(n_857),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1149),
.B(n_1164),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1159),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1160),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1167),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1254),
.B(n_871),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1169),
.Y(n_1393)
);

XOR2xp5_ASAP7_75t_L g1394 ( 
.A(n_931),
.B(n_893),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_870),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1025),
.B(n_916),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1178),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1076),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1180),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1184),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1187),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1231),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1188),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_880),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_885),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1191),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1192),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1165),
.B(n_950),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1137),
.B(n_1139),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_886),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1168),
.B(n_1183),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1234),
.B(n_1240),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1201),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1203),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1154),
.B(n_1155),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1206),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_929),
.B(n_961),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1208),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1209),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1212),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1161),
.B(n_1176),
.Y(n_1421)
);

XNOR2xp5_ASAP7_75t_L g1422 ( 
.A(n_1269),
.B(n_995),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1221),
.B(n_1229),
.Y(n_1423)
);

XOR2xp5_ASAP7_75t_L g1424 ( 
.A(n_943),
.B(n_816),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1253),
.B(n_1248),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1250),
.B(n_1255),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1262),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1062),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1062),
.B(n_1124),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1261),
.B(n_1270),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1273),
.B(n_1274),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1215),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1217),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1228),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1233),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1237),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1238),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_927),
.B(n_1119),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1119),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_846),
.B(n_838),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1239),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1241),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1245),
.Y(n_1443)
);

XOR2xp5_ASAP7_75t_L g1444 ( 
.A(n_1074),
.B(n_1103),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1246),
.Y(n_1445)
);

XOR2xp5_ASAP7_75t_L g1446 ( 
.A(n_1018),
.B(n_888),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1130),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_887),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_817),
.B(n_823),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_SL g1450 ( 
.A(n_1130),
.B(n_1141),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1116),
.B(n_1218),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1126),
.B(n_815),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_874),
.B(n_889),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_892),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1247),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1251),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_905),
.B(n_915),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_824),
.B(n_826),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1265),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1266),
.Y(n_1460)
);

INVxp33_ASAP7_75t_L g1461 ( 
.A(n_1141),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1181),
.B(n_1182),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_919),
.B(n_928),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1268),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_930),
.B(n_848),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_863),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_966),
.A2(n_936),
.B(n_1048),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1181),
.Y(n_1468)
);

XOR2xp5_ASAP7_75t_L g1469 ( 
.A(n_1132),
.B(n_1016),
.Y(n_1469)
);

XOR2xp5_ASAP7_75t_L g1470 ( 
.A(n_1182),
.B(n_1194),
.Y(n_1470)
);

XOR2xp5_ASAP7_75t_L g1471 ( 
.A(n_1194),
.B(n_1219),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_939),
.B(n_1219),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1048),
.A2(n_866),
.B(n_865),
.Y(n_1473)
);

INVxp33_ASAP7_75t_SL g1474 ( 
.A(n_1009),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_872),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_876),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1260),
.B(n_963),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_940),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_890),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_898),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_910),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_912),
.B(n_1260),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1015),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_978),
.B(n_985),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_938),
.Y(n_1485)
);

BUFx8_ASAP7_75t_L g1486 ( 
.A(n_897),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_994),
.B(n_1033),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_941),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_881),
.B(n_900),
.Y(n_1489)
);

CKINVDCx14_ASAP7_75t_R g1490 ( 
.A(n_1163),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_908),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_897),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_1124),
.B(n_1162),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_949),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1116),
.A2(n_1218),
.B(n_1045),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_906),
.B(n_923),
.Y(n_1496)
);

XNOR2xp5_ASAP7_75t_L g1497 ( 
.A(n_1225),
.B(n_858),
.Y(n_1497)
);

XOR2xp5_ASAP7_75t_L g1498 ( 
.A(n_954),
.B(n_1066),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1087),
.B(n_1100),
.Y(n_1499)
);

AND2x6_ASAP7_75t_L g1500 ( 
.A(n_982),
.B(n_1044),
.Y(n_1500)
);

XOR2xp5_ASAP7_75t_L g1501 ( 
.A(n_1107),
.B(n_1117),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_956),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1162),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_836),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_959),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_968),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_925),
.B(n_812),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_970),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_947),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_948),
.Y(n_1510)
);

INVxp33_ASAP7_75t_L g1511 ( 
.A(n_908),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_974),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_977),
.Y(n_1513)
);

CKINVDCx20_ASAP7_75t_R g1514 ( 
.A(n_1147),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_990),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_998),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1001),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_952),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1046),
.A2(n_903),
.B(n_1022),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_813),
.B(n_1064),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_988),
.A2(n_969),
.B(n_946),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1197),
.B(n_1272),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1065),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1069),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1072),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1082),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_953),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1083),
.B(n_1089),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1091),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1093),
.B(n_1094),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1098),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1116),
.B(n_1218),
.Y(n_1532)
);

INVx8_ASAP7_75t_L g1533 ( 
.A(n_921),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1102),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1104),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_975),
.A2(n_937),
.B(n_1006),
.Y(n_1536)
);

XOR2xp5_ASAP7_75t_L g1537 ( 
.A(n_1259),
.B(n_1264),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1112),
.Y(n_1538)
);

XOR2xp5_ASAP7_75t_L g1539 ( 
.A(n_884),
.B(n_932),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1118),
.Y(n_1540)
);

INVxp33_ASAP7_75t_L g1541 ( 
.A(n_932),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1121),
.B(n_1127),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1071),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1136),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_935),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_955),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1145),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1148),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_852),
.B(n_1151),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1153),
.B(n_1157),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1172),
.B(n_1175),
.Y(n_1551)
);

XOR2xp5_ASAP7_75t_L g1552 ( 
.A(n_935),
.B(n_960),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1177),
.A2(n_1186),
.B(n_1267),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_960),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_958),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1179),
.B(n_1189),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1198),
.Y(n_1557)
);

INVx3_ASAP7_75t_R g1558 ( 
.A(n_1035),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1210),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_839),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1211),
.B(n_1223),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1224),
.B(n_1226),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1227),
.B(n_1230),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_965),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1236),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1031),
.B(n_1256),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1257),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_844),
.B(n_1051),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1263),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_981),
.Y(n_1570)
);

XOR2xp5_ASAP7_75t_L g1571 ( 
.A(n_986),
.B(n_1014),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_987),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1003),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1012),
.B(n_1026),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_852),
.B(n_967),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1029),
.B(n_921),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1004),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_851),
.B(n_860),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_971),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_852),
.B(n_973),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1007),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_976),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_855),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_921),
.B(n_1271),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_894),
.B(n_1020),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_979),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_980),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1021),
.B(n_1024),
.Y(n_1588)
);

XNOR2xp5_ASAP7_75t_L g1589 ( 
.A(n_996),
.B(n_1170),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_997),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1059),
.B(n_1252),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_984),
.Y(n_1592)
);

CKINVDCx16_ASAP7_75t_R g1593 ( 
.A(n_1027),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_989),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1028),
.B(n_1002),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_SL g1596 ( 
.A(n_1041),
.B(n_1030),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_909),
.B(n_972),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1096),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_991),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_993),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1000),
.B(n_1005),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1034),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_951),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_SL g1604 ( 
.A(n_1023),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1019),
.Y(n_1605)
);

XNOR2xp5_ASAP7_75t_L g1606 ( 
.A(n_1101),
.B(n_1193),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_918),
.B(n_1011),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_945),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_1115),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1008),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_933),
.B(n_944),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1010),
.Y(n_1612)
);

XNOR2xp5_ASAP7_75t_L g1613 ( 
.A(n_1123),
.B(n_1173),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1039),
.Y(n_1614)
);

NOR2xp67_ASAP7_75t_L g1615 ( 
.A(n_1150),
.B(n_1032),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_850),
.A2(n_869),
.B(n_1190),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_962),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_999),
.Y(n_1618)
);

XOR2xp5_ASAP7_75t_L g1619 ( 
.A(n_1043),
.B(n_1040),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1017),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1092),
.B(n_1243),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_992),
.B(n_1036),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1038),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1037),
.B(n_837),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_821),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_821),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_942),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_821),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_842),
.B(n_964),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_842),
.B(n_964),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_821),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_821),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_942),
.Y(n_1633)
);

INVxp67_ASAP7_75t_SL g1634 ( 
.A(n_842),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1129),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_832),
.B(n_818),
.Y(n_1636)
);

XOR2xp5_ASAP7_75t_L g1637 ( 
.A(n_983),
.B(n_656),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_821),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_821),
.Y(n_1639)
);

BUFx6f_ASAP7_75t_SL g1640 ( 
.A(n_836),
.Y(n_1640)
);

OR2x6_ASAP7_75t_L g1641 ( 
.A(n_1129),
.B(n_596),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_821),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_821),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_R g1644 ( 
.A(n_924),
.B(n_613),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_821),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_821),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_842),
.B(n_964),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_821),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1128),
.A2(n_840),
.B(n_832),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_832),
.B(n_818),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_831),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_820),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_821),
.Y(n_1654)
);

XNOR2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1242),
.B(n_656),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_821),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_820),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_832),
.B(n_818),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1129),
.Y(n_1660)
);

XNOR2x2_ASAP7_75t_L g1661 ( 
.A(n_814),
.B(n_1081),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_942),
.Y(n_1662)
);

XNOR2x2_ASAP7_75t_L g1663 ( 
.A(n_814),
.B(n_1081),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_942),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_821),
.Y(n_1665)
);

XOR2xp5_ASAP7_75t_L g1666 ( 
.A(n_983),
.B(n_656),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_821),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_842),
.B(n_964),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_821),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_821),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_837),
.B(n_814),
.Y(n_1671)
);

AND2x2_ASAP7_75t_SL g1672 ( 
.A(n_1275),
.B(n_532),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_831),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_821),
.Y(n_1674)
);

XNOR2x2_ASAP7_75t_L g1675 ( 
.A(n_814),
.B(n_1081),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1085),
.B(n_596),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_821),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_821),
.Y(n_1678)
);

XOR2xp5_ASAP7_75t_L g1679 ( 
.A(n_983),
.B(n_656),
.Y(n_1679)
);

XOR2xp5_ASAP7_75t_L g1680 ( 
.A(n_983),
.B(n_656),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1129),
.Y(n_1681)
);

XOR2xp5_ASAP7_75t_L g1682 ( 
.A(n_983),
.B(n_656),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_821),
.Y(n_1683)
);

XOR2xp5_ASAP7_75t_L g1684 ( 
.A(n_983),
.B(n_656),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_821),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1109),
.B(n_1205),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1129),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_942),
.Y(n_1688)
);

XOR2xp5_ASAP7_75t_L g1689 ( 
.A(n_983),
.B(n_656),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_821),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_942),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_821),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_820),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_821),
.Y(n_1694)
);

CKINVDCx20_ASAP7_75t_R g1695 ( 
.A(n_942),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_821),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_942),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_942),
.Y(n_1698)
);

AND2x6_ASAP7_75t_L g1699 ( 
.A(n_931),
.B(n_957),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_821),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_837),
.B(n_814),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_821),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_821),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_820),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_821),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_821),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_842),
.B(n_964),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_831),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_820),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_821),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_820),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_821),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_821),
.Y(n_1713)
);

CKINVDCx20_ASAP7_75t_R g1714 ( 
.A(n_942),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1129),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_832),
.B(n_818),
.Y(n_1717)
);

CKINVDCx20_ASAP7_75t_R g1718 ( 
.A(n_942),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_821),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_821),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_821),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_821),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_821),
.Y(n_1723)
);

CKINVDCx16_ASAP7_75t_R g1724 ( 
.A(n_847),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_837),
.B(n_814),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_942),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1129),
.Y(n_1727)
);

NAND2x1p5_ASAP7_75t_L g1728 ( 
.A(n_1085),
.B(n_596),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_820),
.Y(n_1729)
);

XOR2xp5_ASAP7_75t_L g1730 ( 
.A(n_983),
.B(n_656),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_942),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_942),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_821),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_821),
.Y(n_1734)
);

XOR2xp5_ASAP7_75t_L g1735 ( 
.A(n_983),
.B(n_656),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_942),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1129),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_837),
.B(n_814),
.Y(n_1738)
);

CKINVDCx20_ASAP7_75t_R g1739 ( 
.A(n_942),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_842),
.B(n_964),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_821),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_821),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_820),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_R g1744 ( 
.A(n_924),
.B(n_613),
.Y(n_1744)
);

NOR2xp33_ASAP7_75t_SL g1745 ( 
.A(n_847),
.B(n_716),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_821),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_821),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_837),
.B(n_814),
.Y(n_1749)
);

INVxp33_ASAP7_75t_L g1750 ( 
.A(n_1073),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_837),
.B(n_814),
.Y(n_1751)
);

INVxp33_ASAP7_75t_L g1752 ( 
.A(n_1073),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_837),
.B(n_814),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1128),
.A2(n_840),
.B(n_832),
.Y(n_1754)
);

CKINVDCx20_ASAP7_75t_R g1755 ( 
.A(n_942),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1073),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_821),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_821),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_821),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1073),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_821),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_842),
.B(n_964),
.Y(n_1762)
);

XOR2xp5_ASAP7_75t_L g1763 ( 
.A(n_983),
.B(n_656),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_821),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_821),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_821),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_821),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1109),
.B(n_1205),
.Y(n_1768)
);

INVxp33_ASAP7_75t_L g1769 ( 
.A(n_1073),
.Y(n_1769)
);

AND2x2_ASAP7_75t_SL g1770 ( 
.A(n_1275),
.B(n_532),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_821),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_842),
.B(n_964),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_821),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_821),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_821),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_832),
.B(n_497),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_821),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_821),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_821),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_820),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_821),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_821),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_821),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_821),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_821),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_821),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_821),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_821),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_821),
.Y(n_1790)
);

XNOR2xp5_ASAP7_75t_L g1791 ( 
.A(n_983),
.B(n_656),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_837),
.B(n_814),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_821),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_831),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_837),
.B(n_814),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_821),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_821),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_821),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_821),
.Y(n_1799)
);

XOR2xp5_ASAP7_75t_L g1800 ( 
.A(n_983),
.B(n_656),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_821),
.Y(n_1801)
);

XOR2xp5_ASAP7_75t_L g1802 ( 
.A(n_983),
.B(n_656),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_821),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_821),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_821),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_821),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_821),
.Y(n_1807)
);

INVxp33_ASAP7_75t_L g1808 ( 
.A(n_1073),
.Y(n_1808)
);

NAND2x1p5_ASAP7_75t_L g1809 ( 
.A(n_1085),
.B(n_596),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_832),
.B(n_818),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_821),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_821),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_821),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_821),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_821),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1816)
);

XOR2xp5_ASAP7_75t_L g1817 ( 
.A(n_983),
.B(n_656),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_942),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_837),
.B(n_814),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_821),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_821),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_821),
.Y(n_1823)
);

INVx2_ASAP7_75t_SL g1824 ( 
.A(n_1129),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_821),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_821),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_842),
.B(n_964),
.Y(n_1827)
);

INVx8_ASAP7_75t_L g1828 ( 
.A(n_1129),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_842),
.B(n_964),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_821),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_821),
.Y(n_1831)
);

XOR2xp5_ASAP7_75t_L g1832 ( 
.A(n_983),
.B(n_656),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_821),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_821),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_820),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_821),
.Y(n_1836)
);

INVx2_ASAP7_75t_SL g1837 ( 
.A(n_1129),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_842),
.B(n_964),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_821),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1129),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_837),
.B(n_814),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_821),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_821),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_821),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1129),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_832),
.B(n_818),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1109),
.B(n_1205),
.Y(n_1847)
);

OAI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1128),
.A2(n_840),
.B(n_832),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_831),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_837),
.B(n_814),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_820),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_821),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_821),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_821),
.Y(n_1854)
);

CKINVDCx16_ASAP7_75t_R g1855 ( 
.A(n_847),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_821),
.Y(n_1856)
);

NOR2xp67_ASAP7_75t_L g1857 ( 
.A(n_1171),
.B(n_423),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_SL g1858 ( 
.A(n_847),
.B(n_716),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1109),
.B(n_1205),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_832),
.B(n_818),
.Y(n_1860)
);

XOR2xp5_ASAP7_75t_L g1861 ( 
.A(n_983),
.B(n_656),
.Y(n_1861)
);

XNOR2xp5_ASAP7_75t_L g1862 ( 
.A(n_983),
.B(n_656),
.Y(n_1862)
);

XOR2xp5_ASAP7_75t_L g1863 ( 
.A(n_983),
.B(n_656),
.Y(n_1863)
);

CKINVDCx20_ASAP7_75t_R g1864 ( 
.A(n_942),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_837),
.B(n_814),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_821),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_821),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_SL g1869 ( 
.A(n_847),
.B(n_716),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_821),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_837),
.B(n_814),
.Y(n_1872)
);

XOR2xp5_ASAP7_75t_L g1873 ( 
.A(n_983),
.B(n_656),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_821),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_821),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_837),
.B(n_814),
.Y(n_1876)
);

INVxp33_ASAP7_75t_L g1877 ( 
.A(n_1073),
.Y(n_1877)
);

OAI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1128),
.A2(n_840),
.B(n_832),
.Y(n_1878)
);

BUFx3_ASAP7_75t_L g1879 ( 
.A(n_1129),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_820),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_821),
.Y(n_1881)
);

XOR2xp5_ASAP7_75t_L g1882 ( 
.A(n_983),
.B(n_656),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1109),
.B(n_1205),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_820),
.Y(n_1884)
);

XNOR2xp5_ASAP7_75t_L g1885 ( 
.A(n_983),
.B(n_656),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_832),
.B(n_818),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_837),
.B(n_814),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_837),
.B(n_814),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1109),
.B(n_1205),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1128),
.A2(n_840),
.B(n_832),
.Y(n_1890)
);

NAND2xp33_ASAP7_75t_R g1891 ( 
.A(n_924),
.B(n_613),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_821),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_821),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_832),
.B(n_818),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_821),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_821),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_821),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_821),
.Y(n_1898)
);

BUFx3_ASAP7_75t_L g1899 ( 
.A(n_1129),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_832),
.B(n_818),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_821),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_821),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_821),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_821),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_820),
.Y(n_1906)
);

AND2x2_ASAP7_75t_SL g1907 ( 
.A(n_1275),
.B(n_532),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_821),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_837),
.B(n_814),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_821),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_821),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_821),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1129),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_821),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_821),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1109),
.B(n_1205),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_820),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_842),
.B(n_964),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_820),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_821),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_842),
.B(n_964),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_821),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_821),
.Y(n_1924)
);

NOR2x1p5_ASAP7_75t_L g1925 ( 
.A(n_1025),
.B(n_405),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_832),
.B(n_818),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_820),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_837),
.B(n_814),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_821),
.Y(n_1929)
);

NAND2x1p5_ASAP7_75t_L g1930 ( 
.A(n_1085),
.B(n_596),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_821),
.Y(n_1931)
);

INVx2_ASAP7_75t_SL g1932 ( 
.A(n_1129),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_821),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_821),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_837),
.B(n_814),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_842),
.B(n_964),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_821),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_821),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_821),
.Y(n_1940)
);

XNOR2x2_ASAP7_75t_L g1941 ( 
.A(n_814),
.B(n_1081),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_821),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_820),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1073),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1129),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_821),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_820),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_821),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_820),
.Y(n_1949)
);

XNOR2xp5_ASAP7_75t_L g1950 ( 
.A(n_983),
.B(n_656),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_821),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_821),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_821),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_821),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_821),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_821),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_821),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_820),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_821),
.Y(n_1959)
);

XOR2x2_ASAP7_75t_L g1960 ( 
.A(n_1170),
.B(n_685),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_821),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1047),
.A2(n_832),
.B(n_840),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1073),
.B(n_1166),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_821),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_821),
.Y(n_1965)
);

INVxp33_ASAP7_75t_L g1966 ( 
.A(n_1073),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_821),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_821),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_821),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_821),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_821),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_821),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_877),
.Y(n_1973)
);

CKINVDCx11_ASAP7_75t_R g1974 ( 
.A(n_836),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_821),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_837),
.B(n_814),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_821),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_821),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_821),
.Y(n_1979)
);

OAI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1128),
.A2(n_840),
.B(n_832),
.Y(n_1980)
);

XOR2x2_ASAP7_75t_L g1981 ( 
.A(n_1170),
.B(n_685),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_821),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_832),
.B(n_818),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_832),
.B(n_497),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_837),
.B(n_814),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_821),
.Y(n_1986)
);

XOR2xp5_ASAP7_75t_L g1987 ( 
.A(n_983),
.B(n_656),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_821),
.Y(n_1988)
);

XOR2xp5_ASAP7_75t_L g1989 ( 
.A(n_983),
.B(n_656),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_821),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_821),
.Y(n_1991)
);

XNOR2x2_ASAP7_75t_L g1992 ( 
.A(n_814),
.B(n_1081),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1073),
.Y(n_1993)
);

INVxp33_ASAP7_75t_L g1994 ( 
.A(n_1073),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1047),
.A2(n_832),
.B(n_840),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_821),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_821),
.Y(n_1997)
);

INVxp33_ASAP7_75t_L g1998 ( 
.A(n_1073),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_832),
.B(n_818),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_821),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_821),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1073),
.B(n_1166),
.Y(n_2002)
);

AND2x2_ASAP7_75t_SL g2003 ( 
.A(n_1275),
.B(n_532),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_942),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1073),
.B(n_1166),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_842),
.B(n_964),
.Y(n_2006)
);

XNOR2xp5_ASAP7_75t_L g2007 ( 
.A(n_983),
.B(n_656),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2009)
);

OAI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1650),
.A2(n_1848),
.B(n_1754),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1367),
.B(n_1368),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1878),
.B(n_1890),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1486),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1646),
.B(n_1658),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1380),
.A2(n_1474),
.B1(n_1701),
.B2(n_1671),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_1725),
.B(n_1738),
.Y(n_2017)
);

A2O1A1Ixp33_ASAP7_75t_L g2018 ( 
.A1(n_1369),
.A2(n_1749),
.B(n_1753),
.C(n_1751),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1980),
.B(n_1314),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1277),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1281),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1792),
.B(n_1795),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1382),
.B(n_1415),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1819),
.B(n_1841),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1421),
.A2(n_1426),
.B1(n_1423),
.B2(n_1409),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1430),
.B(n_1651),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1850),
.B(n_1865),
.Y(n_2027)
);

INVxp67_ASAP7_75t_L g2028 ( 
.A(n_1686),
.Y(n_2028)
);

NAND2x1p5_ASAP7_75t_L g2029 ( 
.A(n_1576),
.B(n_1584),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1860),
.B(n_1999),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1282),
.Y(n_2031)
);

INVxp67_ASAP7_75t_L g2032 ( 
.A(n_1768),
.Y(n_2032)
);

INVx4_ASAP7_75t_L g2033 ( 
.A(n_1828),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1810),
.B(n_1636),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1872),
.A2(n_1876),
.B1(n_1888),
.B2(n_1887),
.Y(n_2035)
);

OAI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_1909),
.A2(n_1928),
.B1(n_1985),
.B2(n_1976),
.C(n_1935),
.Y(n_2036)
);

NOR2xp67_ASAP7_75t_SL g2037 ( 
.A(n_1724),
.B(n_1855),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1983),
.B(n_1659),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1457),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1283),
.Y(n_2040)
);

BUFx3_ASAP7_75t_L g2041 ( 
.A(n_1486),
.Y(n_2041)
);

BUFx8_ASAP7_75t_L g2042 ( 
.A(n_1640),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1717),
.A2(n_1886),
.B1(n_1894),
.B2(n_1846),
.Y(n_2043)
);

INVx2_ASAP7_75t_SL g2044 ( 
.A(n_1641),
.Y(n_2044)
);

INVx2_ASAP7_75t_SL g2045 ( 
.A(n_1641),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1715),
.B(n_1748),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1425),
.B(n_1900),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1926),
.B(n_1297),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1463),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1458),
.B(n_1452),
.Y(n_2050)
);

AND2x4_ASAP7_75t_L g2051 ( 
.A(n_1584),
.B(n_1318),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1326),
.A2(n_1770),
.B1(n_1907),
.B2(n_1672),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1466),
.B(n_1475),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_1828),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1284),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1286),
.Y(n_2056)
);

O2A1O1Ixp33_ASAP7_75t_L g2057 ( 
.A1(n_1312),
.A2(n_1319),
.B(n_1984),
.C(n_1776),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1476),
.B(n_1479),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_1847),
.B(n_1859),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1624),
.B(n_1449),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1287),
.Y(n_2061)
);

O2A1O1Ixp33_ASAP7_75t_L g2062 ( 
.A1(n_1496),
.A2(n_1292),
.B(n_1388),
.C(n_1376),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1480),
.B(n_1481),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1295),
.B(n_1440),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1785),
.B(n_1816),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2002),
.B(n_2005),
.Y(n_2066)
);

BUFx3_ASAP7_75t_L g2067 ( 
.A(n_1514),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_2003),
.A2(n_1868),
.B1(n_1870),
.B2(n_1820),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1903),
.B(n_1916),
.Y(n_2069)
);

INVx3_ASAP7_75t_L g2070 ( 
.A(n_1533),
.Y(n_2070)
);

INVx4_ASAP7_75t_L g2071 ( 
.A(n_1462),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1937),
.B(n_1963),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1515),
.B(n_1516),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1411),
.A2(n_1412),
.B1(n_1590),
.B2(n_1571),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1288),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1517),
.B(n_1487),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1289),
.Y(n_2077)
);

OR2x6_ASAP7_75t_L g2078 ( 
.A(n_1533),
.B(n_1361),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_1883),
.B(n_1889),
.Y(n_2079)
);

NAND2xp33_ASAP7_75t_L g2080 ( 
.A(n_1699),
.B(n_1402),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1303),
.B(n_1473),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1294),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1616),
.B(n_1536),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1313),
.B(n_1917),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1699),
.B(n_1482),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1699),
.B(n_1483),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1621),
.A2(n_1387),
.B1(n_1620),
.B2(n_1618),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_1438),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1296),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1699),
.B(n_1453),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1962),
.B(n_1995),
.Y(n_2091)
);

AND2x4_ASAP7_75t_L g2092 ( 
.A(n_1318),
.B(n_1629),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1298),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1623),
.B(n_1993),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_1750),
.B(n_1752),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1769),
.B(n_1808),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1629),
.B(n_1630),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1285),
.B(n_1756),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1760),
.B(n_1944),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1521),
.B(n_1495),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1520),
.B(n_1530),
.Y(n_2101)
);

AOI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_1300),
.A2(n_1394),
.B1(n_1877),
.B2(n_1994),
.C(n_1966),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1299),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1542),
.B(n_1550),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1556),
.B(n_1563),
.Y(n_2105)
);

O2A1O1Ixp5_ASAP7_75t_L g2106 ( 
.A1(n_1467),
.A2(n_1451),
.B(n_1532),
.C(n_1322),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1745),
.B(n_1858),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1869),
.B(n_1311),
.Y(n_2108)
);

NOR2xp33_ASAP7_75t_L g2109 ( 
.A(n_1998),
.B(n_1324),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1304),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1305),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1522),
.B(n_1561),
.Y(n_2112)
);

BUFx3_ASAP7_75t_L g2113 ( 
.A(n_1609),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1562),
.B(n_1307),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1308),
.B(n_1310),
.Y(n_2115)
);

BUFx6f_ASAP7_75t_L g2116 ( 
.A(n_1652),
.Y(n_2116)
);

INVx2_ASAP7_75t_SL g2117 ( 
.A(n_1438),
.Y(n_2117)
);

OAI221xp5_ASAP7_75t_L g2118 ( 
.A1(n_1446),
.A2(n_1981),
.B1(n_1960),
.B2(n_1891),
.C(n_1744),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_1992),
.A2(n_1661),
.B1(n_1675),
.B2(n_1663),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_1349),
.B(n_1279),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1316),
.A2(n_1328),
.B1(n_1329),
.B2(n_1323),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1332),
.B(n_1351),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1321),
.B(n_1973),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1330),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1549),
.B(n_1519),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1333),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1334),
.Y(n_2127)
);

AOI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_1644),
.A2(n_1278),
.B1(n_1355),
.B2(n_1293),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_1941),
.A2(n_1331),
.B1(n_1488),
.B2(n_1485),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1337),
.B(n_1339),
.Y(n_2130)
);

A2O1A1Ixp33_ASAP7_75t_L g2131 ( 
.A1(n_1507),
.A2(n_1603),
.B(n_1574),
.C(n_1580),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1342),
.B(n_1344),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1345),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_1371),
.B(n_1427),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1346),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1347),
.Y(n_2136)
);

INVx2_ASAP7_75t_SL g2137 ( 
.A(n_1396),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1348),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_SL g2139 ( 
.A(n_1575),
.B(n_1553),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1352),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1354),
.Y(n_2141)
);

BUFx12f_ASAP7_75t_L g2142 ( 
.A(n_1974),
.Y(n_2142)
);

INVx3_ASAP7_75t_L g2143 ( 
.A(n_1576),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1359),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_1343),
.B(n_1350),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1363),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_1317),
.B(n_1610),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_1612),
.B(n_1622),
.Y(n_2148)
);

BUFx12f_ASAP7_75t_L g2149 ( 
.A(n_1360),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_1461),
.B(n_1511),
.Y(n_2150)
);

AND2x6_ASAP7_75t_SL g2151 ( 
.A(n_1396),
.B(n_1392),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_1566),
.B(n_1422),
.Y(n_2152)
);

BUFx8_ASAP7_75t_L g2153 ( 
.A(n_1604),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_1541),
.B(n_1306),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1338),
.B(n_1484),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1366),
.B(n_1370),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_1327),
.B(n_1336),
.Y(n_2157)
);

INVx2_ASAP7_75t_SL g2158 ( 
.A(n_1681),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_1687),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1373),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_1340),
.B(n_1341),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1374),
.B(n_1375),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1377),
.B(n_1378),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1379),
.Y(n_2164)
);

AOI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_1385),
.A2(n_1648),
.B1(n_1668),
.B2(n_1630),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1383),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_1648),
.A2(n_1707),
.B1(n_1740),
.B2(n_1668),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1386),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1389),
.B(n_1390),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_1652),
.Y(n_2170)
);

CKINVDCx20_ASAP7_75t_R g2171 ( 
.A(n_1325),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1391),
.B(n_1393),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1397),
.B(n_1399),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1566),
.Y(n_2174)
);

AND2x4_ASAP7_75t_SL g2175 ( 
.A(n_1291),
.B(n_1384),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_1356),
.B(n_1358),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1465),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_1583),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1400),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_1465),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1401),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1403),
.B(n_1406),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1407),
.B(n_1413),
.Y(n_2183)
);

O2A1O1Ixp33_ASAP7_75t_L g2184 ( 
.A1(n_1602),
.A2(n_1502),
.B(n_1505),
.C(n_1494),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1414),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1416),
.B(n_1418),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1419),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1420),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1432),
.B(n_1433),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1434),
.B(n_1435),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1436),
.B(n_1437),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1362),
.B(n_1381),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1395),
.B(n_1404),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_1405),
.B(n_1410),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1441),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_1707),
.A2(n_1740),
.B1(n_1772),
.B2(n_1762),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1442),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1443),
.B(n_1445),
.Y(n_2198)
);

OR2x6_ASAP7_75t_L g2199 ( 
.A(n_1361),
.B(n_1291),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1455),
.B(n_1456),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1448),
.B(n_1454),
.Y(n_2201)
);

AOI22xp33_ASAP7_75t_L g2202 ( 
.A1(n_1506),
.A2(n_1512),
.B1(n_1513),
.B2(n_1508),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_1633),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1459),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_L g2205 ( 
.A(n_1596),
.B(n_1615),
.C(n_1589),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_1762),
.B(n_1772),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_1447),
.Y(n_2207)
);

AOI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_1827),
.A2(n_1838),
.B1(n_1919),
.B2(n_1829),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_1653),
.B(n_1657),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_1693),
.B(n_1704),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1460),
.B(n_1464),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_1827),
.B(n_1829),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1625),
.B(n_1626),
.Y(n_2213)
);

INVx2_ASAP7_75t_SL g2214 ( 
.A(n_1727),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1709),
.B(n_1711),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1628),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1631),
.B(n_1632),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1729),
.B(n_1743),
.Y(n_2218)
);

AOI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_1838),
.A2(n_1922),
.B1(n_1936),
.B2(n_1919),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1638),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_1528),
.A2(n_1551),
.B(n_1601),
.Y(n_2221)
);

INVx4_ASAP7_75t_L g2222 ( 
.A(n_1462),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1780),
.B(n_1835),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1639),
.Y(n_2224)
);

AND2x4_ASAP7_75t_SL g2225 ( 
.A(n_1384),
.B(n_1392),
.Y(n_2225)
);

NOR2xp33_ASAP7_75t_L g2226 ( 
.A(n_1851),
.B(n_1880),
.Y(n_2226)
);

O2A1O1Ixp33_ASAP7_75t_L g2227 ( 
.A1(n_1642),
.A2(n_1645),
.B(n_1647),
.C(n_1643),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1884),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_1906),
.B(n_1918),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_1920),
.B(n_1927),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_SL g2231 ( 
.A(n_1943),
.B(n_1947),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1949),
.B(n_1958),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1649),
.B(n_1654),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1656),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_1570),
.B(n_1572),
.Y(n_2235)
);

INVx8_ASAP7_75t_L g2236 ( 
.A(n_1652),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_1922),
.A2(n_2006),
.B1(n_1936),
.B2(n_1444),
.Y(n_2237)
);

AOI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_2006),
.A2(n_1302),
.B1(n_1666),
.B2(n_1637),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1665),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1667),
.Y(n_2240)
);

AOI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_1679),
.A2(n_1680),
.B1(n_1684),
.B2(n_1682),
.Y(n_2241)
);

HB1xp67_ASAP7_75t_L g2242 ( 
.A(n_1470),
.Y(n_2242)
);

NOR2xp33_ASAP7_75t_L g2243 ( 
.A(n_1669),
.B(n_1670),
.Y(n_2243)
);

AOI22xp33_ASAP7_75t_L g2244 ( 
.A1(n_1674),
.A2(n_1678),
.B1(n_1683),
.B2(n_1677),
.Y(n_2244)
);

INVx8_ASAP7_75t_L g2245 ( 
.A(n_1673),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1685),
.B(n_1690),
.Y(n_2246)
);

INVx2_ASAP7_75t_SL g2247 ( 
.A(n_1879),
.Y(n_2247)
);

BUFx3_ASAP7_75t_L g2248 ( 
.A(n_1899),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1692),
.B(n_1694),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1696),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1700),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_1477),
.B(n_1472),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1702),
.B(n_1703),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1705),
.Y(n_2254)
);

NAND3xp33_ASAP7_75t_SL g2255 ( 
.A(n_1598),
.B(n_1365),
.C(n_1469),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1706),
.B(n_1710),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1712),
.B(n_1713),
.Y(n_2257)
);

AOI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_1689),
.A2(n_1730),
.B1(n_1763),
.B2(n_1735),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1719),
.B(n_1720),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_1408),
.B(n_1417),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1721),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1722),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1723),
.B(n_1733),
.Y(n_2263)
);

OR2x6_ASAP7_75t_L g2264 ( 
.A(n_1676),
.B(n_1728),
.Y(n_2264)
);

INVx1_ASAP7_75t_SL g2265 ( 
.A(n_1539),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_1734),
.B(n_1741),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_1471),
.Y(n_2267)
);

INVx3_ASAP7_75t_L g2268 ( 
.A(n_1478),
.Y(n_2268)
);

NOR3xp33_ASAP7_75t_L g2269 ( 
.A(n_1593),
.B(n_1490),
.C(n_1634),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_1573),
.B(n_1577),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_1581),
.B(n_1742),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1746),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1747),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_1757),
.B(n_1758),
.Y(n_2274)
);

OAI22xp33_ASAP7_75t_L g2275 ( 
.A1(n_1759),
.A2(n_1764),
.B1(n_1765),
.B2(n_1761),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_1766),
.B(n_1767),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1771),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1773),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1774),
.B(n_1775),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1777),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_L g2281 ( 
.A(n_1778),
.B(n_1779),
.Y(n_2281)
);

O2A1O1Ixp5_ASAP7_75t_L g2282 ( 
.A1(n_1335),
.A2(n_1781),
.B(n_1783),
.C(n_1782),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_1784),
.B(n_1786),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1787),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_R g2285 ( 
.A(n_1543),
.B(n_1664),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1788),
.B(n_1789),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_1800),
.A2(n_1817),
.B1(n_1832),
.B2(n_1802),
.Y(n_2287)
);

BUFx8_ASAP7_75t_L g2288 ( 
.A(n_1468),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_1790),
.B(n_1793),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_1796),
.B(n_1797),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1798),
.B(n_1799),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_1489),
.B(n_1499),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1801),
.B(n_1803),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1804),
.B(n_1805),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1806),
.B(n_1807),
.Y(n_2295)
);

AND2x4_ASAP7_75t_L g2296 ( 
.A(n_1408),
.B(n_1417),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_1913),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1811),
.Y(n_2298)
);

NAND2xp33_ASAP7_75t_L g2299 ( 
.A(n_1812),
.B(n_1813),
.Y(n_2299)
);

O2A1O1Ixp33_ASAP7_75t_L g2300 ( 
.A1(n_1814),
.A2(n_1821),
.B(n_1822),
.C(n_1815),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1823),
.B(n_1825),
.Y(n_2301)
);

OAI221xp5_ASAP7_75t_L g2302 ( 
.A1(n_1497),
.A2(n_2007),
.B1(n_1885),
.B2(n_1950),
.C(n_1791),
.Y(n_2302)
);

INVx3_ASAP7_75t_L g2303 ( 
.A(n_1509),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_1826),
.B(n_1830),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1831),
.Y(n_2305)
);

AO221x1_ASAP7_75t_L g2306 ( 
.A1(n_1833),
.A2(n_1979),
.B1(n_1940),
.B2(n_2001),
.C(n_1939),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1834),
.Y(n_2307)
);

OAI22xp33_ASAP7_75t_L g2308 ( 
.A1(n_1836),
.A2(n_1959),
.B1(n_1874),
.B2(n_2000),
.Y(n_2308)
);

A2O1A1Ixp33_ASAP7_75t_L g2309 ( 
.A1(n_1605),
.A2(n_1569),
.B(n_1567),
.C(n_1565),
.Y(n_2309)
);

AND2x6_ASAP7_75t_L g2310 ( 
.A(n_1839),
.B(n_1842),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1843),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_1844),
.Y(n_2312)
);

NOR2xp67_ASAP7_75t_L g2313 ( 
.A(n_1737),
.B(n_1857),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1852),
.B(n_1853),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_1854),
.B(n_1856),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_L g2316 ( 
.A1(n_1866),
.A2(n_1965),
.B1(n_1964),
.B2(n_1961),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1867),
.B(n_1871),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_1875),
.B(n_1881),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1892),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1893),
.B(n_1895),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_1617),
.B(n_1673),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1896),
.Y(n_2322)
);

NOR2xp67_ASAP7_75t_L g2323 ( 
.A(n_1568),
.B(n_1429),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1897),
.Y(n_2324)
);

OAI22xp33_ASAP7_75t_L g2325 ( 
.A1(n_1898),
.A2(n_1914),
.B1(n_1912),
.B2(n_1911),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_1901),
.B(n_1902),
.Y(n_2326)
);

NAND2xp33_ASAP7_75t_L g2327 ( 
.A(n_1904),
.B(n_1905),
.Y(n_2327)
);

INVx2_ASAP7_75t_SL g2328 ( 
.A(n_1945),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_1908),
.B(n_1910),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_1915),
.B(n_1921),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_1923),
.B(n_1924),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_1861),
.A2(n_1873),
.B1(n_1882),
.B2(n_1863),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_L g2333 ( 
.A(n_1929),
.B(n_1931),
.Y(n_2333)
);

INVxp67_ASAP7_75t_L g2334 ( 
.A(n_1554),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1933),
.B(n_1934),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_1938),
.A2(n_1954),
.B1(n_1942),
.B2(n_1997),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_1946),
.B(n_1948),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_1951),
.B(n_1952),
.Y(n_2338)
);

NAND2x1p5_ASAP7_75t_L g2339 ( 
.A(n_1953),
.B(n_1955),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1956),
.B(n_1957),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_1967),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_1968),
.B(n_1969),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1970),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_SL g2344 ( 
.A(n_1971),
.B(n_1972),
.Y(n_2344)
);

O2A1O1Ixp33_ASAP7_75t_L g2345 ( 
.A1(n_1975),
.A2(n_1988),
.B(n_1996),
.C(n_1991),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1977),
.B(n_1978),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_1510),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_R g2348 ( 
.A(n_1691),
.B(n_1697),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_1982),
.B(n_1986),
.Y(n_2349)
);

AOI22xp33_ASAP7_75t_L g2350 ( 
.A1(n_1990),
.A2(n_1544),
.B1(n_1535),
.B2(n_1534),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1523),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_1524),
.B(n_1525),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1518),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1526),
.B(n_1529),
.Y(n_2354)
);

AOI22xp33_ASAP7_75t_L g2355 ( 
.A1(n_1531),
.A2(n_1538),
.B1(n_1540),
.B2(n_1559),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_1547),
.B(n_1548),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_1557),
.B(n_1582),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_1586),
.A2(n_1599),
.B1(n_1600),
.B2(n_1587),
.Y(n_2358)
);

NAND2x1_ASAP7_75t_L g2359 ( 
.A(n_1500),
.B(n_1594),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1527),
.B(n_1546),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_1987),
.B(n_1989),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1673),
.B(n_1708),
.Y(n_2362)
);

INVx2_ASAP7_75t_SL g2363 ( 
.A(n_1708),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_1862),
.B(n_1555),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_1564),
.Y(n_2365)
);

AOI22xp5_ASAP7_75t_L g2366 ( 
.A1(n_1619),
.A2(n_1424),
.B1(n_1925),
.B2(n_1498),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1579),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1592),
.B(n_1588),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_1595),
.B(n_1607),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_1708),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1614),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_L g2372 ( 
.A(n_1608),
.B(n_1492),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_1552),
.B(n_1560),
.Y(n_2373)
);

INVx2_ASAP7_75t_SL g2374 ( 
.A(n_1794),
.Y(n_2374)
);

A2O1A1Ixp33_ASAP7_75t_L g2375 ( 
.A1(n_1578),
.A2(n_1611),
.B(n_1597),
.C(n_1585),
.Y(n_2375)
);

BUFx3_ASAP7_75t_L g2376 ( 
.A(n_1794),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_1794),
.Y(n_2377)
);

AOI22xp33_ASAP7_75t_L g2378 ( 
.A1(n_1500),
.A2(n_1450),
.B1(n_1353),
.B2(n_1591),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_1591),
.B(n_1545),
.Y(n_2379)
);

AND2x2_ASAP7_75t_SL g2380 ( 
.A(n_1655),
.B(n_1439),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1500),
.Y(n_2381)
);

BUFx12f_ASAP7_75t_L g2382 ( 
.A(n_1726),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_1357),
.B(n_1606),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1613),
.B(n_1491),
.Y(n_2384)
);

BUFx3_ASAP7_75t_L g2385 ( 
.A(n_1849),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_1849),
.B(n_1809),
.Y(n_2386)
);

HB1xp67_ASAP7_75t_L g2387 ( 
.A(n_1493),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1500),
.Y(n_2388)
);

AOI22xp5_ASAP7_75t_L g2389 ( 
.A1(n_1501),
.A2(n_1537),
.B1(n_1732),
.B2(n_2004),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_1398),
.B(n_1849),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_1930),
.B(n_1315),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1320),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_1372),
.B(n_1558),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_1932),
.B(n_1301),
.Y(n_2394)
);

INVx3_ASAP7_75t_L g2395 ( 
.A(n_1635),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1660),
.B(n_1840),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_1716),
.B(n_1845),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_1824),
.B(n_1837),
.Y(n_2398)
);

OR2x6_ASAP7_75t_L g2399 ( 
.A(n_1504),
.B(n_1428),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_1503),
.B(n_1627),
.Y(n_2400)
);

OAI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_1662),
.A2(n_1864),
.B1(n_1695),
.B2(n_1698),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_1688),
.B(n_1714),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1718),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_1731),
.B(n_1736),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_1818),
.Y(n_2405)
);

AND2x6_ASAP7_75t_L g2406 ( 
.A(n_1739),
.B(n_1755),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1277),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_1277),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1277),
.Y(n_2413)
);

OAI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_1431),
.A2(n_1314),
.B1(n_1415),
.B2(n_1382),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_1277),
.Y(n_2417)
);

NAND2xp33_ASAP7_75t_L g2418 ( 
.A(n_1314),
.B(n_1382),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_1277),
.Y(n_2419)
);

HB1xp67_ASAP7_75t_L g2420 ( 
.A(n_1427),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1277),
.Y(n_2421)
);

NOR3x1_ASAP7_75t_L g2422 ( 
.A(n_1634),
.B(n_857),
.C(n_616),
.Y(n_2422)
);

AOI22xp33_ASAP7_75t_L g2423 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_SL g2424 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2424)
);

OR2x2_ASAP7_75t_L g2425 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2427)
);

A2O1A1Ixp33_ASAP7_75t_L g2428 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1277),
.Y(n_2429)
);

INVx2_ASAP7_75t_SL g2430 ( 
.A(n_1486),
.Y(n_2430)
);

NOR2xp33_ASAP7_75t_SL g2431 ( 
.A(n_1745),
.B(n_716),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_1427),
.Y(n_2432)
);

OAI22xp5_ASAP7_75t_L g2433 ( 
.A1(n_1431),
.A2(n_1314),
.B1(n_1415),
.B2(n_1382),
.Y(n_2433)
);

NOR3xp33_ASAP7_75t_L g2434 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_1533),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_1277),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_1457),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_SL g2444 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2444)
);

INVxp67_ASAP7_75t_L g2445 ( 
.A(n_1686),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_1277),
.Y(n_2447)
);

O2A1O1Ixp33_ASAP7_75t_L g2448 ( 
.A1(n_1326),
.A2(n_1128),
.B(n_747),
.C(n_750),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2450)
);

OR2x2_ASAP7_75t_L g2451 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2451)
);

INVx2_ASAP7_75t_SL g2452 ( 
.A(n_1486),
.Y(n_2452)
);

INVx8_ASAP7_75t_L g2453 ( 
.A(n_1828),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2454)
);

NOR2xp67_ASAP7_75t_L g2455 ( 
.A(n_1349),
.B(n_716),
.Y(n_2455)
);

O2A1O1Ixp33_ASAP7_75t_L g2456 ( 
.A1(n_1326),
.A2(n_1128),
.B(n_747),
.C(n_750),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1277),
.Y(n_2457)
);

INVxp67_ASAP7_75t_L g2458 ( 
.A(n_1686),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1277),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_1457),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2464)
);

INVx8_ASAP7_75t_L g2465 ( 
.A(n_1828),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_SL g2466 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2470)
);

INVx2_ASAP7_75t_SL g2471 ( 
.A(n_1486),
.Y(n_2471)
);

OAI221xp5_ASAP7_75t_L g2472 ( 
.A1(n_1309),
.A2(n_1196),
.B1(n_567),
.B2(n_763),
.C(n_685),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_L g2473 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2473)
);

AOI22xp33_ASAP7_75t_L g2474 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_L g2475 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2478)
);

INVxp67_ASAP7_75t_L g2479 ( 
.A(n_1686),
.Y(n_2479)
);

INVxp67_ASAP7_75t_SL g2480 ( 
.A(n_1431),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2482)
);

AOI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_1277),
.Y(n_2484)
);

INVx4_ASAP7_75t_L g2485 ( 
.A(n_1828),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_SL g2487 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_1277),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_1277),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_1457),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_1277),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2497)
);

O2A1O1Ixp5_ASAP7_75t_L g2498 ( 
.A1(n_1319),
.A2(n_1128),
.B(n_840),
.C(n_1081),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_1457),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_1277),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2501)
);

NOR2xp33_ASAP7_75t_SL g2502 ( 
.A(n_1745),
.B(n_716),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_SL g2506 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_1457),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_L g2510 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_1277),
.Y(n_2514)
);

AND2x6_ASAP7_75t_SL g2515 ( 
.A(n_1313),
.B(n_625),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_SL g2516 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_1457),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2520)
);

BUFx3_ASAP7_75t_L g2521 ( 
.A(n_1486),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2522)
);

NOR2xp33_ASAP7_75t_L g2523 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2523)
);

NOR2x1p5_ASAP7_75t_L g2524 ( 
.A(n_1681),
.B(n_405),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_1277),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2526)
);

AOI22xp33_ASAP7_75t_SL g2527 ( 
.A1(n_1309),
.A2(n_1275),
.B1(n_1770),
.B2(n_1672),
.Y(n_2527)
);

OAI221xp5_ASAP7_75t_L g2528 ( 
.A1(n_1309),
.A2(n_1196),
.B1(n_567),
.B2(n_763),
.C(n_685),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1277),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2530)
);

AOI22xp33_ASAP7_75t_L g2531 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_1277),
.Y(n_2533)
);

AOI22xp33_ASAP7_75t_L g2534 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2534)
);

NAND2xp33_ASAP7_75t_L g2535 ( 
.A(n_1314),
.B(n_1382),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2536)
);

NAND2xp33_ASAP7_75t_L g2537 ( 
.A(n_1314),
.B(n_1382),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_1277),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2542)
);

OAI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2546)
);

BUFx3_ASAP7_75t_L g2547 ( 
.A(n_1486),
.Y(n_2547)
);

AOI22xp33_ASAP7_75t_L g2548 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_1457),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_1457),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_L g2554 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_1457),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2556)
);

AND2x6_ASAP7_75t_SL g2557 ( 
.A(n_1313),
.B(n_625),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_SL g2558 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2559)
);

AND2x6_ASAP7_75t_L g2560 ( 
.A(n_1451),
.B(n_931),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_1277),
.Y(n_2561)
);

AOI22xp33_ASAP7_75t_L g2562 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2562)
);

AOI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2565)
);

A2O1A1Ixp33_ASAP7_75t_L g2566 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_1277),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_1277),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2571)
);

AOI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_1303),
.A2(n_1995),
.B(n_1962),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1277),
.Y(n_2573)
);

INVxp67_ASAP7_75t_L g2574 ( 
.A(n_1686),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_1277),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_1277),
.Y(n_2576)
);

NAND2xp33_ASAP7_75t_L g2577 ( 
.A(n_1314),
.B(n_1382),
.Y(n_2577)
);

NOR2xp67_ASAP7_75t_L g2578 ( 
.A(n_1349),
.B(n_716),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_1277),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_1457),
.Y(n_2580)
);

OAI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_2581)
);

CKINVDCx5p33_ASAP7_75t_R g2582 ( 
.A(n_1633),
.Y(n_2582)
);

INVx3_ASAP7_75t_L g2583 ( 
.A(n_1533),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2584)
);

AND3x1_ASAP7_75t_L g2585 ( 
.A(n_1309),
.B(n_924),
.C(n_1170),
.Y(n_2585)
);

AOI22xp5_ASAP7_75t_L g2586 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_1457),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_1457),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_L g2591 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2592)
);

BUFx6f_ASAP7_75t_SL g2593 ( 
.A(n_1384),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_1457),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_1277),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2597)
);

AND2x6_ASAP7_75t_L g2598 ( 
.A(n_1451),
.B(n_931),
.Y(n_2598)
);

A2O1A1Ixp33_ASAP7_75t_L g2599 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_1277),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_1277),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_SL g2603 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_1457),
.Y(n_2604)
);

A2O1A1Ixp33_ASAP7_75t_L g2605 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_2605)
);

AOI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_1457),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_1457),
.Y(n_2608)
);

INVx1_ASAP7_75t_SL g2609 ( 
.A(n_1279),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_1277),
.Y(n_2610)
);

O2A1O1Ixp5_ASAP7_75t_L g2611 ( 
.A1(n_1319),
.A2(n_1128),
.B(n_840),
.C(n_1081),
.Y(n_2611)
);

OAI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_1431),
.A2(n_1314),
.B1(n_1415),
.B2(n_1382),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_1277),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2615)
);

OR2x2_ASAP7_75t_L g2616 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2617)
);

A2O1A1Ixp33_ASAP7_75t_L g2618 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_1277),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2621)
);

AOI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2622)
);

INVx4_ASAP7_75t_L g2623 ( 
.A(n_1828),
.Y(n_2623)
);

OAI22xp5_ASAP7_75t_SL g2624 ( 
.A1(n_1380),
.A2(n_1196),
.B1(n_685),
.B2(n_763),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_SL g2626 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_1457),
.Y(n_2628)
);

OAI22xp33_ASAP7_75t_L g2629 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_2629)
);

BUFx3_ASAP7_75t_L g2630 ( 
.A(n_1486),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2631)
);

INVx5_ASAP7_75t_L g2632 ( 
.A(n_1533),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_1457),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_1277),
.Y(n_2634)
);

O2A1O1Ixp33_ASAP7_75t_L g2635 ( 
.A1(n_1326),
.A2(n_1128),
.B(n_747),
.C(n_750),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_1277),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_1277),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_SL g2641 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_SL g2642 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_1457),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_1457),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_1277),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_1277),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_SL g2652 ( 
.A(n_1745),
.B(n_716),
.Y(n_2652)
);

INVxp67_ASAP7_75t_SL g2653 ( 
.A(n_1431),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_1457),
.Y(n_2654)
);

INVx3_ASAP7_75t_L g2655 ( 
.A(n_1533),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_1533),
.Y(n_2656)
);

OAI22xp33_ASAP7_75t_L g2657 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_1277),
.Y(n_2659)
);

OAI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_2660)
);

BUFx3_ASAP7_75t_L g2661 ( 
.A(n_1486),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_1277),
.Y(n_2662)
);

AOI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_1303),
.A2(n_1995),
.B(n_1962),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_SL g2665 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_SL g2666 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_1457),
.Y(n_2667)
);

NOR2xp33_ASAP7_75t_L g2668 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2672)
);

BUFx8_ASAP7_75t_L g2673 ( 
.A(n_1640),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_1277),
.Y(n_2674)
);

BUFx2_ASAP7_75t_L g2675 ( 
.A(n_1343),
.Y(n_2675)
);

AOI221xp5_ASAP7_75t_L g2676 ( 
.A1(n_1309),
.A2(n_567),
.B1(n_1701),
.B2(n_1671),
.C(n_1276),
.Y(n_2676)
);

INVx4_ASAP7_75t_L g2677 ( 
.A(n_1828),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_1277),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2680)
);

BUFx6f_ASAP7_75t_L g2681 ( 
.A(n_1533),
.Y(n_2681)
);

AOI22xp33_ASAP7_75t_L g2682 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_1277),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2684)
);

O2A1O1Ixp33_ASAP7_75t_L g2685 ( 
.A1(n_1326),
.A2(n_1128),
.B(n_747),
.C(n_750),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_1277),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_1457),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_SL g2691 ( 
.A(n_1745),
.B(n_716),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_1277),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2694)
);

OAI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_2695)
);

NOR2xp33_ASAP7_75t_L g2696 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2697)
);

NAND3xp33_ASAP7_75t_L g2698 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2698)
);

AOI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_L g2701 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2701)
);

AOI22xp33_ASAP7_75t_L g2702 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_1277),
.Y(n_2703)
);

BUFx3_ASAP7_75t_L g2704 ( 
.A(n_1486),
.Y(n_2704)
);

INVx2_ASAP7_75t_SL g2705 ( 
.A(n_1486),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2706)
);

AOI21x1_ASAP7_75t_L g2707 ( 
.A1(n_1451),
.A2(n_1042),
.B(n_1532),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_1584),
.B(n_1318),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_1457),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_1457),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2714)
);

INVx2_ASAP7_75t_SL g2715 ( 
.A(n_1486),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2716)
);

BUFx3_ASAP7_75t_L g2717 ( 
.A(n_1486),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2718)
);

AOI22xp33_ASAP7_75t_L g2719 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2720)
);

NOR2xp33_ASAP7_75t_L g2721 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2722)
);

INVxp33_ASAP7_75t_L g2723 ( 
.A(n_1313),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_1633),
.Y(n_2724)
);

AND2x4_ASAP7_75t_L g2725 ( 
.A(n_1584),
.B(n_1318),
.Y(n_2725)
);

AOI22xp33_ASAP7_75t_L g2726 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_1457),
.Y(n_2727)
);

AOI221xp5_ASAP7_75t_L g2728 ( 
.A1(n_1309),
.A2(n_567),
.B1(n_1701),
.B2(n_1671),
.C(n_1276),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_SL g2729 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_1533),
.Y(n_2730)
);

INVx4_ASAP7_75t_L g2731 ( 
.A(n_1828),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_SL g2732 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_SL g2734 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_1277),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_1277),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_SL g2741 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2741)
);

NOR3xp33_ASAP7_75t_L g2742 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2742)
);

OAI22xp5_ASAP7_75t_SL g2743 ( 
.A1(n_1380),
.A2(n_1196),
.B1(n_685),
.B2(n_763),
.Y(n_2743)
);

BUFx6f_ASAP7_75t_L g2744 ( 
.A(n_1533),
.Y(n_2744)
);

O2A1O1Ixp33_ASAP7_75t_L g2745 ( 
.A1(n_1326),
.A2(n_1128),
.B(n_747),
.C(n_750),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2746)
);

A2O1A1Ixp33_ASAP7_75t_L g2747 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_2747)
);

AND2x4_ASAP7_75t_L g2748 ( 
.A(n_1584),
.B(n_1318),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_1277),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_1277),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_SL g2752 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2752)
);

OR2x2_ASAP7_75t_L g2753 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2753)
);

AOI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2754)
);

O2A1O1Ixp33_ASAP7_75t_L g2755 ( 
.A1(n_1326),
.A2(n_1128),
.B(n_747),
.C(n_750),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_1277),
.Y(n_2756)
);

NOR3xp33_ASAP7_75t_L g2757 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2761)
);

AOI22xp33_ASAP7_75t_L g2762 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_1277),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2766)
);

NOR3xp33_ASAP7_75t_L g2767 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2767)
);

INVxp33_ASAP7_75t_L g2768 ( 
.A(n_1313),
.Y(n_2768)
);

INVx2_ASAP7_75t_SL g2769 ( 
.A(n_1486),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2773)
);

BUFx3_ASAP7_75t_L g2774 ( 
.A(n_1486),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2777)
);

OAI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_SL g2780 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2782)
);

O2A1O1Ixp5_ASAP7_75t_L g2783 ( 
.A1(n_1319),
.A2(n_1128),
.B(n_840),
.C(n_1081),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2784)
);

NOR2xp33_ASAP7_75t_L g2785 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_1277),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_1457),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_1457),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_1457),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_1277),
.Y(n_2796)
);

AOI22xp33_ASAP7_75t_L g2797 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2798)
);

NAND2xp5_ASAP7_75t_L g2799 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2799)
);

NOR2xp33_ASAP7_75t_R g2800 ( 
.A(n_1490),
.B(n_716),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_1457),
.Y(n_2801)
);

INVx2_ASAP7_75t_SL g2802 ( 
.A(n_1486),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_SL g2803 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2803)
);

AOI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2804)
);

NAND3xp33_ASAP7_75t_L g2805 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2807)
);

A2O1A1Ixp33_ASAP7_75t_L g2808 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_1457),
.Y(n_2809)
);

INVxp67_ASAP7_75t_L g2810 ( 
.A(n_1686),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2811)
);

INVx2_ASAP7_75t_SL g2812 ( 
.A(n_1486),
.Y(n_2812)
);

AOI22xp33_ASAP7_75t_L g2813 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2814)
);

OR2x6_ASAP7_75t_L g2815 ( 
.A(n_1533),
.B(n_1129),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2818)
);

BUFx3_ASAP7_75t_L g2819 ( 
.A(n_1486),
.Y(n_2819)
);

INVx3_ASAP7_75t_L g2820 ( 
.A(n_1533),
.Y(n_2820)
);

INVx2_ASAP7_75t_SL g2821 ( 
.A(n_1486),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_SL g2822 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_1277),
.Y(n_2823)
);

NOR3xp33_ASAP7_75t_L g2824 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2825)
);

O2A1O1Ixp33_ASAP7_75t_L g2826 ( 
.A1(n_1326),
.A2(n_1128),
.B(n_747),
.C(n_750),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_1457),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_1277),
.Y(n_2828)
);

AOI221xp5_ASAP7_75t_L g2829 ( 
.A1(n_1309),
.A2(n_567),
.B1(n_1701),
.B2(n_1671),
.C(n_1276),
.Y(n_2829)
);

AOI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_1277),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_SL g2834 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2834)
);

AOI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_1303),
.A2(n_1995),
.B(n_1962),
.Y(n_2835)
);

AOI22xp33_ASAP7_75t_L g2836 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_1457),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_SL g2838 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_SL g2839 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2840)
);

NOR2xp33_ASAP7_75t_L g2841 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_SL g2843 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_1277),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_1457),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_SL g2846 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_SL g2848 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2848)
);

O2A1O1Ixp5_ASAP7_75t_L g2849 ( 
.A1(n_1319),
.A2(n_1128),
.B(n_840),
.C(n_1081),
.Y(n_2849)
);

INVx2_ASAP7_75t_SL g2850 ( 
.A(n_1486),
.Y(n_2850)
);

INVxp67_ASAP7_75t_SL g2851 ( 
.A(n_1431),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_SL g2853 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2853)
);

BUFx6f_ASAP7_75t_L g2854 ( 
.A(n_1533),
.Y(n_2854)
);

NOR2xp33_ASAP7_75t_L g2855 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2855)
);

OR2x6_ASAP7_75t_L g2856 ( 
.A(n_1533),
.B(n_1129),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_1303),
.A2(n_1995),
.B(n_1962),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_1457),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_1277),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2863)
);

OAI221xp5_ASAP7_75t_L g2864 ( 
.A1(n_1309),
.A2(n_1196),
.B1(n_567),
.B2(n_763),
.C(n_685),
.Y(n_2864)
);

BUFx3_ASAP7_75t_L g2865 ( 
.A(n_1486),
.Y(n_2865)
);

NOR2xp33_ASAP7_75t_L g2866 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2866)
);

OAI22x1_ASAP7_75t_SL g2867 ( 
.A1(n_1633),
.A2(n_1691),
.B1(n_1697),
.B2(n_1664),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2868)
);

AND2x4_ASAP7_75t_SL g2869 ( 
.A(n_1641),
.B(n_1095),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_1486),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_1457),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_1457),
.Y(n_2872)
);

BUFx6f_ASAP7_75t_SL g2873 ( 
.A(n_1384),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_1457),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2875)
);

NAND2xp33_ASAP7_75t_L g2876 ( 
.A(n_1314),
.B(n_1382),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_1457),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_SL g2879 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2879)
);

OR2x6_ASAP7_75t_L g2880 ( 
.A(n_1533),
.B(n_1129),
.Y(n_2880)
);

NOR2xp33_ASAP7_75t_L g2881 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_1277),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2884)
);

OAI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_1431),
.A2(n_1314),
.B1(n_1415),
.B2(n_1382),
.Y(n_2885)
);

AOI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2886)
);

NAND2xp33_ASAP7_75t_L g2887 ( 
.A(n_1314),
.B(n_1382),
.Y(n_2887)
);

AOI22xp33_ASAP7_75t_L g2888 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2890)
);

OR2x2_ASAP7_75t_L g2891 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2894)
);

INVx2_ASAP7_75t_SL g2895 ( 
.A(n_1486),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2897)
);

AND2x6_ASAP7_75t_SL g2898 ( 
.A(n_1313),
.B(n_625),
.Y(n_2898)
);

NOR3xp33_ASAP7_75t_L g2899 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2899)
);

AND2x4_ASAP7_75t_L g2900 ( 
.A(n_1584),
.B(n_1318),
.Y(n_2900)
);

NAND3xp33_ASAP7_75t_L g2901 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_1277),
.Y(n_2902)
);

BUFx6f_ASAP7_75t_L g2903 ( 
.A(n_1533),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_1277),
.Y(n_2905)
);

NOR3xp33_ASAP7_75t_L g2906 ( 
.A(n_1309),
.B(n_1081),
.C(n_814),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_SL g2907 ( 
.A(n_1745),
.B(n_716),
.Y(n_2907)
);

OR2x2_ASAP7_75t_L g2908 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_1277),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_1457),
.Y(n_2910)
);

AOI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2913)
);

OR2x2_ASAP7_75t_L g2914 ( 
.A(n_1686),
.B(n_1768),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_1457),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2916)
);

BUFx3_ASAP7_75t_L g2917 ( 
.A(n_1486),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2919)
);

AOI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2921)
);

AOI22xp33_ASAP7_75t_L g2922 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_2922)
);

AOI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2923)
);

OAI221xp5_ASAP7_75t_L g2924 ( 
.A1(n_1309),
.A2(n_1196),
.B1(n_567),
.B2(n_763),
.C(n_685),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_1457),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_1277),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2929)
);

INVxp67_ASAP7_75t_L g2930 ( 
.A(n_1686),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2931)
);

NOR2xp33_ASAP7_75t_L g2932 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_1457),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_1277),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2937)
);

AOI22xp5_ASAP7_75t_L g2938 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_SL g2939 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2939)
);

NOR2xp67_ASAP7_75t_SL g2940 ( 
.A(n_1724),
.B(n_407),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_1457),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_1745),
.B(n_1858),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2944)
);

OAI22xp5_ASAP7_75t_L g2945 ( 
.A1(n_1431),
.A2(n_1314),
.B1(n_1415),
.B2(n_1382),
.Y(n_2945)
);

INVxp67_ASAP7_75t_SL g2946 ( 
.A(n_1431),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_1457),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2948)
);

INVx2_ASAP7_75t_SL g2949 ( 
.A(n_1486),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2950)
);

AND2x2_ASAP7_75t_SL g2951 ( 
.A(n_2003),
.B(n_1275),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_1277),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_1277),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_1457),
.Y(n_2957)
);

OAI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_1431),
.A2(n_1128),
.B(n_840),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_1277),
.Y(n_2962)
);

BUFx3_ASAP7_75t_L g2963 ( 
.A(n_1486),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_1457),
.Y(n_2964)
);

INVx3_ASAP7_75t_L g2965 ( 
.A(n_1533),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2966)
);

NAND2xp33_ASAP7_75t_L g2967 ( 
.A(n_1314),
.B(n_1382),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2968)
);

NOR2xp33_ASAP7_75t_L g2969 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_1457),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_1457),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_1457),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_L g2975 ( 
.A(n_1309),
.B(n_1276),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_1457),
.Y(n_2977)
);

BUFx3_ASAP7_75t_L g2978 ( 
.A(n_1486),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_1290),
.B(n_1280),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2980)
);

INVxp67_ASAP7_75t_L g2981 ( 
.A(n_1686),
.Y(n_2981)
);

NAND2x1_ASAP7_75t_L g2982 ( 
.A(n_1576),
.B(n_1500),
.Y(n_2982)
);

OR2x2_ASAP7_75t_SL g2983 ( 
.A(n_1724),
.B(n_1855),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_1457),
.Y(n_2984)
);

INVx2_ASAP7_75t_SL g2985 ( 
.A(n_1486),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_SL g2988 ( 
.A(n_1650),
.B(n_1754),
.Y(n_2988)
);

OAI22xp5_ASAP7_75t_L g2989 ( 
.A1(n_1431),
.A2(n_1314),
.B1(n_1415),
.B2(n_1382),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_1457),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_1277),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_1277),
.Y(n_2993)
);

AND2x4_ASAP7_75t_L g2994 ( 
.A(n_1584),
.B(n_1318),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_1431),
.B(n_1364),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_1457),
.Y(n_2996)
);

OAI221xp5_ASAP7_75t_L g2997 ( 
.A1(n_1309),
.A2(n_1196),
.B1(n_567),
.B2(n_763),
.C(n_685),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_1277),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_1277),
.Y(n_2999)
);

OAI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_1431),
.A2(n_1314),
.B1(n_1415),
.B2(n_1382),
.Y(n_3000)
);

O2A1O1Ixp33_ASAP7_75t_L g3001 ( 
.A1(n_1326),
.A2(n_1128),
.B(n_747),
.C(n_750),
.Y(n_3001)
);

NOR2xp33_ASAP7_75t_L g3002 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_SL g3003 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3003)
);

AOI22xp33_ASAP7_75t_L g3004 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3006)
);

AOI22xp33_ASAP7_75t_L g3007 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_1277),
.Y(n_3008)
);

INVxp67_ASAP7_75t_SL g3009 ( 
.A(n_1431),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_1277),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_L g3014 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3015)
);

AOI22xp33_ASAP7_75t_L g3016 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3016)
);

OR2x6_ASAP7_75t_L g3017 ( 
.A(n_1533),
.B(n_1129),
.Y(n_3017)
);

NAND2xp33_ASAP7_75t_L g3018 ( 
.A(n_1314),
.B(n_1382),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_1457),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_1457),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3024)
);

AOI22xp33_ASAP7_75t_L g3025 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_1277),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_1457),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_1457),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_SL g3030 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3030)
);

CKINVDCx11_ASAP7_75t_R g3031 ( 
.A(n_1325),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_1277),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_SL g3034 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3034)
);

OAI22xp33_ASAP7_75t_L g3035 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_3035)
);

BUFx3_ASAP7_75t_L g3036 ( 
.A(n_1486),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_1457),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_L g3038 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3038)
);

AND2x6_ASAP7_75t_SL g3039 ( 
.A(n_1313),
.B(n_625),
.Y(n_3039)
);

AOI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_SL g3041 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3041)
);

NOR2x1p5_ASAP7_75t_L g3042 ( 
.A(n_1681),
.B(n_405),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_1457),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_1457),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_1277),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_1277),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_1277),
.Y(n_3048)
);

BUFx8_ASAP7_75t_L g3049 ( 
.A(n_1640),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_1290),
.B(n_1280),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_1277),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3052)
);

AO221x1_ASAP7_75t_L g3053 ( 
.A1(n_1292),
.A2(n_763),
.B1(n_685),
.B2(n_395),
.C(n_1056),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3054)
);

INVx8_ASAP7_75t_L g3055 ( 
.A(n_1828),
.Y(n_3055)
);

INVx1_ASAP7_75t_SL g3056 ( 
.A(n_1279),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_1457),
.Y(n_3057)
);

AND2x4_ASAP7_75t_L g3058 ( 
.A(n_1584),
.B(n_1318),
.Y(n_3058)
);

INVx3_ASAP7_75t_L g3059 ( 
.A(n_1533),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_1277),
.Y(n_3061)
);

OR2x2_ASAP7_75t_L g3062 ( 
.A(n_1686),
.B(n_1768),
.Y(n_3062)
);

INVx2_ASAP7_75t_SL g3063 ( 
.A(n_1486),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_1277),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_1290),
.B(n_1280),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_1290),
.B(n_1280),
.Y(n_3067)
);

NOR2x1p5_ASAP7_75t_L g3068 ( 
.A(n_1681),
.B(n_405),
.Y(n_3068)
);

AOI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3069)
);

INVx2_ASAP7_75t_SL g3070 ( 
.A(n_1486),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_1277),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3076)
);

AOI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_1277),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_1277),
.Y(n_3079)
);

INVx2_ASAP7_75t_SL g3080 ( 
.A(n_1486),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3082)
);

AOI22xp5_ASAP7_75t_L g3083 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_SL g3085 ( 
.A(n_1745),
.B(n_716),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_SL g3087 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_SL g3088 ( 
.A(n_1745),
.B(n_716),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3089)
);

INVx4_ASAP7_75t_L g3090 ( 
.A(n_1828),
.Y(n_3090)
);

NAND2x1_ASAP7_75t_L g3091 ( 
.A(n_1576),
.B(n_1500),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3092)
);

INVxp67_ASAP7_75t_L g3093 ( 
.A(n_1686),
.Y(n_3093)
);

AND2x6_ASAP7_75t_L g3094 ( 
.A(n_1451),
.B(n_931),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_SL g3095 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_L g3097 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_1457),
.Y(n_3099)
);

NOR2xp33_ASAP7_75t_L g3100 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_1457),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3102)
);

BUFx6f_ASAP7_75t_L g3103 ( 
.A(n_1533),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3104)
);

INVx3_ASAP7_75t_L g3105 ( 
.A(n_1533),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_SL g3107 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_1457),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3109)
);

A2O1A1Ixp33_ASAP7_75t_L g3110 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_L g3111 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_1277),
.Y(n_3112)
);

INVx5_ASAP7_75t_L g3113 ( 
.A(n_1533),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_1745),
.B(n_1858),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3117)
);

BUFx6f_ASAP7_75t_L g3118 ( 
.A(n_1533),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_1277),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_R g3121 ( 
.A(n_1490),
.B(n_716),
.Y(n_3121)
);

NAND2xp33_ASAP7_75t_SL g3122 ( 
.A(n_1558),
.B(n_613),
.Y(n_3122)
);

BUFx6f_ASAP7_75t_L g3123 ( 
.A(n_1533),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_SL g3125 ( 
.A(n_1745),
.B(n_1858),
.Y(n_3125)
);

AOI22xp33_ASAP7_75t_L g3126 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_1745),
.B(n_1858),
.Y(n_3127)
);

OAI221xp5_ASAP7_75t_L g3128 ( 
.A1(n_1309),
.A2(n_1196),
.B1(n_567),
.B2(n_763),
.C(n_685),
.Y(n_3128)
);

AOI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_SL g3130 ( 
.A(n_1745),
.B(n_1858),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_1290),
.B(n_1280),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_1457),
.Y(n_3132)
);

AND2x4_ASAP7_75t_L g3133 ( 
.A(n_1584),
.B(n_1318),
.Y(n_3133)
);

OAI22xp33_ASAP7_75t_L g3134 ( 
.A1(n_1314),
.A2(n_1415),
.B1(n_1421),
.B2(n_1382),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_L g3136 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3137)
);

INVx3_ASAP7_75t_L g3138 ( 
.A(n_1533),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_1277),
.Y(n_3142)
);

INVxp67_ASAP7_75t_SL g3143 ( 
.A(n_1431),
.Y(n_3143)
);

BUFx6f_ASAP7_75t_L g3144 ( 
.A(n_1533),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_SL g3145 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3146)
);

AOI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_1277),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_1457),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_1290),
.B(n_1280),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_1457),
.Y(n_3151)
);

AOI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_1290),
.B(n_1280),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_1277),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_1277),
.Y(n_3155)
);

NOR2x1p5_ASAP7_75t_L g3156 ( 
.A(n_1681),
.B(n_405),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3157)
);

INVx2_ASAP7_75t_SL g3158 ( 
.A(n_1486),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_1457),
.Y(n_3159)
);

BUFx8_ASAP7_75t_L g3160 ( 
.A(n_1640),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_1277),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_1290),
.B(n_1280),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_1457),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_SL g3166 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_1277),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_1457),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3171)
);

A2O1A1Ixp33_ASAP7_75t_L g3172 ( 
.A1(n_1431),
.A2(n_1369),
.B(n_1128),
.C(n_1276),
.Y(n_3172)
);

AND2x4_ASAP7_75t_L g3173 ( 
.A(n_1584),
.B(n_1318),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_1277),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3175)
);

NOR2xp33_ASAP7_75t_L g3176 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_SL g3178 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3178)
);

NAND2xp33_ASAP7_75t_SL g3179 ( 
.A(n_1558),
.B(n_613),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3180)
);

AOI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_1309),
.A2(n_867),
.B1(n_837),
.B2(n_1380),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_1457),
.Y(n_3182)
);

NOR2xp67_ASAP7_75t_L g3183 ( 
.A(n_1349),
.B(n_716),
.Y(n_3183)
);

AOI22xp33_ASAP7_75t_L g3184 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3185)
);

NAND2x1p5_ASAP7_75t_L g3186 ( 
.A(n_1576),
.B(n_1584),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_1457),
.Y(n_3189)
);

INVx4_ASAP7_75t_L g3190 ( 
.A(n_1828),
.Y(n_3190)
);

INVxp67_ASAP7_75t_L g3191 ( 
.A(n_1686),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_1457),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3193)
);

INVxp67_ASAP7_75t_L g3194 ( 
.A(n_1686),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_1277),
.Y(n_3198)
);

NOR2xp67_ASAP7_75t_L g3199 ( 
.A(n_1349),
.B(n_716),
.Y(n_3199)
);

AOI22xp33_ASAP7_75t_L g3200 ( 
.A1(n_1326),
.A2(n_1312),
.B1(n_1671),
.B2(n_1276),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_1457),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_1277),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_SL g3203 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_SL g3205 ( 
.A(n_1650),
.B(n_1754),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_1457),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_1277),
.Y(n_3208)
);

NOR2xp33_ASAP7_75t_L g3209 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_L g3210 ( 
.A(n_1309),
.B(n_1276),
.Y(n_3210)
);

OR2x2_ASAP7_75t_L g3211 ( 
.A(n_1686),
.B(n_1768),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_1457),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_1457),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_1277),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_1431),
.B(n_1364),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_1277),
.Y(n_3218)
);

BUFx6f_ASAP7_75t_L g3219 ( 
.A(n_2707),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2414),
.B(n_2433),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_2036),
.B(n_2011),
.Y(n_3221)
);

O2A1O1Ixp33_ASAP7_75t_L g3222 ( 
.A1(n_2018),
.A2(n_2566),
.B(n_2599),
.C(n_2428),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_SL g3223 ( 
.A(n_2543),
.B(n_2581),
.Y(n_3223)
);

A2O1A1Ixp33_ASAP7_75t_L g3224 ( 
.A1(n_2958),
.A2(n_2618),
.B(n_2747),
.C(n_2605),
.Y(n_3224)
);

AOI22xp33_ASAP7_75t_L g3225 ( 
.A1(n_2017),
.A2(n_2022),
.B1(n_2027),
.B2(n_2024),
.Y(n_3225)
);

NOR2xp33_ASAP7_75t_L g3226 ( 
.A(n_2011),
.B(n_2408),
.Y(n_3226)
);

NAND2x1p5_ASAP7_75t_L g3227 ( 
.A(n_2083),
.B(n_2081),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2091),
.Y(n_3228)
);

BUFx2_ASAP7_75t_L g3229 ( 
.A(n_2010),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2282),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_2543),
.B(n_2581),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_2808),
.B(n_3110),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2612),
.B(n_2885),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2945),
.B(n_2989),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2306),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_2408),
.B(n_2416),
.Y(n_3236)
);

INVx2_ASAP7_75t_SL g3237 ( 
.A(n_2381),
.Y(n_3237)
);

OAI22xp33_ASAP7_75t_L g3238 ( 
.A1(n_2035),
.A2(n_2622),
.B1(n_2699),
.B2(n_2586),
.Y(n_3238)
);

BUFx6f_ASAP7_75t_L g3239 ( 
.A(n_2388),
.Y(n_3239)
);

BUFx3_ASAP7_75t_L g3240 ( 
.A(n_2175),
.Y(n_3240)
);

BUFx6f_ASAP7_75t_L g3241 ( 
.A(n_2359),
.Y(n_3241)
);

HB1xp67_ASAP7_75t_L g3242 ( 
.A(n_2292),
.Y(n_3242)
);

AOI22xp5_ASAP7_75t_L g3243 ( 
.A1(n_2416),
.A2(n_2473),
.B1(n_2481),
.B2(n_2454),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3000),
.B(n_2629),
.Y(n_3244)
);

BUFx3_ASAP7_75t_L g3245 ( 
.A(n_2175),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2629),
.B(n_2657),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2020),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_SL g3248 ( 
.A(n_2657),
.B(n_2660),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2660),
.B(n_2695),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2021),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_2454),
.B(n_2473),
.Y(n_3251)
);

NOR2xp33_ASAP7_75t_L g3252 ( 
.A(n_2481),
.B(n_2482),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_2560),
.Y(n_3253)
);

INVx3_ASAP7_75t_L g3254 ( 
.A(n_2310),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2695),
.B(n_2778),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2778),
.B(n_3035),
.Y(n_3256)
);

A2O1A1Ixp33_ASAP7_75t_L g3257 ( 
.A1(n_3172),
.A2(n_2017),
.B(n_2024),
.C(n_2022),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2031),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3035),
.B(n_3134),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2125),
.Y(n_3260)
);

NOR2xp33_ASAP7_75t_L g3261 ( 
.A(n_2482),
.B(n_2504),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2040),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3134),
.B(n_2043),
.Y(n_3263)
);

AOI22xp33_ASAP7_75t_L g3264 ( 
.A1(n_2027),
.A2(n_2510),
.B1(n_2517),
.B2(n_2504),
.Y(n_3264)
);

NAND3xp33_ASAP7_75t_SL g3265 ( 
.A(n_2676),
.B(n_2829),
.C(n_2728),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2025),
.B(n_2023),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_2125),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_2083),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_2423),
.B(n_2474),
.Y(n_3269)
);

INVx4_ASAP7_75t_L g3270 ( 
.A(n_2310),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2055),
.Y(n_3271)
);

BUFx2_ASAP7_75t_L g3272 ( 
.A(n_2090),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2075),
.Y(n_3273)
);

INVx3_ASAP7_75t_L g3274 ( 
.A(n_2310),
.Y(n_3274)
);

OAI21xp33_ASAP7_75t_L g3275 ( 
.A1(n_3210),
.A2(n_2517),
.B(n_2510),
.Y(n_3275)
);

AOI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_2518),
.A2(n_2554),
.B1(n_2564),
.B2(n_2523),
.Y(n_3276)
);

INVx2_ASAP7_75t_SL g3277 ( 
.A(n_2982),
.Y(n_3277)
);

INVxp67_ASAP7_75t_SL g3278 ( 
.A(n_2299),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2030),
.B(n_2034),
.Y(n_3279)
);

OAI22xp5_ASAP7_75t_L g3280 ( 
.A1(n_2009),
.A2(n_2407),
.B1(n_2411),
.B2(n_2410),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2077),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2111),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2518),
.B(n_2523),
.Y(n_3283)
);

INVx5_ASAP7_75t_L g3284 ( 
.A(n_2310),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2038),
.B(n_2423),
.Y(n_3285)
);

INVx2_ASAP7_75t_L g3286 ( 
.A(n_2106),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_SL g3287 ( 
.A(n_2474),
.B(n_2483),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2124),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_SL g3289 ( 
.A(n_2483),
.B(n_2531),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_2013),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2531),
.B(n_2534),
.Y(n_3291)
);

BUFx2_ASAP7_75t_L g3292 ( 
.A(n_2560),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_2534),
.B(n_2548),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2126),
.Y(n_3294)
);

BUFx6f_ASAP7_75t_L g3295 ( 
.A(n_3094),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_2013),
.Y(n_3296)
);

NAND2x1p5_ASAP7_75t_L g3297 ( 
.A(n_2081),
.B(n_2100),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2127),
.Y(n_3298)
);

OAI22xp5_ASAP7_75t_L g3299 ( 
.A1(n_2426),
.A2(n_2435),
.B1(n_2440),
.B2(n_2427),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_SL g3300 ( 
.A(n_2548),
.B(n_2562),
.Y(n_3300)
);

AND2x4_ASAP7_75t_L g3301 ( 
.A(n_2143),
.B(n_2560),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_2441),
.A2(n_2446),
.B1(n_2449),
.B2(n_2443),
.Y(n_3302)
);

NAND2x1p5_ASAP7_75t_L g3303 ( 
.A(n_2100),
.B(n_2424),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_2562),
.B(n_2563),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_2563),
.B(n_2606),
.Y(n_3305)
);

NOR2xp33_ASAP7_75t_L g3306 ( 
.A(n_2554),
.B(n_2564),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2140),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_2606),
.B(n_2682),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_L g3309 ( 
.A(n_2591),
.B(n_2597),
.Y(n_3309)
);

AOI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_2572),
.A2(n_2835),
.B(n_2663),
.Y(n_3310)
);

HB1xp67_ASAP7_75t_L g3311 ( 
.A(n_2420),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_2141),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_2682),
.B(n_2702),
.Y(n_3313)
);

INVx4_ASAP7_75t_L g3314 ( 
.A(n_2310),
.Y(n_3314)
);

AOI22xp5_ASAP7_75t_L g3315 ( 
.A1(n_2591),
.A2(n_2597),
.B1(n_2668),
.B2(n_2664),
.Y(n_3315)
);

AOI22xp5_ASAP7_75t_L g3316 ( 
.A1(n_2664),
.A2(n_2668),
.B1(n_2696),
.B2(n_2669),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_L g3317 ( 
.A(n_2669),
.B(n_2696),
.Y(n_3317)
);

AOI22xp33_ASAP7_75t_L g3318 ( 
.A1(n_2701),
.A2(n_2736),
.B1(n_2760),
.B2(n_2721),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_L g3319 ( 
.A(n_2701),
.B(n_2721),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_2702),
.B(n_2713),
.Y(n_3320)
);

CKINVDCx5p33_ASAP7_75t_R g3321 ( 
.A(n_3031),
.Y(n_3321)
);

OAI22xp33_ASAP7_75t_L g3322 ( 
.A1(n_2754),
.A2(n_2830),
.B1(n_2886),
.B2(n_2781),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_2424),
.Y(n_3323)
);

AO22x1_ASAP7_75t_L g3324 ( 
.A1(n_2736),
.A2(n_2779),
.B1(n_2785),
.B2(n_2760),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2713),
.B(n_2719),
.Y(n_3325)
);

NOR2xp33_ASAP7_75t_L g3326 ( 
.A(n_2779),
.B(n_2785),
.Y(n_3326)
);

INVx2_ASAP7_75t_SL g3327 ( 
.A(n_3091),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2439),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_2818),
.A2(n_2855),
.B1(n_2866),
.B2(n_2841),
.Y(n_3329)
);

AOI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2818),
.A2(n_2855),
.B1(n_2866),
.B2(n_2841),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2144),
.Y(n_3331)
);

BUFx2_ASAP7_75t_L g3332 ( 
.A(n_2560),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_2439),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2719),
.B(n_2726),
.Y(n_3334)
);

AOI22xp5_ASAP7_75t_L g3335 ( 
.A1(n_2881),
.A2(n_2894),
.B1(n_2897),
.B2(n_2893),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2726),
.B(n_2762),
.Y(n_3336)
);

AND2x6_ASAP7_75t_SL g3337 ( 
.A(n_2881),
.B(n_2893),
.Y(n_3337)
);

INVx1_ASAP7_75t_L g3338 ( 
.A(n_2146),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2168),
.Y(n_3339)
);

INVx2_ASAP7_75t_SL g3340 ( 
.A(n_2339),
.Y(n_3340)
);

AOI22xp5_ASAP7_75t_L g3341 ( 
.A1(n_2894),
.A2(n_2913),
.B1(n_2916),
.B2(n_2897),
.Y(n_3341)
);

INVx2_ASAP7_75t_SL g3342 ( 
.A(n_2339),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2179),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_2913),
.B(n_2916),
.Y(n_3344)
);

INVx3_ASAP7_75t_L g3345 ( 
.A(n_2560),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2185),
.Y(n_3346)
);

OR2x2_ASAP7_75t_SL g3347 ( 
.A(n_2698),
.B(n_2805),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_2762),
.B(n_2797),
.Y(n_3348)
);

BUFx6f_ASAP7_75t_L g3349 ( 
.A(n_2598),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2797),
.B(n_2804),
.Y(n_3350)
);

INVx3_ASAP7_75t_L g3351 ( 
.A(n_2598),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_2804),
.B(n_2813),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_SL g3353 ( 
.A(n_2813),
.B(n_2836),
.Y(n_3353)
);

AOI22xp33_ASAP7_75t_L g3354 ( 
.A1(n_2931),
.A2(n_2956),
.B1(n_2959),
.B2(n_2932),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_2836),
.B(n_2842),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2188),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2195),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_2931),
.B(n_2932),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_2956),
.A2(n_2968),
.B1(n_2969),
.B2(n_2959),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_SL g3360 ( 
.A1(n_2968),
.A2(n_3038),
.B1(n_3210),
.B2(n_2969),
.Y(n_3360)
);

INVx2_ASAP7_75t_SL g3361 ( 
.A(n_2086),
.Y(n_3361)
);

AOI22xp5_ASAP7_75t_L g3362 ( 
.A1(n_2975),
.A2(n_3014),
.B1(n_3015),
.B2(n_3002),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_2444),
.Y(n_3363)
);

BUFx6f_ASAP7_75t_SL g3364 ( 
.A(n_2598),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_2842),
.B(n_2888),
.Y(n_3365)
);

AO22x1_ASAP7_75t_L g3366 ( 
.A1(n_2975),
.A2(n_3014),
.B1(n_3015),
.B2(n_3002),
.Y(n_3366)
);

INVx2_ASAP7_75t_SL g3367 ( 
.A(n_2598),
.Y(n_3367)
);

NOR2xp33_ASAP7_75t_L g3368 ( 
.A(n_3022),
.B(n_3038),
.Y(n_3368)
);

INVx2_ASAP7_75t_L g3369 ( 
.A(n_2444),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_3022),
.B(n_3096),
.Y(n_3370)
);

BUFx6f_ASAP7_75t_L g3371 ( 
.A(n_2598),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_3096),
.B(n_3097),
.Y(n_3372)
);

INVx3_ASAP7_75t_L g3373 ( 
.A(n_3094),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2197),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_2888),
.B(n_2922),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_SL g3376 ( 
.A1(n_3176),
.A2(n_3209),
.B1(n_3193),
.B2(n_3100),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_2922),
.B(n_3004),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3004),
.B(n_3006),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3006),
.B(n_3007),
.Y(n_3379)
);

INVx4_ASAP7_75t_L g3380 ( 
.A(n_2632),
.Y(n_3380)
);

AND2x4_ASAP7_75t_L g3381 ( 
.A(n_2143),
.B(n_3094),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_3097),
.B(n_3100),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3007),
.B(n_3016),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_3016),
.B(n_3025),
.Y(n_3384)
);

NOR2x1_ASAP7_75t_R g3385 ( 
.A(n_2142),
.B(n_2041),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_2466),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2204),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_3025),
.B(n_3069),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_2466),
.Y(n_3389)
);

AND3x2_ASAP7_75t_SL g3390 ( 
.A(n_2119),
.B(n_3126),
.C(n_3069),
.Y(n_3390)
);

AOI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3102),
.A2(n_3136),
.B1(n_3170),
.B2(n_3111),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3126),
.B(n_3147),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3147),
.B(n_3184),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_2234),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_2240),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_2470),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_2470),
.Y(n_3397)
);

AND2x4_ASAP7_75t_L g3398 ( 
.A(n_3094),
.B(n_2050),
.Y(n_3398)
);

BUFx2_ASAP7_75t_L g3399 ( 
.A(n_3094),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2251),
.Y(n_3400)
);

NAND3xp33_ASAP7_75t_SL g3401 ( 
.A(n_2911),
.B(n_2923),
.C(n_2920),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3184),
.B(n_3200),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3200),
.B(n_2048),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2254),
.Y(n_3404)
);

BUFx6f_ASAP7_75t_L g3405 ( 
.A(n_2478),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_2478),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2261),
.Y(n_3407)
);

INVx3_ASAP7_75t_L g3408 ( 
.A(n_2632),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_2859),
.A2(n_2491),
.B(n_2487),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_2062),
.B(n_2119),
.Y(n_3410)
);

INVx4_ASAP7_75t_L g3411 ( 
.A(n_2632),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2262),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2272),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_3102),
.B(n_3111),
.Y(n_3414)
);

BUFx12f_ASAP7_75t_L g3415 ( 
.A(n_2042),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3136),
.B(n_3170),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_2278),
.Y(n_3417)
);

BUFx6f_ASAP7_75t_L g3418 ( 
.A(n_2487),
.Y(n_3418)
);

NOR2xp33_ASAP7_75t_L g3419 ( 
.A(n_3176),
.B(n_3180),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_2048),
.B(n_2450),
.Y(n_3420)
);

NOR2x2_ASAP7_75t_L g3421 ( 
.A(n_2199),
.B(n_2078),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2280),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_SL g3423 ( 
.A(n_2434),
.B(n_2475),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2461),
.B(n_2463),
.Y(n_3424)
);

CKINVDCx5p33_ASAP7_75t_R g3425 ( 
.A(n_2800),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_2491),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_2495),
.Y(n_3427)
);

BUFx6f_ASAP7_75t_L g3428 ( 
.A(n_2495),
.Y(n_3428)
);

AND2x4_ASAP7_75t_L g3429 ( 
.A(n_2050),
.B(n_2632),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_L g3430 ( 
.A(n_3180),
.B(n_3193),
.Y(n_3430)
);

INVx2_ASAP7_75t_SL g3431 ( 
.A(n_2276),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_2298),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_2305),
.Y(n_3433)
);

OR2x2_ASAP7_75t_L g3434 ( 
.A(n_2496),
.B(n_2501),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_2496),
.Y(n_3435)
);

A2O1A1Ixp33_ASAP7_75t_L g3436 ( 
.A1(n_3209),
.A2(n_3196),
.B(n_3195),
.C(n_2611),
.Y(n_3436)
);

HB1xp67_ASAP7_75t_L g3437 ( 
.A(n_2432),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_SL g3438 ( 
.A(n_2742),
.B(n_2757),
.Y(n_3438)
);

AND2x4_ASAP7_75t_L g3439 ( 
.A(n_3113),
.B(n_2019),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_SL g3440 ( 
.A(n_2767),
.B(n_2824),
.Y(n_3440)
);

NAND2x1p5_ASAP7_75t_L g3441 ( 
.A(n_2501),
.B(n_2503),
.Y(n_3441)
);

INVx3_ASAP7_75t_L g3442 ( 
.A(n_3113),
.Y(n_3442)
);

BUFx3_ASAP7_75t_L g3443 ( 
.A(n_2453),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_SL g3444 ( 
.A(n_2899),
.B(n_2906),
.Y(n_3444)
);

NOR2xp33_ASAP7_75t_L g3445 ( 
.A(n_3195),
.B(n_3196),
.Y(n_3445)
);

INVx3_ASAP7_75t_L g3446 ( 
.A(n_3113),
.Y(n_3446)
);

AOI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_2934),
.A2(n_3040),
.B1(n_3077),
.B2(n_2938),
.Y(n_3447)
);

INVx6_ASAP7_75t_L g3448 ( 
.A(n_3113),
.Y(n_3448)
);

BUFx2_ASAP7_75t_L g3449 ( 
.A(n_2085),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_2307),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_2464),
.B(n_2467),
.Y(n_3451)
);

CKINVDCx5p33_ASAP7_75t_R g3452 ( 
.A(n_2800),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2468),
.B(n_2469),
.Y(n_3453)
);

BUFx3_ASAP7_75t_L g3454 ( 
.A(n_2453),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_R g3455 ( 
.A(n_3122),
.B(n_3179),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_2311),
.Y(n_3456)
);

BUFx12f_ASAP7_75t_L g3457 ( 
.A(n_2042),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_2476),
.B(n_2477),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_SL g3459 ( 
.A(n_2057),
.B(n_2901),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_2019),
.B(n_2503),
.Y(n_3460)
);

INVxp67_ASAP7_75t_L g3461 ( 
.A(n_2120),
.Y(n_3461)
);

XOR2x2_ASAP7_75t_L g3462 ( 
.A(n_2624),
.B(n_2743),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_SL g3463 ( 
.A(n_2074),
.B(n_2486),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_2506),
.Y(n_3464)
);

AOI22x1_ASAP7_75t_L g3465 ( 
.A1(n_2480),
.A2(n_2653),
.B1(n_2946),
.B2(n_2851),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2324),
.Y(n_3466)
);

INVxp67_ASAP7_75t_SL g3467 ( 
.A(n_2327),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_2506),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_2488),
.B(n_2492),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_2409),
.Y(n_3470)
);

BUFx3_ASAP7_75t_L g3471 ( 
.A(n_2453),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_2511),
.Y(n_3472)
);

AOI21xp5_ASAP7_75t_L g3473 ( 
.A1(n_2511),
.A2(n_2536),
.B(n_2516),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_2412),
.Y(n_3474)
);

BUFx3_ASAP7_75t_L g3475 ( 
.A(n_2465),
.Y(n_3475)
);

AOI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_2516),
.A2(n_2538),
.B(n_2536),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_2497),
.B(n_2505),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_2538),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_2546),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_2546),
.Y(n_3480)
);

HB1xp67_ASAP7_75t_L g3481 ( 
.A(n_2551),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_2507),
.B(n_2509),
.Y(n_3482)
);

AOI22xp5_ASAP7_75t_L g3483 ( 
.A1(n_3083),
.A2(n_3129),
.B1(n_3152),
.B2(n_3098),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_R g3484 ( 
.A(n_2431),
.B(n_2502),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_SL g3485 ( 
.A(n_2513),
.B(n_2520),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_2551),
.A2(n_2569),
.B(n_2558),
.Y(n_3486)
);

CKINVDCx5p33_ASAP7_75t_R g3487 ( 
.A(n_3121),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_2522),
.B(n_2526),
.Y(n_3488)
);

AND2x4_ASAP7_75t_L g3489 ( 
.A(n_2174),
.B(n_2051),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2530),
.B(n_2539),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_2413),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_2417),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_L g3493 ( 
.A1(n_3053),
.A2(n_2528),
.B1(n_2864),
.B2(n_2472),
.Y(n_3493)
);

BUFx12f_ASAP7_75t_L g3494 ( 
.A(n_2673),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_SL g3495 ( 
.A(n_2541),
.B(n_2542),
.Y(n_3495)
);

NOR3xp33_ASAP7_75t_SL g3496 ( 
.A(n_2924),
.B(n_3128),
.C(n_2997),
.Y(n_3496)
);

OR2x2_ASAP7_75t_L g3497 ( 
.A(n_2558),
.B(n_2569),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_2544),
.B(n_2545),
.Y(n_3498)
);

BUFx2_ASAP7_75t_L g3499 ( 
.A(n_2199),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_2552),
.B(n_2553),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_2603),
.Y(n_3501)
);

AOI22xp33_ASAP7_75t_L g3502 ( 
.A1(n_3181),
.A2(n_3143),
.B1(n_3009),
.B2(n_2418),
.Y(n_3502)
);

BUFx12f_ASAP7_75t_L g3503 ( 
.A(n_2673),
.Y(n_3503)
);

CKINVDCx5p33_ASAP7_75t_R g3504 ( 
.A(n_3121),
.Y(n_3504)
);

NOR2xp33_ASAP7_75t_L g3505 ( 
.A(n_2723),
.B(n_2768),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_2419),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_2556),
.B(n_2559),
.Y(n_3507)
);

INVx3_ASAP7_75t_L g3508 ( 
.A(n_2029),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_2421),
.Y(n_3509)
);

AOI22xp33_ASAP7_75t_L g3510 ( 
.A1(n_2535),
.A2(n_2537),
.B1(n_2876),
.B2(n_2577),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_2567),
.B(n_2571),
.Y(n_3511)
);

INVx2_ASAP7_75t_SL g3512 ( 
.A(n_2276),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_2429),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_2603),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_2584),
.B(n_2587),
.Y(n_3515)
);

NAND3xp33_ASAP7_75t_L g3516 ( 
.A(n_2498),
.B(n_2849),
.C(n_2783),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_2588),
.B(n_2592),
.Y(n_3517)
);

AOI22xp5_ASAP7_75t_L g3518 ( 
.A1(n_2585),
.A2(n_2016),
.B1(n_2967),
.B2(n_2887),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_2617),
.Y(n_3519)
);

HB1xp67_ASAP7_75t_L g3520 ( 
.A(n_2617),
.Y(n_3520)
);

BUFx6f_ASAP7_75t_L g3521 ( 
.A(n_2621),
.Y(n_3521)
);

NAND3xp33_ASAP7_75t_SL g3522 ( 
.A(n_2448),
.B(n_2635),
.C(n_2456),
.Y(n_3522)
);

INVx3_ASAP7_75t_L g3523 ( 
.A(n_2029),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_2594),
.B(n_2602),
.Y(n_3524)
);

AND2x4_ASAP7_75t_L g3525 ( 
.A(n_2174),
.B(n_2051),
.Y(n_3525)
);

INVx4_ASAP7_75t_L g3526 ( 
.A(n_2436),
.Y(n_3526)
);

INVx4_ASAP7_75t_L g3527 ( 
.A(n_2436),
.Y(n_3527)
);

AOI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_2621),
.A2(n_2626),
.B(n_2625),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_2437),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_2614),
.B(n_2615),
.Y(n_3530)
);

BUFx6f_ASAP7_75t_L g3531 ( 
.A(n_2625),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_2626),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_2620),
.B(n_2645),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_2631),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_2447),
.Y(n_3535)
);

INVx4_ASAP7_75t_L g3536 ( 
.A(n_2436),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_2646),
.B(n_2647),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_L g3538 ( 
.A(n_2649),
.B(n_2658),
.Y(n_3538)
);

INVx5_ASAP7_75t_L g3539 ( 
.A(n_2078),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_2671),
.B(n_2679),
.Y(n_3540)
);

BUFx3_ASAP7_75t_L g3541 ( 
.A(n_2951),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_2684),
.B(n_2687),
.Y(n_3542)
);

AOI22xp5_ASAP7_75t_L g3543 ( 
.A1(n_3018),
.A2(n_2068),
.B1(n_2690),
.B2(n_2688),
.Y(n_3543)
);

INVx2_ASAP7_75t_SL g3544 ( 
.A(n_2283),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_2692),
.B(n_2694),
.Y(n_3545)
);

BUFx3_ASAP7_75t_L g3546 ( 
.A(n_2951),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_2457),
.Y(n_3547)
);

AND2x4_ASAP7_75t_SL g3548 ( 
.A(n_2078),
.B(n_2436),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_2631),
.Y(n_3549)
);

NAND2xp33_ASAP7_75t_SL g3550 ( 
.A(n_3213),
.B(n_3215),
.Y(n_3550)
);

NOR2x2_ASAP7_75t_L g3551 ( 
.A(n_2199),
.B(n_2399),
.Y(n_3551)
);

NOR2xp33_ASAP7_75t_L g3552 ( 
.A(n_2697),
.B(n_2700),
.Y(n_3552)
);

INVx3_ASAP7_75t_L g3553 ( 
.A(n_3186),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_2706),
.B(n_2709),
.Y(n_3554)
);

INVx2_ASAP7_75t_L g3555 ( 
.A(n_2636),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_SL g3556 ( 
.A(n_2710),
.B(n_2716),
.Y(n_3556)
);

OAI21xp5_ASAP7_75t_L g3557 ( 
.A1(n_2636),
.A2(n_3205),
.B(n_3203),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_2720),
.B(n_2722),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_2735),
.B(n_2738),
.Y(n_3559)
);

AOI22xp5_ASAP7_75t_L g3560 ( 
.A1(n_2739),
.A2(n_2746),
.B1(n_2761),
.B2(n_2758),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_2638),
.A2(n_2642),
.B(n_2641),
.Y(n_3561)
);

CKINVDCx5p33_ASAP7_75t_R g3562 ( 
.A(n_2348),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_2459),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_2763),
.B(n_2765),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_SL g3565 ( 
.A(n_2766),
.B(n_2770),
.Y(n_3565)
);

BUFx3_ASAP7_75t_L g3566 ( 
.A(n_2465),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_2638),
.A2(n_2642),
.B(n_2641),
.Y(n_3567)
);

AND2x4_ASAP7_75t_L g3568 ( 
.A(n_2708),
.B(n_2725),
.Y(n_3568)
);

INVxp67_ASAP7_75t_SL g3569 ( 
.A(n_2275),
.Y(n_3569)
);

OR2x2_ASAP7_75t_L g3570 ( 
.A(n_2665),
.B(n_2666),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_2771),
.B(n_2772),
.Y(n_3571)
);

OR2x6_ASAP7_75t_L g3572 ( 
.A(n_2665),
.B(n_2666),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_L g3573 ( 
.A(n_2775),
.B(n_2776),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_2777),
.B(n_2784),
.Y(n_3574)
);

AND2x2_ASAP7_75t_L g3575 ( 
.A(n_2672),
.B(n_2714),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_2484),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_2790),
.B(n_2792),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_2489),
.Y(n_3578)
);

BUFx2_ASAP7_75t_L g3579 ( 
.A(n_2490),
.Y(n_3579)
);

AOI22xp33_ASAP7_75t_L g3580 ( 
.A1(n_2672),
.A2(n_2718),
.B1(n_2729),
.B2(n_2714),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_2718),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_2494),
.Y(n_3582)
);

BUFx6f_ASAP7_75t_L g3583 ( 
.A(n_2729),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_2732),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3203),
.B(n_3205),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_2732),
.Y(n_3586)
);

INVx2_ASAP7_75t_L g3587 ( 
.A(n_2733),
.Y(n_3587)
);

INVxp67_ASAP7_75t_SL g3588 ( 
.A(n_2275),
.Y(n_3588)
);

AND2x2_ASAP7_75t_L g3589 ( 
.A(n_2733),
.B(n_2734),
.Y(n_3589)
);

INVx2_ASAP7_75t_SL g3590 ( 
.A(n_2283),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_2734),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_2795),
.B(n_2798),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_SL g3593 ( 
.A(n_2799),
.B(n_2806),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_2500),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_2514),
.Y(n_3595)
);

AOI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_2807),
.A2(n_2811),
.B1(n_2816),
.B2(n_2814),
.Y(n_3596)
);

CKINVDCx5p33_ASAP7_75t_R g3597 ( 
.A(n_2348),
.Y(n_3597)
);

OAI22xp33_ASAP7_75t_L g3598 ( 
.A1(n_2833),
.A2(n_2840),
.B1(n_2857),
.B2(n_2852),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_2525),
.Y(n_3599)
);

AOI22xp5_ASAP7_75t_L g3600 ( 
.A1(n_2858),
.A2(n_2863),
.B1(n_2883),
.B2(n_2877),
.Y(n_3600)
);

INVx1_ASAP7_75t_SL g3601 ( 
.A(n_2145),
.Y(n_3601)
);

BUFx4f_ASAP7_75t_L g3602 ( 
.A(n_2681),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_SL g3603 ( 
.A(n_2884),
.B(n_2890),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_2741),
.Y(n_3604)
);

BUFx3_ASAP7_75t_L g3605 ( 
.A(n_2983),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_2741),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_2896),
.B(n_2904),
.Y(n_3607)
);

NOR2x2_ASAP7_75t_L g3608 ( 
.A(n_2399),
.B(n_2264),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_2912),
.B(n_2918),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_2529),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_2533),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_2750),
.Y(n_3612)
);

OR2x6_ASAP7_75t_L g3613 ( 
.A(n_2750),
.B(n_2752),
.Y(n_3613)
);

AOI22xp33_ASAP7_75t_L g3614 ( 
.A1(n_2752),
.A2(n_2773),
.B1(n_2780),
.B2(n_2759),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_2540),
.Y(n_3615)
);

A2O1A1Ixp33_ASAP7_75t_L g3616 ( 
.A1(n_2685),
.A2(n_2755),
.B(n_2826),
.C(n_2745),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_2759),
.A2(n_2780),
.B(n_2773),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_2782),
.A2(n_2793),
.B(n_2787),
.Y(n_3618)
);

AND2x4_ASAP7_75t_L g3619 ( 
.A(n_2708),
.B(n_2725),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_2561),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_SL g3621 ( 
.A(n_2925),
.B(n_2926),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_SL g3622 ( 
.A(n_2929),
.B(n_2937),
.Y(n_3622)
);

OR2x4_ASAP7_75t_L g3623 ( 
.A(n_2255),
.B(n_2148),
.Y(n_3623)
);

A2O1A1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_3001),
.A2(n_2948),
.B(n_2952),
.C(n_2944),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_2966),
.B(n_2970),
.Y(n_3625)
);

BUFx8_ASAP7_75t_L g3626 ( 
.A(n_2593),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_2782),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_2973),
.B(n_2976),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_2980),
.B(n_2986),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_2568),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_2987),
.B(n_2990),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_L g3632 ( 
.A(n_2995),
.B(n_3005),
.Y(n_3632)
);

CKINVDCx5p33_ASAP7_75t_R g3633 ( 
.A(n_2285),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_2787),
.B(n_2793),
.Y(n_3634)
);

AOI22xp5_ASAP7_75t_L g3635 ( 
.A1(n_3010),
.A2(n_3011),
.B1(n_3019),
.B2(n_3013),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_2570),
.Y(n_3636)
);

INVx5_ASAP7_75t_L g3637 ( 
.A(n_2151),
.Y(n_3637)
);

AND2x4_ASAP7_75t_L g3638 ( 
.A(n_2748),
.B(n_2900),
.Y(n_3638)
);

HB1xp67_ASAP7_75t_L g3639 ( 
.A(n_2803),
.Y(n_3639)
);

AOI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_2803),
.A2(n_2832),
.B(n_2822),
.Y(n_3640)
);

BUFx6f_ASAP7_75t_L g3641 ( 
.A(n_2822),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_2573),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3021),
.B(n_3024),
.Y(n_3643)
);

CKINVDCx20_ASAP7_75t_R g3644 ( 
.A(n_2171),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_2832),
.Y(n_3645)
);

INVx2_ASAP7_75t_L g3646 ( 
.A(n_2834),
.Y(n_3646)
);

BUFx6f_ASAP7_75t_L g3647 ( 
.A(n_2834),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_2575),
.Y(n_3648)
);

INVx2_ASAP7_75t_L g3649 ( 
.A(n_2838),
.Y(n_3649)
);

INVx2_ASAP7_75t_SL g3650 ( 
.A(n_2289),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_SL g3651 ( 
.A(n_3027),
.B(n_3032),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_L g3652 ( 
.A(n_3046),
.B(n_3052),
.Y(n_3652)
);

INVx3_ASAP7_75t_L g3653 ( 
.A(n_3186),
.Y(n_3653)
);

INVx2_ASAP7_75t_SL g3654 ( 
.A(n_2289),
.Y(n_3654)
);

CKINVDCx5p33_ASAP7_75t_R g3655 ( 
.A(n_2285),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_2576),
.Y(n_3656)
);

NAND3xp33_ASAP7_75t_L g3657 ( 
.A(n_3054),
.B(n_3066),
.C(n_3060),
.Y(n_3657)
);

AOI22xp5_ASAP7_75t_L g3658 ( 
.A1(n_3071),
.A2(n_3073),
.B1(n_3076),
.B2(n_3074),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3081),
.B(n_3082),
.Y(n_3659)
);

AOI22xp33_ASAP7_75t_L g3660 ( 
.A1(n_2838),
.A2(n_2843),
.B1(n_2846),
.B2(n_2839),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3086),
.B(n_3089),
.Y(n_3661)
);

INVx5_ASAP7_75t_L g3662 ( 
.A(n_2681),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_SL g3663 ( 
.A(n_3092),
.B(n_3104),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_2579),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3106),
.B(n_3109),
.Y(n_3665)
);

AOI22xp5_ASAP7_75t_L g3666 ( 
.A1(n_3114),
.A2(n_3116),
.B1(n_3120),
.B2(n_3117),
.Y(n_3666)
);

BUFx2_ASAP7_75t_L g3667 ( 
.A(n_2596),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3124),
.B(n_3135),
.Y(n_3668)
);

BUFx6f_ASAP7_75t_L g3669 ( 
.A(n_2839),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_2600),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_2601),
.Y(n_3671)
);

NAND2x1_ASAP7_75t_L g3672 ( 
.A(n_2221),
.B(n_2351),
.Y(n_3672)
);

BUFx3_ASAP7_75t_L g3673 ( 
.A(n_2465),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_2610),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_2613),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3137),
.B(n_3139),
.Y(n_3676)
);

AND2x6_ASAP7_75t_SL g3677 ( 
.A(n_2361),
.B(n_2079),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3140),
.B(n_3141),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_2619),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_2634),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3146),
.B(n_3157),
.Y(n_3681)
);

AOI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3161),
.A2(n_3165),
.B1(n_3175),
.B2(n_3168),
.Y(n_3682)
);

AOI22xp33_ASAP7_75t_L g3683 ( 
.A1(n_2843),
.A2(n_2848),
.B1(n_2853),
.B2(n_2846),
.Y(n_3683)
);

AND2x4_ASAP7_75t_L g3684 ( 
.A(n_2748),
.B(n_2900),
.Y(n_3684)
);

INVx3_ASAP7_75t_L g3685 ( 
.A(n_2681),
.Y(n_3685)
);

AOI22xp33_ASAP7_75t_L g3686 ( 
.A1(n_2848),
.A2(n_2875),
.B1(n_2879),
.B2(n_2853),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3177),
.B(n_3185),
.Y(n_3687)
);

INVx2_ASAP7_75t_SL g3688 ( 
.A(n_2304),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_2875),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_2879),
.Y(n_3690)
);

NAND2xp33_ASAP7_75t_L g3691 ( 
.A(n_3188),
.B(n_3204),
.Y(n_3691)
);

AND2x6_ASAP7_75t_L g3692 ( 
.A(n_2052),
.B(n_2422),
.Y(n_3692)
);

INVx2_ASAP7_75t_SL g3693 ( 
.A(n_2304),
.Y(n_3693)
);

OAI22xp33_ASAP7_75t_L g3694 ( 
.A1(n_3187),
.A2(n_3217),
.B1(n_3207),
.B2(n_2026),
.Y(n_3694)
);

OAI22xp5_ASAP7_75t_SL g3695 ( 
.A1(n_2527),
.A2(n_2118),
.B1(n_2129),
.B2(n_2128),
.Y(n_3695)
);

INVxp33_ASAP7_75t_SL g3696 ( 
.A(n_2401),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_2047),
.B(n_2012),
.Y(n_3697)
);

CKINVDCx5p33_ASAP7_75t_R g3698 ( 
.A(n_2203),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_L g3699 ( 
.A(n_2064),
.B(n_2059),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_2637),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_2639),
.Y(n_3701)
);

BUFx6f_ASAP7_75t_L g3702 ( 
.A(n_2919),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_SL g3703 ( 
.A(n_2047),
.B(n_2129),
.Y(n_3703)
);

NOR2xp67_ASAP7_75t_L g3704 ( 
.A(n_2053),
.B(n_2058),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_2919),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_SL g3706 ( 
.A(n_2060),
.B(n_2101),
.Y(n_3706)
);

BUFx8_ASAP7_75t_L g3707 ( 
.A(n_2593),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_2060),
.B(n_2063),
.Y(n_3708)
);

NOR2xp67_ASAP7_75t_L g3709 ( 
.A(n_2073),
.B(n_2070),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_2921),
.B(n_3041),
.Y(n_3710)
);

INVx3_ASAP7_75t_L g3711 ( 
.A(n_2681),
.Y(n_3711)
);

BUFx8_ASAP7_75t_SL g3712 ( 
.A(n_2149),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_2988),
.B(n_3030),
.Y(n_3713)
);

BUFx2_ASAP7_75t_L g3714 ( 
.A(n_2648),
.Y(n_3714)
);

NOR3xp33_ASAP7_75t_SL g3715 ( 
.A(n_2205),
.B(n_2087),
.C(n_2107),
.Y(n_3715)
);

NOR2xp33_ASAP7_75t_L g3716 ( 
.A(n_2425),
.B(n_2442),
.Y(n_3716)
);

OR2x2_ASAP7_75t_L g3717 ( 
.A(n_2921),
.B(n_2933),
.Y(n_3717)
);

NAND2x1p5_ASAP7_75t_L g3718 ( 
.A(n_2933),
.B(n_2939),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_L g3719 ( 
.A1(n_2939),
.A2(n_2960),
.B1(n_2988),
.B2(n_2954),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_2960),
.B(n_3197),
.Y(n_3720)
);

AND2x4_ASAP7_75t_L g3721 ( 
.A(n_2994),
.B(n_3058),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_2650),
.Y(n_3722)
);

CKINVDCx5p33_ASAP7_75t_R g3723 ( 
.A(n_2582),
.Y(n_3723)
);

O2A1O1Ixp5_ASAP7_75t_L g3724 ( 
.A1(n_2954),
.A2(n_3030),
.B(n_3034),
.C(n_3003),
.Y(n_3724)
);

INVx3_ASAP7_75t_L g3725 ( 
.A(n_2744),
.Y(n_3725)
);

NAND2xp33_ASAP7_75t_L g3726 ( 
.A(n_2104),
.B(n_2105),
.Y(n_3726)
);

CKINVDCx5p33_ASAP7_75t_R g3727 ( 
.A(n_2724),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_SL g3728 ( 
.A1(n_2652),
.A2(n_2691),
.B1(n_3085),
.B2(n_2907),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_2659),
.Y(n_3729)
);

AOI22xp5_ASAP7_75t_L g3730 ( 
.A1(n_2084),
.A2(n_2079),
.B1(n_2415),
.B2(n_2008),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_2131),
.B(n_2375),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_2462),
.A2(n_2512),
.B1(n_2627),
.B2(n_2532),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3095),
.B(n_3003),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_2662),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3178),
.B(n_3034),
.Y(n_3735)
);

AND3x2_ASAP7_75t_SL g3736 ( 
.A(n_3041),
.B(n_3084),
.C(n_3072),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_3072),
.Y(n_3737)
);

AOI22xp5_ASAP7_75t_L g3738 ( 
.A1(n_2670),
.A2(n_2680),
.B1(n_2817),
.B2(n_2791),
.Y(n_3738)
);

BUFx6f_ASAP7_75t_L g3739 ( 
.A(n_3084),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_2674),
.Y(n_3740)
);

CKINVDCx8_ASAP7_75t_R g3741 ( 
.A(n_2515),
.Y(n_3741)
);

NOR2xp33_ASAP7_75t_L g3742 ( 
.A(n_2451),
.B(n_2565),
.Y(n_3742)
);

BUFx3_ASAP7_75t_L g3743 ( 
.A(n_3055),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3087),
.B(n_3171),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_SL g3745 ( 
.A(n_2148),
.B(n_3087),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_2678),
.Y(n_3746)
);

INVx4_ASAP7_75t_L g3747 ( 
.A(n_2744),
.Y(n_3747)
);

AOI22xp33_ASAP7_75t_L g3748 ( 
.A1(n_3095),
.A2(n_3145),
.B1(n_3166),
.B2(n_3107),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3107),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_SL g3750 ( 
.A(n_3145),
.B(n_3166),
.Y(n_3750)
);

INVx5_ASAP7_75t_L g3751 ( 
.A(n_2744),
.Y(n_3751)
);

INVx3_ASAP7_75t_L g3752 ( 
.A(n_2744),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_2616),
.B(n_2640),
.Y(n_3753)
);

AND2x2_ASAP7_75t_L g3754 ( 
.A(n_3197),
.B(n_3171),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3178),
.B(n_2139),
.Y(n_3755)
);

BUFx6f_ASAP7_75t_L g3756 ( 
.A(n_2139),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_2683),
.Y(n_3757)
);

INVx1_ASAP7_75t_SL g3758 ( 
.A(n_2651),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_2076),
.B(n_2308),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_2943),
.A2(n_3125),
.B(n_3115),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_2686),
.Y(n_3761)
);

AND2x4_ASAP7_75t_L g3762 ( 
.A(n_2994),
.B(n_3058),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_2308),
.B(n_2325),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_2325),
.B(n_2326),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_2326),
.B(n_2330),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_L g3766 ( 
.A(n_2753),
.B(n_2891),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_SL g3767 ( 
.A(n_3088),
.B(n_3127),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_2693),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_2703),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_2330),
.B(n_2344),
.Y(n_3770)
);

NOR2xp33_ASAP7_75t_L g3771 ( 
.A(n_2908),
.B(n_2914),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_SL g3772 ( 
.A(n_3130),
.B(n_2112),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_2737),
.Y(n_3773)
);

AOI22xp5_ASAP7_75t_L g3774 ( 
.A1(n_2825),
.A2(n_2847),
.B1(n_2868),
.B2(n_2862),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_2740),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_2355),
.B(n_2358),
.Y(n_3776)
);

BUFx2_ASAP7_75t_L g3777 ( 
.A(n_2749),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_2344),
.B(n_2349),
.Y(n_3778)
);

INVx2_ASAP7_75t_SL g3779 ( 
.A(n_2349),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_2243),
.B(n_2246),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_2751),
.Y(n_3781)
);

AOI22xp33_ASAP7_75t_L g3782 ( 
.A1(n_2152),
.A2(n_3211),
.B1(n_3062),
.B2(n_2028),
.Y(n_3782)
);

BUFx6f_ASAP7_75t_L g3783 ( 
.A(n_2854),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_2243),
.B(n_2246),
.Y(n_3784)
);

BUFx6f_ASAP7_75t_L g3785 ( 
.A(n_2854),
.Y(n_3785)
);

NOR2xp33_ASAP7_75t_L g3786 ( 
.A(n_2108),
.B(n_2889),
.Y(n_3786)
);

INVx1_ASAP7_75t_SL g3787 ( 
.A(n_2609),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_2756),
.Y(n_3788)
);

NOR2x1_ASAP7_75t_R g3789 ( 
.A(n_2041),
.B(n_2521),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_2764),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_2152),
.A2(n_2032),
.B1(n_2458),
.B2(n_2445),
.Y(n_3791)
);

INVxp67_ASAP7_75t_L g3792 ( 
.A(n_2120),
.Y(n_3792)
);

INVx2_ASAP7_75t_SL g3793 ( 
.A(n_2056),
.Y(n_3793)
);

HB1xp67_ASAP7_75t_L g3794 ( 
.A(n_2271),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_2061),
.B(n_2082),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_2266),
.B(n_2274),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_2786),
.Y(n_3797)
);

INVxp67_ASAP7_75t_L g3798 ( 
.A(n_2123),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_2796),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_2266),
.B(n_2274),
.Y(n_3800)
);

NAND2xp5_ASAP7_75t_L g3801 ( 
.A(n_2281),
.B(n_2318),
.Y(n_3801)
);

CKINVDCx5p33_ASAP7_75t_R g3802 ( 
.A(n_2867),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_2823),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_SL g3804 ( 
.A(n_2355),
.B(n_2309),
.Y(n_3804)
);

INVx3_ASAP7_75t_L g3805 ( 
.A(n_2854),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_2281),
.B(n_2318),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_2329),
.B(n_2331),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_2828),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_2831),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_2844),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_2329),
.B(n_2331),
.Y(n_3811)
);

NOR2xp33_ASAP7_75t_L g3812 ( 
.A(n_2892),
.B(n_2942),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_2861),
.Y(n_3813)
);

OAI22xp5_ASAP7_75t_L g3814 ( 
.A1(n_2333),
.A2(n_2342),
.B1(n_2337),
.B2(n_2244),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_2333),
.B(n_2337),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_2342),
.B(n_2271),
.Y(n_3816)
);

NOR2xp67_ASAP7_75t_L g3817 ( 
.A(n_2070),
.B(n_2583),
.Y(n_3817)
);

AOI22xp5_ASAP7_75t_L g3818 ( 
.A1(n_2950),
.A2(n_2979),
.B1(n_3050),
.B2(n_2961),
.Y(n_3818)
);

NOR2xp33_ASAP7_75t_R g3819 ( 
.A(n_3055),
.B(n_2380),
.Y(n_3819)
);

INVxp67_ASAP7_75t_L g3820 ( 
.A(n_2123),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_2235),
.B(n_2270),
.Y(n_3821)
);

BUFx6f_ASAP7_75t_L g3822 ( 
.A(n_2854),
.Y(n_3822)
);

OR2x6_ASAP7_75t_L g3823 ( 
.A(n_2235),
.B(n_2270),
.Y(n_3823)
);

INVx1_ASAP7_75t_L g3824 ( 
.A(n_2882),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_SL g3825 ( 
.A(n_2350),
.B(n_3065),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_L g3826 ( 
.A(n_2902),
.B(n_2905),
.Y(n_3826)
);

INVx3_ASAP7_75t_L g3827 ( 
.A(n_2903),
.Y(n_3827)
);

AND2x4_ASAP7_75t_L g3828 ( 
.A(n_3133),
.B(n_3173),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_2080),
.A2(n_2227),
.B(n_2184),
.Y(n_3829)
);

BUFx3_ASAP7_75t_L g3830 ( 
.A(n_2903),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_2909),
.B(n_2928),
.Y(n_3831)
);

CKINVDCx20_ASAP7_75t_R g3832 ( 
.A(n_3049),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_2936),
.B(n_2953),
.Y(n_3833)
);

INVx2_ASAP7_75t_L g3834 ( 
.A(n_2955),
.Y(n_3834)
);

BUFx2_ASAP7_75t_L g3835 ( 
.A(n_2962),
.Y(n_3835)
);

OR2x2_ASAP7_75t_L g3836 ( 
.A(n_2479),
.B(n_2574),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_2992),
.Y(n_3837)
);

AOI22xp33_ASAP7_75t_L g3838 ( 
.A1(n_2810),
.A2(n_2981),
.B1(n_3093),
.B2(n_2930),
.Y(n_3838)
);

HB1xp67_ASAP7_75t_L g3839 ( 
.A(n_2993),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_2350),
.B(n_3067),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_2998),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_2999),
.Y(n_3842)
);

AND2x4_ASAP7_75t_L g3843 ( 
.A(n_3133),
.B(n_3173),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3008),
.Y(n_3844)
);

AND2x4_ASAP7_75t_L g3845 ( 
.A(n_2260),
.B(n_2296),
.Y(n_3845)
);

BUFx3_ASAP7_75t_L g3846 ( 
.A(n_3055),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3012),
.B(n_3026),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3033),
.Y(n_3848)
);

INVx2_ASAP7_75t_SL g3849 ( 
.A(n_2089),
.Y(n_3849)
);

OAI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_2176),
.A2(n_2194),
.B(n_2193),
.Y(n_3850)
);

BUFx6f_ASAP7_75t_L g3851 ( 
.A(n_2903),
.Y(n_3851)
);

OR2x2_ASAP7_75t_L g3852 ( 
.A(n_3191),
.B(n_3194),
.Y(n_3852)
);

O2A1O1Ixp5_ASAP7_75t_L g3853 ( 
.A1(n_2121),
.A2(n_2336),
.B(n_2193),
.C(n_2194),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3045),
.B(n_3047),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3048),
.B(n_3051),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_SL g3856 ( 
.A(n_3131),
.B(n_3150),
.Y(n_3856)
);

NAND3xp33_ASAP7_75t_SL g3857 ( 
.A(n_2165),
.B(n_2102),
.C(n_2378),
.Y(n_3857)
);

HB1xp67_ASAP7_75t_L g3858 ( 
.A(n_3061),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3064),
.B(n_3075),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3078),
.B(n_3079),
.Y(n_3860)
);

INVx3_ASAP7_75t_L g3861 ( 
.A(n_2903),
.Y(n_3861)
);

BUFx3_ASAP7_75t_L g3862 ( 
.A(n_2288),
.Y(n_3862)
);

AOI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3153),
.A2(n_3163),
.B1(n_2049),
.B2(n_2438),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3112),
.B(n_3119),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3142),
.Y(n_3865)
);

AND2x4_ASAP7_75t_L g3866 ( 
.A(n_2260),
.B(n_2296),
.Y(n_3866)
);

INVx2_ASAP7_75t_SL g3867 ( 
.A(n_2093),
.Y(n_3867)
);

BUFx3_ASAP7_75t_L g3868 ( 
.A(n_2288),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_SL g3869 ( 
.A(n_2039),
.B(n_2460),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3148),
.B(n_3154),
.Y(n_3870)
);

BUFx3_ASAP7_75t_L g3871 ( 
.A(n_2225),
.Y(n_3871)
);

AND2x4_ASAP7_75t_L g3872 ( 
.A(n_2583),
.B(n_2655),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3155),
.Y(n_3873)
);

NOR2xp33_ASAP7_75t_L g3874 ( 
.A(n_2066),
.B(n_2069),
.Y(n_3874)
);

BUFx3_ASAP7_75t_L g3875 ( 
.A(n_2225),
.Y(n_3875)
);

BUFx4f_ASAP7_75t_L g3876 ( 
.A(n_3103),
.Y(n_3876)
);

AND2x6_ASAP7_75t_L g3877 ( 
.A(n_3103),
.B(n_3118),
.Y(n_3877)
);

CKINVDCx5p33_ASAP7_75t_R g3878 ( 
.A(n_2382),
.Y(n_3878)
);

INVx3_ASAP7_75t_L g3879 ( 
.A(n_3103),
.Y(n_3879)
);

AND2x6_ASAP7_75t_L g3880 ( 
.A(n_3103),
.B(n_3118),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3162),
.Y(n_3881)
);

AND2x4_ASAP7_75t_L g3882 ( 
.A(n_2655),
.B(n_2656),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3167),
.Y(n_3883)
);

BUFx4f_ASAP7_75t_L g3884 ( 
.A(n_3118),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3174),
.Y(n_3885)
);

AOI21xp5_ASAP7_75t_L g3886 ( 
.A1(n_2300),
.A2(n_2345),
.B(n_2130),
.Y(n_3886)
);

INVx2_ASAP7_75t_SL g3887 ( 
.A(n_2103),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3198),
.B(n_3202),
.Y(n_3888)
);

INVx2_ASAP7_75t_SL g3889 ( 
.A(n_2110),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_2133),
.B(n_2135),
.Y(n_3890)
);

OR2x6_ASAP7_75t_L g3891 ( 
.A(n_3118),
.B(n_3123),
.Y(n_3891)
);

NAND2xp33_ASAP7_75t_SL g3892 ( 
.A(n_2940),
.B(n_3123),
.Y(n_3892)
);

AOI22xp33_ASAP7_75t_L g3893 ( 
.A1(n_2493),
.A2(n_2499),
.B1(n_2519),
.B2(n_2508),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_SL g3894 ( 
.A(n_2549),
.B(n_2550),
.Y(n_3894)
);

INVx2_ASAP7_75t_SL g3895 ( 
.A(n_2136),
.Y(n_3895)
);

OAI22xp5_ASAP7_75t_L g3896 ( 
.A1(n_2202),
.A2(n_2316),
.B1(n_2244),
.B2(n_2132),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3208),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_SL g3898 ( 
.A(n_2555),
.B(n_2580),
.Y(n_3898)
);

NOR2xp33_ASAP7_75t_L g3899 ( 
.A(n_2072),
.B(n_2015),
.Y(n_3899)
);

INVx4_ASAP7_75t_L g3900 ( 
.A(n_3123),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3216),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3218),
.B(n_2202),
.Y(n_3902)
);

AOI22xp5_ASAP7_75t_L g3903 ( 
.A1(n_2046),
.A2(n_2065),
.B1(n_2364),
.B2(n_2147),
.Y(n_3903)
);

BUFx6f_ASAP7_75t_SL g3904 ( 
.A(n_2521),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_SL g3905 ( 
.A(n_2589),
.B(n_2590),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_SL g3906 ( 
.A(n_2595),
.B(n_2604),
.Y(n_3906)
);

INVx1_ASAP7_75t_SL g3907 ( 
.A(n_3056),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_2316),
.B(n_2138),
.Y(n_3908)
);

HB1xp67_ASAP7_75t_L g3909 ( 
.A(n_2160),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_2164),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_2364),
.A2(n_2147),
.B1(n_2096),
.B2(n_2095),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_2115),
.Y(n_3912)
);

AOI22xp33_ASAP7_75t_L g3913 ( 
.A1(n_2607),
.A2(n_2628),
.B1(n_2633),
.B2(n_2608),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_SL g3914 ( 
.A(n_2643),
.B(n_2644),
.Y(n_3914)
);

INVx5_ASAP7_75t_L g3915 ( 
.A(n_3123),
.Y(n_3915)
);

OAI22xp5_ASAP7_75t_L g3916 ( 
.A1(n_2156),
.A2(n_2162),
.B1(n_2169),
.B2(n_2163),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_2654),
.B(n_2667),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_2166),
.B(n_2181),
.Y(n_3918)
);

OAI22xp5_ASAP7_75t_L g3919 ( 
.A1(n_2172),
.A2(n_2173),
.B1(n_2183),
.B2(n_2182),
.Y(n_3919)
);

BUFx6f_ASAP7_75t_SL g3920 ( 
.A(n_2547),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_2186),
.Y(n_3921)
);

NOR2xp33_ASAP7_75t_L g3922 ( 
.A(n_2252),
.B(n_2383),
.Y(n_3922)
);

NAND2x1p5_ASAP7_75t_L g3923 ( 
.A(n_2656),
.B(n_2730),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_2689),
.B(n_2711),
.Y(n_3924)
);

AND2x6_ASAP7_75t_SL g3925 ( 
.A(n_2361),
.B(n_2402),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_2189),
.Y(n_3926)
);

AND3x1_ASAP7_75t_SL g3927 ( 
.A(n_2302),
.B(n_3042),
.C(n_2524),
.Y(n_3927)
);

BUFx6f_ASAP7_75t_L g3928 ( 
.A(n_3144),
.Y(n_3928)
);

HB1xp67_ASAP7_75t_L g3929 ( 
.A(n_2187),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_2216),
.Y(n_3930)
);

BUFx3_ASAP7_75t_L g3931 ( 
.A(n_2675),
.Y(n_3931)
);

BUFx2_ASAP7_75t_L g3932 ( 
.A(n_2371),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_2220),
.B(n_2224),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_2239),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_2250),
.B(n_2273),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_SL g3936 ( 
.A(n_2712),
.B(n_2727),
.Y(n_3936)
);

NOR2xp67_ASAP7_75t_L g3937 ( 
.A(n_2730),
.B(n_2820),
.Y(n_3937)
);

BUFx6f_ASAP7_75t_L g3938 ( 
.A(n_3144),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_2190),
.Y(n_3939)
);

O2A1O1Ixp33_ASAP7_75t_L g3940 ( 
.A1(n_2176),
.A2(n_2209),
.B(n_2210),
.C(n_2201),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_2277),
.B(n_2284),
.Y(n_3941)
);

OR2x6_ASAP7_75t_L g3942 ( 
.A(n_3144),
.B(n_2820),
.Y(n_3942)
);

OAI22xp5_ASAP7_75t_L g3943 ( 
.A1(n_2191),
.A2(n_2198),
.B1(n_2211),
.B2(n_2200),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_2213),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_2312),
.Y(n_3945)
);

NOR2xp33_ASAP7_75t_L g3946 ( 
.A(n_2095),
.B(n_2096),
.Y(n_3946)
);

BUFx6f_ASAP7_75t_L g3947 ( 
.A(n_3144),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_2319),
.Y(n_3948)
);

AND2x2_ASAP7_75t_L g3949 ( 
.A(n_2322),
.B(n_2341),
.Y(n_3949)
);

AND2x4_ASAP7_75t_L g3950 ( 
.A(n_2965),
.B(n_3059),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_2343),
.B(n_2788),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_2789),
.B(n_2794),
.Y(n_3952)
);

A2O1A1Ixp33_ASAP7_75t_L g3953 ( 
.A1(n_2356),
.A2(n_2161),
.B(n_2192),
.C(n_2157),
.Y(n_3953)
);

INVx1_ASAP7_75t_L g3954 ( 
.A(n_2217),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_2233),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_2801),
.B(n_2809),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_2827),
.B(n_2837),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_2249),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_2845),
.B(n_2860),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_SL g3960 ( 
.A1(n_2380),
.A2(n_2113),
.B1(n_2630),
.B2(n_2547),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_2871),
.B(n_2872),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_2874),
.B(n_2878),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_2253),
.Y(n_3963)
);

NAND2xp5_ASAP7_75t_L g3964 ( 
.A(n_2910),
.B(n_2915),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_2927),
.B(n_2935),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_2256),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_SL g3967 ( 
.A(n_2941),
.B(n_2947),
.Y(n_3967)
);

INVx5_ASAP7_75t_L g3968 ( 
.A(n_2965),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_2957),
.B(n_2964),
.Y(n_3969)
);

AOI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_2037),
.A2(n_2155),
.B1(n_2237),
.B2(n_2109),
.Y(n_3970)
);

AOI22xp5_ASAP7_75t_L g3971 ( 
.A1(n_2109),
.A2(n_2161),
.B1(n_2192),
.B2(n_2157),
.Y(n_3971)
);

INVx4_ASAP7_75t_L g3972 ( 
.A(n_3059),
.Y(n_3972)
);

INVx2_ASAP7_75t_L g3973 ( 
.A(n_2257),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_2971),
.B(n_2972),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_2259),
.Y(n_3975)
);

AOI22xp5_ASAP7_75t_L g3976 ( 
.A1(n_2223),
.A2(n_2230),
.B1(n_2226),
.B2(n_2134),
.Y(n_3976)
);

OR2x2_ASAP7_75t_L g3977 ( 
.A(n_2263),
.B(n_2279),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_2286),
.Y(n_3978)
);

AND2x2_ASAP7_75t_SL g3979 ( 
.A(n_2378),
.B(n_3105),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_2290),
.Y(n_3980)
);

A2O1A1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_2356),
.A2(n_2223),
.B(n_2230),
.C(n_2226),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_2974),
.B(n_2977),
.Y(n_3982)
);

AND2x4_ASAP7_75t_L g3983 ( 
.A(n_3105),
.B(n_3138),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_2291),
.Y(n_3984)
);

BUFx3_ASAP7_75t_L g3985 ( 
.A(n_2370),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_2134),
.A2(n_2991),
.B1(n_2996),
.B2(n_2984),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_2293),
.Y(n_3987)
);

OAI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_2201),
.A2(n_2210),
.B(n_2209),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_2294),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3020),
.B(n_3023),
.Y(n_3990)
);

OAI22x1_ASAP7_75t_R g3991 ( 
.A1(n_2403),
.A2(n_2405),
.B1(n_2265),
.B2(n_2406),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_2295),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3028),
.B(n_3029),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3037),
.B(n_3043),
.Y(n_3994)
);

NAND2x1p5_ASAP7_75t_L g3995 ( 
.A(n_3138),
.B(n_2215),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_2301),
.Y(n_3996)
);

NOR2xp33_ASAP7_75t_L g3997 ( 
.A(n_2122),
.B(n_2098),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_2314),
.Y(n_3998)
);

NOR2x2_ASAP7_75t_L g3999 ( 
.A(n_2399),
.B(n_2264),
.Y(n_3999)
);

CKINVDCx5p33_ASAP7_75t_R g4000 ( 
.A(n_3049),
.Y(n_4000)
);

OAI21xp5_ASAP7_75t_L g4001 ( 
.A1(n_2215),
.A2(n_2229),
.B(n_2218),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3044),
.B(n_3057),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_2315),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_2317),
.Y(n_4004)
);

INVxp67_ASAP7_75t_L g4005 ( 
.A(n_2154),
.Y(n_4005)
);

AOI22xp33_ASAP7_75t_L g4006 ( 
.A1(n_3099),
.A2(n_3151),
.B1(n_3212),
.B2(n_3206),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_2320),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_2335),
.Y(n_4008)
);

BUFx2_ASAP7_75t_L g4009 ( 
.A(n_2177),
.Y(n_4009)
);

AND2x4_ASAP7_75t_L g4010 ( 
.A(n_2177),
.B(n_2180),
.Y(n_4010)
);

INVx3_ASAP7_75t_L g4011 ( 
.A(n_2180),
.Y(n_4011)
);

BUFx3_ASAP7_75t_L g4012 ( 
.A(n_2370),
.Y(n_4012)
);

BUFx3_ASAP7_75t_L g4013 ( 
.A(n_2376),
.Y(n_4013)
);

CKINVDCx5p33_ASAP7_75t_R g4014 ( 
.A(n_3160),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_2338),
.Y(n_4015)
);

INVxp67_ASAP7_75t_SL g4016 ( 
.A(n_2340),
.Y(n_4016)
);

NOR2xp33_ASAP7_75t_R g4017 ( 
.A(n_2207),
.B(n_2248),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_2346),
.Y(n_4018)
);

BUFx6f_ASAP7_75t_L g4019 ( 
.A(n_2116),
.Y(n_4019)
);

BUFx3_ASAP7_75t_L g4020 ( 
.A(n_2376),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_2218),
.A2(n_2231),
.B(n_2229),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_2352),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_2354),
.Y(n_4023)
);

CKINVDCx5p33_ASAP7_75t_R g4024 ( 
.A(n_3160),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_2367),
.Y(n_4025)
);

AND2x4_ASAP7_75t_L g4026 ( 
.A(n_2092),
.B(n_2097),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_2353),
.Y(n_4027)
);

NOR3xp33_ASAP7_75t_SL g4028 ( 
.A(n_2321),
.B(n_2391),
.C(n_2400),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3101),
.B(n_3108),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3132),
.B(n_3149),
.Y(n_4030)
);

NAND3xp33_ASAP7_75t_L g4031 ( 
.A(n_3159),
.B(n_3169),
.C(n_3164),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_2357),
.Y(n_4032)
);

BUFx3_ASAP7_75t_L g4033 ( 
.A(n_2385),
.Y(n_4033)
);

NOR2xp33_ASAP7_75t_L g4034 ( 
.A(n_2099),
.B(n_2094),
.Y(n_4034)
);

OAI22xp33_ASAP7_75t_L g4035 ( 
.A1(n_3182),
.A2(n_3214),
.B1(n_3201),
.B2(n_3192),
.Y(n_4035)
);

INVx5_ASAP7_75t_L g4036 ( 
.A(n_2815),
.Y(n_4036)
);

BUFx8_ASAP7_75t_L g4037 ( 
.A(n_2873),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_2114),
.Y(n_4038)
);

INVx3_ASAP7_75t_L g4039 ( 
.A(n_2228),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_2365),
.Y(n_4040)
);

INVx3_ASAP7_75t_L g4041 ( 
.A(n_2228),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_SL g4042 ( 
.A(n_3189),
.B(n_2455),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_2360),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_2578),
.B(n_3183),
.Y(n_4044)
);

BUFx3_ASAP7_75t_L g4045 ( 
.A(n_2116),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_2369),
.B(n_2268),
.Y(n_4046)
);

INVx5_ASAP7_75t_L g4047 ( 
.A(n_2815),
.Y(n_4047)
);

NOR2xp33_ASAP7_75t_L g4048 ( 
.A(n_2384),
.B(n_2373),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_2268),
.B(n_2303),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_2231),
.Y(n_4050)
);

BUFx6f_ASAP7_75t_L g4051 ( 
.A(n_2116),
.Y(n_4051)
);

INVx3_ASAP7_75t_L g4052 ( 
.A(n_2303),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_2347),
.B(n_2232),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_2232),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_SL g4055 ( 
.A(n_3199),
.B(n_2368),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_2347),
.B(n_2154),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_2362),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_2377),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_2372),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_2379),
.B(n_2372),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_2386),
.B(n_2391),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_SL g4062 ( 
.A(n_2167),
.B(n_2196),
.Y(n_4062)
);

NAND2xp33_ASAP7_75t_SL g4063 ( 
.A(n_2873),
.B(n_3190),
.Y(n_4063)
);

AOI21xp5_ASAP7_75t_L g4064 ( 
.A1(n_2394),
.A2(n_2264),
.B(n_3017),
.Y(n_4064)
);

BUFx4f_ASAP7_75t_L g4065 ( 
.A(n_2815),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_2208),
.B(n_2219),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_2116),
.B(n_2170),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_2170),
.B(n_2092),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_2170),
.Y(n_4069)
);

O2A1O1Ixp33_ASAP7_75t_L g4070 ( 
.A1(n_2394),
.A2(n_2334),
.B(n_2117),
.C(n_2088),
.Y(n_4070)
);

INVx3_ASAP7_75t_L g4071 ( 
.A(n_2170),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_2097),
.B(n_2206),
.Y(n_4072)
);

AOI22xp33_ASAP7_75t_L g4073 ( 
.A1(n_2269),
.A2(n_2113),
.B1(n_2178),
.B2(n_2067),
.Y(n_4073)
);

AND2x2_ASAP7_75t_L g4074 ( 
.A(n_2206),
.B(n_2212),
.Y(n_4074)
);

HB1xp67_ASAP7_75t_L g4075 ( 
.A(n_2385),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_2212),
.B(n_2071),
.Y(n_4076)
);

CKINVDCx6p67_ASAP7_75t_R g4077 ( 
.A(n_2630),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_2137),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_2071),
.B(n_2222),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_SL g4080 ( 
.A(n_2323),
.B(n_2313),
.Y(n_4080)
);

AOI21xp5_ASAP7_75t_L g4081 ( 
.A1(n_2856),
.A2(n_2880),
.B(n_3017),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_2222),
.B(n_2363),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_2374),
.Y(n_4083)
);

NOR2xp33_ASAP7_75t_L g4084 ( 
.A(n_2373),
.B(n_2241),
.Y(n_4084)
);

AOI22xp33_ASAP7_75t_L g4085 ( 
.A1(n_2178),
.A2(n_2067),
.B1(n_2267),
.B2(n_2242),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_2395),
.Y(n_4086)
);

NAND2x1p5_ASAP7_75t_L g4087 ( 
.A(n_2033),
.B(n_3190),
.Y(n_4087)
);

OAI22xp5_ASAP7_75t_L g4088 ( 
.A1(n_2366),
.A2(n_2880),
.B1(n_3017),
.B2(n_2856),
.Y(n_4088)
);

AOI22xp33_ASAP7_75t_L g4089 ( 
.A1(n_2406),
.A2(n_3036),
.B1(n_2978),
.B2(n_2963),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_2150),
.B(n_2395),
.Y(n_4090)
);

AOI22xp5_ASAP7_75t_L g4091 ( 
.A1(n_2258),
.A2(n_2332),
.B1(n_2287),
.B2(n_2238),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_SL g4092 ( 
.A(n_2044),
.B(n_2045),
.Y(n_4092)
);

AOI22xp33_ASAP7_75t_L g4093 ( 
.A1(n_2406),
.A2(n_2704),
.B1(n_3036),
.B2(n_2978),
.Y(n_4093)
);

BUFx12f_ASAP7_75t_L g4094 ( 
.A(n_2153),
.Y(n_4094)
);

AOI21xp5_ASAP7_75t_L g4095 ( 
.A1(n_2856),
.A2(n_2880),
.B(n_2869),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_2150),
.B(n_2236),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_2236),
.B(n_2245),
.Y(n_4097)
);

HB1xp67_ASAP7_75t_L g4098 ( 
.A(n_2390),
.Y(n_4098)
);

OAI22xp5_ASAP7_75t_SL g4099 ( 
.A1(n_2557),
.A2(n_3039),
.B1(n_2898),
.B2(n_2917),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_2869),
.B(n_2390),
.Y(n_4100)
);

INVx3_ASAP7_75t_L g4101 ( 
.A(n_2236),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_2392),
.Y(n_4102)
);

INVx4_ASAP7_75t_L g4103 ( 
.A(n_2245),
.Y(n_4103)
);

NOR2x2_ASAP7_75t_L g4104 ( 
.A(n_3068),
.B(n_3156),
.Y(n_4104)
);

INVx2_ASAP7_75t_SL g4105 ( 
.A(n_2245),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_2207),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_2398),
.Y(n_4107)
);

OR2x6_ASAP7_75t_L g4108 ( 
.A(n_2033),
.B(n_3090),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_SL g4109 ( 
.A(n_2396),
.B(n_2397),
.Y(n_4109)
);

INVx8_ASAP7_75t_L g4110 ( 
.A(n_2406),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_2387),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_2248),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_2396),
.Y(n_4113)
);

CKINVDCx20_ASAP7_75t_R g4114 ( 
.A(n_2153),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_2054),
.B(n_2731),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_2485),
.B(n_2731),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_2158),
.Y(n_4117)
);

INVx1_ASAP7_75t_SL g4118 ( 
.A(n_2159),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_2485),
.B(n_3090),
.Y(n_4119)
);

AND2x4_ASAP7_75t_L g4120 ( 
.A(n_2623),
.B(n_2677),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_2393),
.Y(n_4121)
);

OAI22xp5_ASAP7_75t_L g4122 ( 
.A1(n_2393),
.A2(n_2963),
.B1(n_2917),
.B2(n_2870),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_2214),
.Y(n_4123)
);

INVxp67_ASAP7_75t_L g4124 ( 
.A(n_2247),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_2297),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_2623),
.B(n_2677),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_2328),
.Y(n_4127)
);

AND2x4_ASAP7_75t_L g4128 ( 
.A(n_2661),
.B(n_2870),
.Y(n_4128)
);

INVx2_ASAP7_75t_SL g4129 ( 
.A(n_2661),
.Y(n_4129)
);

NOR2xp33_ASAP7_75t_L g4130 ( 
.A(n_2389),
.B(n_2014),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_2704),
.Y(n_4131)
);

INVx3_ASAP7_75t_L g4132 ( 
.A(n_2717),
.Y(n_4132)
);

INVx2_ASAP7_75t_SL g4133 ( 
.A(n_2717),
.Y(n_4133)
);

NAND3xp33_ASAP7_75t_SL g4134 ( 
.A(n_2404),
.B(n_2406),
.C(n_2819),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_SL g4135 ( 
.A(n_2774),
.B(n_2865),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_2774),
.Y(n_4136)
);

INVx3_ASAP7_75t_L g4137 ( 
.A(n_2819),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_2865),
.Y(n_4138)
);

INVx2_ASAP7_75t_L g4139 ( 
.A(n_2430),
.Y(n_4139)
);

BUFx8_ASAP7_75t_SL g4140 ( 
.A(n_2452),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_2471),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_2705),
.Y(n_4142)
);

INVxp67_ASAP7_75t_L g4143 ( 
.A(n_2715),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_SL g4144 ( 
.A(n_2769),
.B(n_2802),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_2812),
.Y(n_4145)
);

INVx2_ASAP7_75t_L g4146 ( 
.A(n_2821),
.Y(n_4146)
);

AND2x4_ASAP7_75t_L g4147 ( 
.A(n_2850),
.B(n_2895),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_2949),
.B(n_2985),
.Y(n_4148)
);

CKINVDCx5p33_ASAP7_75t_R g4149 ( 
.A(n_3063),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_3070),
.Y(n_4150)
);

NOR2xp33_ASAP7_75t_L g4151 ( 
.A(n_3080),
.B(n_3158),
.Y(n_4151)
);

AOI22xp5_ASAP7_75t_L g4152 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4152)
);

AOI21xp5_ASAP7_75t_L g4153 ( 
.A1(n_2081),
.A2(n_2663),
.B(n_2572),
.Y(n_4153)
);

INVx2_ASAP7_75t_L g4154 ( 
.A(n_2707),
.Y(n_4154)
);

BUFx3_ASAP7_75t_L g4155 ( 
.A(n_2175),
.Y(n_4155)
);

INVx2_ASAP7_75t_L g4156 ( 
.A(n_2707),
.Y(n_4156)
);

NOR2xp33_ASAP7_75t_L g4157 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4159)
);

HB1xp67_ASAP7_75t_L g4160 ( 
.A(n_2381),
.Y(n_4160)
);

NOR2xp33_ASAP7_75t_L g4161 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4161)
);

BUFx2_ASAP7_75t_L g4162 ( 
.A(n_2010),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4163)
);

AND2x2_ASAP7_75t_L g4164 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_2282),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_2282),
.Y(n_4167)
);

INVx5_ASAP7_75t_L g4168 ( 
.A(n_2310),
.Y(n_4168)
);

OR2x2_ASAP7_75t_L g4169 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_2707),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_2282),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_2707),
.Y(n_4172)
);

INVx2_ASAP7_75t_L g4173 ( 
.A(n_2707),
.Y(n_4173)
);

CKINVDCx20_ASAP7_75t_R g4174 ( 
.A(n_3031),
.Y(n_4174)
);

INVx1_ASAP7_75t_SL g4175 ( 
.A(n_2145),
.Y(n_4175)
);

INVx5_ASAP7_75t_L g4176 ( 
.A(n_2310),
.Y(n_4176)
);

NOR2x1p5_ASAP7_75t_L g4177 ( 
.A(n_2480),
.B(n_2653),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4179)
);

OR2x2_ASAP7_75t_L g4180 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_SL g4181 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4181)
);

INVx4_ASAP7_75t_L g4182 ( 
.A(n_2310),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_2282),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_2282),
.Y(n_4184)
);

AOI22xp33_ASAP7_75t_L g4185 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4185)
);

INVx8_ASAP7_75t_L g4186 ( 
.A(n_2310),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_SL g4187 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_2282),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_SL g4189 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_2282),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_2282),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_SL g4192 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4192)
);

INVx5_ASAP7_75t_L g4193 ( 
.A(n_2310),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_2282),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_2282),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_2707),
.Y(n_4196)
);

HB1xp67_ASAP7_75t_L g4197 ( 
.A(n_2381),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_2282),
.Y(n_4198)
);

INVx2_ASAP7_75t_SL g4199 ( 
.A(n_2381),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_2282),
.Y(n_4200)
);

AND2x6_ASAP7_75t_SL g4201 ( 
.A(n_2011),
.B(n_2408),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_SL g4202 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4202)
);

BUFx2_ASAP7_75t_L g4203 ( 
.A(n_2010),
.Y(n_4203)
);

BUFx4f_ASAP7_75t_L g4204 ( 
.A(n_2310),
.Y(n_4204)
);

INVx2_ASAP7_75t_SL g4205 ( 
.A(n_2381),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_SL g4206 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_2282),
.Y(n_4207)
);

AND2x2_ASAP7_75t_SL g4208 ( 
.A(n_2119),
.B(n_1275),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4209)
);

NOR3xp33_ASAP7_75t_SL g4210 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_L g4212 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4213)
);

AOI22xp33_ASAP7_75t_L g4214 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4214)
);

NAND2xp33_ASAP7_75t_SL g4215 ( 
.A(n_2023),
.B(n_2030),
.Y(n_4215)
);

NOR3xp33_ASAP7_75t_SL g4216 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4216)
);

INVx5_ASAP7_75t_L g4217 ( 
.A(n_2310),
.Y(n_4217)
);

BUFx3_ASAP7_75t_L g4218 ( 
.A(n_2175),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_SL g4219 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4219)
);

AOI22xp5_ASAP7_75t_L g4220 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_2707),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4222)
);

NAND3xp33_ASAP7_75t_SL g4223 ( 
.A(n_2676),
.B(n_2829),
.C(n_2728),
.Y(n_4223)
);

OAI22xp5_ASAP7_75t_L g4224 ( 
.A1(n_2009),
.A2(n_2410),
.B1(n_2411),
.B2(n_2407),
.Y(n_4224)
);

INVx2_ASAP7_75t_SL g4225 ( 
.A(n_2381),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_2707),
.Y(n_4228)
);

A2O1A1Ixp33_ASAP7_75t_L g4229 ( 
.A1(n_2958),
.A2(n_2428),
.B(n_2599),
.C(n_2566),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_2282),
.Y(n_4230)
);

INVx2_ASAP7_75t_SL g4231 ( 
.A(n_2381),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_L g4232 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4232)
);

AND2x4_ASAP7_75t_L g4233 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_2282),
.Y(n_4234)
);

NOR3xp33_ASAP7_75t_SL g4235 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_2707),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4238)
);

AOI22xp33_ASAP7_75t_L g4239 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_SL g4240 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_2282),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_2282),
.Y(n_4242)
);

NOR2xp33_ASAP7_75t_L g4243 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_2282),
.Y(n_4245)
);

INVx4_ASAP7_75t_L g4246 ( 
.A(n_2310),
.Y(n_4246)
);

AOI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_2081),
.A2(n_2663),
.B(n_2572),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4248)
);

NAND3xp33_ASAP7_75t_SL g4249 ( 
.A(n_2676),
.B(n_2829),
.C(n_2728),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4250)
);

BUFx12f_ASAP7_75t_L g4251 ( 
.A(n_3031),
.Y(n_4251)
);

CKINVDCx5p33_ASAP7_75t_R g4252 ( 
.A(n_3031),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4254)
);

AOI22xp33_ASAP7_75t_L g4255 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4255)
);

NOR2x2_ASAP7_75t_L g4256 ( 
.A(n_2199),
.B(n_2078),
.Y(n_4256)
);

CKINVDCx5p33_ASAP7_75t_R g4257 ( 
.A(n_3031),
.Y(n_4257)
);

AOI22xp5_ASAP7_75t_L g4258 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4258)
);

AOI21xp5_ASAP7_75t_L g4259 ( 
.A1(n_2081),
.A2(n_2663),
.B(n_2572),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4260)
);

INVx5_ASAP7_75t_L g4261 ( 
.A(n_2310),
.Y(n_4261)
);

HB1xp67_ASAP7_75t_L g4262 ( 
.A(n_2381),
.Y(n_4262)
);

INVx2_ASAP7_75t_L g4263 ( 
.A(n_2707),
.Y(n_4263)
);

CKINVDCx5p33_ASAP7_75t_R g4264 ( 
.A(n_3031),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_SL g4266 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_2707),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_2282),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_2282),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_2707),
.Y(n_4270)
);

OAI22xp5_ASAP7_75t_L g4271 ( 
.A1(n_2009),
.A2(n_2410),
.B1(n_2411),
.B2(n_2407),
.Y(n_4271)
);

AND2x4_ASAP7_75t_L g4272 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4272)
);

BUFx2_ASAP7_75t_L g4273 ( 
.A(n_2010),
.Y(n_4273)
);

NOR3xp33_ASAP7_75t_L g4274 ( 
.A(n_2036),
.B(n_1081),
.C(n_814),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4276)
);

INVx2_ASAP7_75t_SL g4277 ( 
.A(n_2381),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_SL g4279 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4279)
);

AND2x2_ASAP7_75t_L g4280 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4280)
);

NOR2xp33_ASAP7_75t_L g4281 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4281)
);

NOR3xp33_ASAP7_75t_SL g4282 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4282)
);

BUFx6f_ASAP7_75t_L g4283 ( 
.A(n_2707),
.Y(n_4283)
);

BUFx6f_ASAP7_75t_L g4284 ( 
.A(n_2707),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_2282),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_2707),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_2282),
.Y(n_4287)
);

AOI22xp33_ASAP7_75t_L g4288 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4288)
);

AND2x4_ASAP7_75t_L g4289 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4289)
);

AOI22xp5_ASAP7_75t_L g4290 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4290)
);

BUFx3_ASAP7_75t_L g4291 ( 
.A(n_2175),
.Y(n_4291)
);

AOI22xp33_ASAP7_75t_SL g4292 ( 
.A1(n_2017),
.A2(n_2022),
.B1(n_2027),
.B2(n_2024),
.Y(n_4292)
);

BUFx3_ASAP7_75t_L g4293 ( 
.A(n_2175),
.Y(n_4293)
);

INVx3_ASAP7_75t_L g4294 ( 
.A(n_2707),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4296)
);

INVx1_ASAP7_75t_SL g4297 ( 
.A(n_2145),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_2282),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_2282),
.Y(n_4299)
);

NAND2xp5_ASAP7_75t_L g4300 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4300)
);

NOR2x1p5_ASAP7_75t_L g4301 ( 
.A(n_2480),
.B(n_2653),
.Y(n_4301)
);

AOI22xp33_ASAP7_75t_L g4302 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4302)
);

INVx2_ASAP7_75t_SL g4303 ( 
.A(n_2381),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_SL g4304 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4304)
);

NOR2xp33_ASAP7_75t_L g4305 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4306)
);

INVx2_ASAP7_75t_SL g4307 ( 
.A(n_2381),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_2707),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4310)
);

BUFx6f_ASAP7_75t_L g4311 ( 
.A(n_2707),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_2707),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_L g4313 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4313)
);

INVx4_ASAP7_75t_L g4314 ( 
.A(n_2310),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_2282),
.Y(n_4315)
);

AND2x4_ASAP7_75t_L g4316 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_2707),
.Y(n_4318)
);

INVx4_ASAP7_75t_L g4319 ( 
.A(n_2310),
.Y(n_4319)
);

AOI22xp33_ASAP7_75t_L g4320 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4320)
);

HB1xp67_ASAP7_75t_L g4321 ( 
.A(n_2381),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_2282),
.Y(n_4322)
);

HB1xp67_ASAP7_75t_L g4323 ( 
.A(n_2381),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_2282),
.Y(n_4324)
);

AO22x1_ASAP7_75t_L g4325 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4326)
);

HB1xp67_ASAP7_75t_L g4327 ( 
.A(n_2381),
.Y(n_4327)
);

CKINVDCx5p33_ASAP7_75t_R g4328 ( 
.A(n_3031),
.Y(n_4328)
);

INVx2_ASAP7_75t_SL g4329 ( 
.A(n_2381),
.Y(n_4329)
);

O2A1O1Ixp5_ASAP7_75t_L g4330 ( 
.A1(n_2081),
.A2(n_2010),
.B(n_2958),
.C(n_2424),
.Y(n_4330)
);

OR2x6_ASAP7_75t_L g4331 ( 
.A(n_2010),
.B(n_2572),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_2707),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4333)
);

NOR2xp33_ASAP7_75t_L g4334 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_SL g4336 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4336)
);

INVx2_ASAP7_75t_SL g4337 ( 
.A(n_2381),
.Y(n_4337)
);

NOR2xp33_ASAP7_75t_L g4338 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4338)
);

NOR3xp33_ASAP7_75t_SL g4339 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4339)
);

INVx3_ASAP7_75t_L g4340 ( 
.A(n_2707),
.Y(n_4340)
);

INVx3_ASAP7_75t_L g4341 ( 
.A(n_2707),
.Y(n_4341)
);

BUFx6f_ASAP7_75t_L g4342 ( 
.A(n_2707),
.Y(n_4342)
);

OAI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_2428),
.A2(n_2599),
.B(n_2566),
.Y(n_4343)
);

INVxp67_ASAP7_75t_SL g4344 ( 
.A(n_2299),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_SL g4345 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_2282),
.Y(n_4346)
);

INVx2_ASAP7_75t_SL g4347 ( 
.A(n_2381),
.Y(n_4347)
);

AOI22xp33_ASAP7_75t_L g4348 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4349)
);

BUFx12f_ASAP7_75t_L g4350 ( 
.A(n_3031),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_2707),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_2282),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_SL g4353 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4354)
);

AND2x4_ASAP7_75t_L g4355 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4355)
);

BUFx6f_ASAP7_75t_L g4356 ( 
.A(n_2707),
.Y(n_4356)
);

CKINVDCx5p33_ASAP7_75t_R g4357 ( 
.A(n_3031),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_2282),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_SL g4360 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4360)
);

CKINVDCx20_ASAP7_75t_R g4361 ( 
.A(n_3031),
.Y(n_4361)
);

OR2x6_ASAP7_75t_L g4362 ( 
.A(n_2010),
.B(n_2572),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_2282),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_2707),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_2282),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_2707),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_2707),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_2282),
.Y(n_4368)
);

A2O1A1Ixp33_ASAP7_75t_SL g4369 ( 
.A1(n_2010),
.A2(n_2958),
.B(n_1671),
.C(n_1701),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4371)
);

NAND2xp5_ASAP7_75t_SL g4372 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4372)
);

NAND2x1p5_ASAP7_75t_L g4373 ( 
.A(n_2083),
.B(n_2081),
.Y(n_4373)
);

INVx1_ASAP7_75t_SL g4374 ( 
.A(n_2145),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_SL g4375 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4375)
);

AND2x4_ASAP7_75t_L g4376 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4376)
);

HB1xp67_ASAP7_75t_L g4377 ( 
.A(n_2381),
.Y(n_4377)
);

NAND2xp5_ASAP7_75t_L g4378 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4378)
);

AND2x2_ASAP7_75t_SL g4379 ( 
.A(n_2119),
.B(n_1275),
.Y(n_4379)
);

INVx5_ASAP7_75t_L g4380 ( 
.A(n_2310),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_2707),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4382)
);

NOR2xp33_ASAP7_75t_L g4383 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4383)
);

OAI22xp5_ASAP7_75t_SL g4384 ( 
.A1(n_2743),
.A2(n_2624),
.B1(n_2528),
.B2(n_2472),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4385)
);

OR2x2_ASAP7_75t_SL g4386 ( 
.A(n_2698),
.B(n_814),
.Y(n_4386)
);

HB1xp67_ASAP7_75t_L g4387 ( 
.A(n_2381),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_2707),
.Y(n_4388)
);

BUFx6f_ASAP7_75t_L g4389 ( 
.A(n_2707),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_2282),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_2282),
.Y(n_4391)
);

INVx2_ASAP7_75t_SL g4392 ( 
.A(n_2381),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_2707),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4394)
);

NOR2x1p5_ASAP7_75t_L g4395 ( 
.A(n_2480),
.B(n_2653),
.Y(n_4395)
);

INVx2_ASAP7_75t_SL g4396 ( 
.A(n_2381),
.Y(n_4396)
);

NOR3xp33_ASAP7_75t_L g4397 ( 
.A(n_2036),
.B(n_1081),
.C(n_814),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_2282),
.Y(n_4398)
);

AND2x2_ASAP7_75t_SL g4399 ( 
.A(n_2119),
.B(n_1275),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4400)
);

NOR2xp33_ASAP7_75t_L g4401 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_L g4402 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_2282),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_2282),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_SL g4405 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4405)
);

INVx3_ASAP7_75t_L g4406 ( 
.A(n_2707),
.Y(n_4406)
);

OAI22xp5_ASAP7_75t_L g4407 ( 
.A1(n_2009),
.A2(n_2410),
.B1(n_2411),
.B2(n_2407),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_2707),
.Y(n_4408)
);

AND2x2_ASAP7_75t_L g4409 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4409)
);

INVx2_ASAP7_75t_L g4410 ( 
.A(n_2707),
.Y(n_4410)
);

NOR2xp33_ASAP7_75t_L g4411 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4411)
);

BUFx2_ASAP7_75t_L g4412 ( 
.A(n_2010),
.Y(n_4412)
);

BUFx6f_ASAP7_75t_L g4413 ( 
.A(n_2707),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_2282),
.Y(n_4414)
);

CKINVDCx5p33_ASAP7_75t_R g4415 ( 
.A(n_3031),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_2282),
.Y(n_4416)
);

A2O1A1Ixp33_ASAP7_75t_L g4417 ( 
.A1(n_2958),
.A2(n_2428),
.B(n_2599),
.C(n_2566),
.Y(n_4417)
);

NOR2xp33_ASAP7_75t_L g4418 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4418)
);

NAND2x1p5_ASAP7_75t_L g4419 ( 
.A(n_2083),
.B(n_2081),
.Y(n_4419)
);

INVx1_ASAP7_75t_SL g4420 ( 
.A(n_2145),
.Y(n_4420)
);

INVx2_ASAP7_75t_SL g4421 ( 
.A(n_2381),
.Y(n_4421)
);

NAND2x1p5_ASAP7_75t_L g4422 ( 
.A(n_2083),
.B(n_2081),
.Y(n_4422)
);

AOI22xp5_ASAP7_75t_L g4423 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4423)
);

CKINVDCx5p33_ASAP7_75t_R g4424 ( 
.A(n_3031),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_2282),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_2282),
.Y(n_4427)
);

OR2x2_ASAP7_75t_L g4428 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4428)
);

NOR2x1p5_ASAP7_75t_L g4429 ( 
.A(n_2480),
.B(n_2653),
.Y(n_4429)
);

INVx3_ASAP7_75t_L g4430 ( 
.A(n_2707),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4431)
);

AND3x1_ASAP7_75t_L g4432 ( 
.A(n_2676),
.B(n_924),
.C(n_2728),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_SL g4433 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_2707),
.Y(n_4434)
);

INVx3_ASAP7_75t_L g4435 ( 
.A(n_2707),
.Y(n_4435)
);

OR2x2_ASAP7_75t_L g4436 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_2707),
.Y(n_4437)
);

AOI22xp5_ASAP7_75t_L g4438 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_SL g4439 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_2707),
.Y(n_4440)
);

NOR2x1_ASAP7_75t_L g4441 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4442)
);

CKINVDCx5p33_ASAP7_75t_R g4443 ( 
.A(n_3031),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_SL g4444 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4444)
);

INVxp33_ASAP7_75t_L g4445 ( 
.A(n_2079),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_SL g4446 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4446)
);

INVxp67_ASAP7_75t_SL g4447 ( 
.A(n_2299),
.Y(n_4447)
);

AND2x4_ASAP7_75t_L g4448 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_SL g4450 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4450)
);

OAI21xp5_ASAP7_75t_L g4451 ( 
.A1(n_2428),
.A2(n_2599),
.B(n_2566),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4452)
);

AND2x4_ASAP7_75t_L g4453 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4453)
);

AND2x4_ASAP7_75t_L g4454 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4454)
);

CKINVDCx5p33_ASAP7_75t_R g4455 ( 
.A(n_3031),
.Y(n_4455)
);

NOR3xp33_ASAP7_75t_SL g4456 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4456)
);

INVx3_ASAP7_75t_L g4457 ( 
.A(n_2707),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_2282),
.Y(n_4458)
);

AND2x4_ASAP7_75t_L g4459 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4459)
);

AND2x4_ASAP7_75t_L g4460 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4460)
);

INVx4_ASAP7_75t_L g4461 ( 
.A(n_2310),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_2282),
.Y(n_4462)
);

CKINVDCx8_ASAP7_75t_R g4463 ( 
.A(n_2151),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_SL g4464 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_SL g4465 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4465)
);

NOR2x1p5_ASAP7_75t_L g4466 ( 
.A(n_2480),
.B(n_2653),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_2282),
.Y(n_4468)
);

CKINVDCx5p33_ASAP7_75t_R g4469 ( 
.A(n_3031),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4470)
);

BUFx2_ASAP7_75t_L g4471 ( 
.A(n_2010),
.Y(n_4471)
);

NAND2x1p5_ASAP7_75t_L g4472 ( 
.A(n_2083),
.B(n_2081),
.Y(n_4472)
);

BUFx6f_ASAP7_75t_L g4473 ( 
.A(n_2707),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4475)
);

BUFx3_ASAP7_75t_L g4476 ( 
.A(n_2560),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_2282),
.Y(n_4477)
);

AND2x2_ASAP7_75t_L g4478 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_2282),
.Y(n_4479)
);

BUFx6f_ASAP7_75t_L g4480 ( 
.A(n_2707),
.Y(n_4480)
);

NOR2x2_ASAP7_75t_L g4481 ( 
.A(n_2199),
.B(n_2078),
.Y(n_4481)
);

AOI22xp5_ASAP7_75t_L g4482 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4483)
);

INVx2_ASAP7_75t_L g4484 ( 
.A(n_2707),
.Y(n_4484)
);

AOI22xp33_ASAP7_75t_L g4485 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_2707),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_2282),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4488)
);

NOR2xp33_ASAP7_75t_L g4489 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4491)
);

INVx2_ASAP7_75t_L g4492 ( 
.A(n_2707),
.Y(n_4492)
);

BUFx6f_ASAP7_75t_L g4493 ( 
.A(n_2707),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_SL g4494 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4494)
);

OR2x2_ASAP7_75t_L g4495 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_2282),
.Y(n_4496)
);

NAND3xp33_ASAP7_75t_L g4497 ( 
.A(n_3209),
.B(n_1081),
.C(n_814),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4498)
);

INVx2_ASAP7_75t_L g4499 ( 
.A(n_2707),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_2282),
.Y(n_4500)
);

OR2x6_ASAP7_75t_L g4501 ( 
.A(n_2010),
.B(n_2572),
.Y(n_4501)
);

AND2x6_ASAP7_75t_SL g4502 ( 
.A(n_2011),
.B(n_2408),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_2707),
.Y(n_4503)
);

BUFx6f_ASAP7_75t_L g4504 ( 
.A(n_2707),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_2707),
.Y(n_4505)
);

OR2x6_ASAP7_75t_L g4506 ( 
.A(n_2010),
.B(n_2572),
.Y(n_4506)
);

AND2x6_ASAP7_75t_L g4507 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4507)
);

NOR2xp33_ASAP7_75t_L g4508 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_2282),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_2707),
.Y(n_4510)
);

NOR2xp33_ASAP7_75t_L g4511 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4511)
);

BUFx4f_ASAP7_75t_L g4512 ( 
.A(n_2310),
.Y(n_4512)
);

INVx2_ASAP7_75t_L g4513 ( 
.A(n_2707),
.Y(n_4513)
);

AND2x4_ASAP7_75t_L g4514 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4514)
);

NOR2xp33_ASAP7_75t_R g4515 ( 
.A(n_3122),
.B(n_716),
.Y(n_4515)
);

INVx2_ASAP7_75t_SL g4516 ( 
.A(n_2381),
.Y(n_4516)
);

INVx4_ASAP7_75t_L g4517 ( 
.A(n_2310),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_2707),
.Y(n_4519)
);

BUFx6f_ASAP7_75t_L g4520 ( 
.A(n_2707),
.Y(n_4520)
);

AOI22xp5_ASAP7_75t_L g4521 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_2707),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_2707),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_2282),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_2707),
.Y(n_4525)
);

BUFx6f_ASAP7_75t_SL g4526 ( 
.A(n_2310),
.Y(n_4526)
);

INVx5_ASAP7_75t_L g4527 ( 
.A(n_2310),
.Y(n_4527)
);

AOI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_2282),
.Y(n_4530)
);

AOI22xp5_ASAP7_75t_L g4531 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4531)
);

AOI22xp5_ASAP7_75t_L g4532 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_SL g4534 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4534)
);

OAI22xp5_ASAP7_75t_L g4535 ( 
.A1(n_2009),
.A2(n_2410),
.B1(n_2411),
.B2(n_2407),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_2282),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_SL g4537 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_2282),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_2707),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_2282),
.Y(n_4540)
);

AOI22xp5_ASAP7_75t_L g4541 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_SL g4542 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4542)
);

BUFx6f_ASAP7_75t_L g4543 ( 
.A(n_2707),
.Y(n_4543)
);

INVx3_ASAP7_75t_L g4544 ( 
.A(n_2707),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_2282),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_2282),
.Y(n_4547)
);

INVx3_ASAP7_75t_L g4548 ( 
.A(n_2707),
.Y(n_4548)
);

OAI221xp5_ASAP7_75t_L g4549 ( 
.A1(n_2036),
.A2(n_2035),
.B1(n_2018),
.B2(n_2728),
.C(n_2676),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_2707),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_2282),
.Y(n_4552)
);

NOR2xp33_ASAP7_75t_L g4553 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4554)
);

INVx3_ASAP7_75t_L g4555 ( 
.A(n_2707),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4556)
);

INVx3_ASAP7_75t_L g4557 ( 
.A(n_2707),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4558)
);

INVx1_ASAP7_75t_L g4559 ( 
.A(n_2282),
.Y(n_4559)
);

AOI22xp33_ASAP7_75t_L g4560 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4560)
);

INVx1_ASAP7_75t_SL g4561 ( 
.A(n_2145),
.Y(n_4561)
);

AOI21xp5_ASAP7_75t_L g4562 ( 
.A1(n_2081),
.A2(n_2663),
.B(n_2572),
.Y(n_4562)
);

AND2x2_ASAP7_75t_SL g4563 ( 
.A(n_2119),
.B(n_1275),
.Y(n_4563)
);

NOR2xp33_ASAP7_75t_L g4564 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4564)
);

AND2x2_ASAP7_75t_L g4565 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4565)
);

NAND2xp33_ASAP7_75t_L g4566 ( 
.A(n_2428),
.B(n_2566),
.Y(n_4566)
);

OR2x6_ASAP7_75t_L g4567 ( 
.A(n_2010),
.B(n_2572),
.Y(n_4567)
);

INVx4_ASAP7_75t_L g4568 ( 
.A(n_2310),
.Y(n_4568)
);

OR2x2_ASAP7_75t_L g4569 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4569)
);

NAND2x1p5_ASAP7_75t_L g4570 ( 
.A(n_2083),
.B(n_2081),
.Y(n_4570)
);

AND2x4_ASAP7_75t_L g4571 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_L g4572 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4572)
);

OAI22xp5_ASAP7_75t_L g4573 ( 
.A1(n_2009),
.A2(n_2410),
.B1(n_2411),
.B2(n_2407),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_2707),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_2282),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_2282),
.Y(n_4576)
);

INVx3_ASAP7_75t_L g4577 ( 
.A(n_2707),
.Y(n_4577)
);

A2O1A1Ixp33_ASAP7_75t_L g4578 ( 
.A1(n_2958),
.A2(n_2428),
.B(n_2599),
.C(n_2566),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_2282),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4580)
);

NOR2xp33_ASAP7_75t_L g4581 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4581)
);

AND2x6_ASAP7_75t_SL g4582 ( 
.A(n_2011),
.B(n_2408),
.Y(n_4582)
);

NOR2xp33_ASAP7_75t_R g4583 ( 
.A(n_3122),
.B(n_716),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4584)
);

BUFx2_ASAP7_75t_L g4585 ( 
.A(n_2010),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_SL g4586 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4586)
);

OAI22xp33_ASAP7_75t_L g4587 ( 
.A1(n_2035),
.A2(n_2036),
.B1(n_2622),
.B2(n_2586),
.Y(n_4587)
);

HB1xp67_ASAP7_75t_L g4588 ( 
.A(n_2381),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4589)
);

INVx2_ASAP7_75t_L g4590 ( 
.A(n_2707),
.Y(n_4590)
);

NAND2x1p5_ASAP7_75t_L g4591 ( 
.A(n_2083),
.B(n_2081),
.Y(n_4591)
);

AND2x6_ASAP7_75t_SL g4592 ( 
.A(n_2011),
.B(n_2408),
.Y(n_4592)
);

AOI22xp33_ASAP7_75t_L g4593 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_2282),
.Y(n_4594)
);

BUFx3_ASAP7_75t_L g4595 ( 
.A(n_2175),
.Y(n_4595)
);

OAI21xp33_ASAP7_75t_L g4596 ( 
.A1(n_3209),
.A2(n_2408),
.B(n_2011),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_2282),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4598)
);

OR2x2_ASAP7_75t_L g4599 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4600)
);

INVx2_ASAP7_75t_SL g4601 ( 
.A(n_2381),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4603)
);

A2O1A1Ixp33_ASAP7_75t_L g4604 ( 
.A1(n_2958),
.A2(n_2428),
.B(n_2599),
.C(n_2566),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_2707),
.Y(n_4606)
);

BUFx3_ASAP7_75t_L g4607 ( 
.A(n_2560),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_2282),
.Y(n_4609)
);

INVx3_ASAP7_75t_L g4610 ( 
.A(n_2707),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4611)
);

BUFx6f_ASAP7_75t_L g4612 ( 
.A(n_2707),
.Y(n_4612)
);

INVx1_ASAP7_75t_SL g4613 ( 
.A(n_2145),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_2707),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_2282),
.Y(n_4615)
);

AOI22xp5_ASAP7_75t_L g4616 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4617)
);

AOI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4618)
);

HB1xp67_ASAP7_75t_L g4619 ( 
.A(n_2381),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4620)
);

BUFx3_ASAP7_75t_L g4621 ( 
.A(n_2560),
.Y(n_4621)
);

AOI22xp5_ASAP7_75t_L g4622 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_2282),
.Y(n_4623)
);

AOI22xp33_ASAP7_75t_L g4624 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_SL g4626 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_SL g4628 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_2282),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_2282),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_SL g4631 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_2282),
.Y(n_4633)
);

BUFx3_ASAP7_75t_L g4634 ( 
.A(n_2560),
.Y(n_4634)
);

INVx2_ASAP7_75t_SL g4635 ( 
.A(n_2381),
.Y(n_4635)
);

NAND3xp33_ASAP7_75t_SL g4636 ( 
.A(n_2676),
.B(n_2829),
.C(n_2728),
.Y(n_4636)
);

INVx2_ASAP7_75t_SL g4637 ( 
.A(n_2381),
.Y(n_4637)
);

INVx1_ASAP7_75t_SL g4638 ( 
.A(n_2145),
.Y(n_4638)
);

AND2x4_ASAP7_75t_L g4639 ( 
.A(n_2381),
.B(n_2388),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_2282),
.Y(n_4640)
);

AOI22xp5_ASAP7_75t_L g4641 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_2707),
.Y(n_4642)
);

BUFx5_ASAP7_75t_L g4643 ( 
.A(n_2560),
.Y(n_4643)
);

CKINVDCx20_ASAP7_75t_R g4644 ( 
.A(n_3031),
.Y(n_4644)
);

NOR3xp33_ASAP7_75t_SL g4645 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4645)
);

INVxp67_ASAP7_75t_L g4646 ( 
.A(n_2120),
.Y(n_4646)
);

OAI22xp5_ASAP7_75t_L g4647 ( 
.A1(n_2009),
.A2(n_2410),
.B1(n_2411),
.B2(n_2407),
.Y(n_4647)
);

NAND2xp33_ASAP7_75t_R g4648 ( 
.A(n_2017),
.B(n_2022),
.Y(n_4648)
);

NOR3xp33_ASAP7_75t_SL g4649 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_2282),
.Y(n_4651)
);

INVx5_ASAP7_75t_L g4652 ( 
.A(n_2310),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_2282),
.Y(n_4653)
);

AOI22xp33_ASAP7_75t_L g4654 ( 
.A1(n_2017),
.A2(n_2024),
.B1(n_2027),
.B2(n_2022),
.Y(n_4654)
);

CKINVDCx5p33_ASAP7_75t_R g4655 ( 
.A(n_3031),
.Y(n_4655)
);

NOR2xp33_ASAP7_75t_L g4656 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_2707),
.Y(n_4657)
);

INVx5_ASAP7_75t_L g4658 ( 
.A(n_2310),
.Y(n_4658)
);

BUFx6f_ASAP7_75t_L g4659 ( 
.A(n_2707),
.Y(n_4659)
);

BUFx2_ASAP7_75t_L g4660 ( 
.A(n_2010),
.Y(n_4660)
);

NOR3xp33_ASAP7_75t_SL g4661 ( 
.A(n_2472),
.B(n_1744),
.C(n_1644),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_2707),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_2707),
.Y(n_4663)
);

CKINVDCx5p33_ASAP7_75t_R g4664 ( 
.A(n_3031),
.Y(n_4664)
);

BUFx6f_ASAP7_75t_L g4665 ( 
.A(n_2707),
.Y(n_4665)
);

INVx3_ASAP7_75t_L g4666 ( 
.A(n_2707),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_2707),
.Y(n_4667)
);

BUFx2_ASAP7_75t_R g4668 ( 
.A(n_2041),
.Y(n_4668)
);

NOR2xp33_ASAP7_75t_L g4669 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4669)
);

NOR2xp67_ASAP7_75t_L g4670 ( 
.A(n_2632),
.B(n_3113),
.Y(n_4670)
);

OR2x2_ASAP7_75t_SL g4671 ( 
.A(n_2698),
.B(n_814),
.Y(n_4671)
);

BUFx4f_ASAP7_75t_SL g4672 ( 
.A(n_2149),
.Y(n_4672)
);

NAND3xp33_ASAP7_75t_SL g4673 ( 
.A(n_2676),
.B(n_2829),
.C(n_2728),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4674)
);

AOI22xp5_ASAP7_75t_L g4675 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_2282),
.Y(n_4676)
);

OAI22xp33_ASAP7_75t_L g4677 ( 
.A1(n_2035),
.A2(n_2036),
.B1(n_2622),
.B2(n_2586),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_2282),
.Y(n_4678)
);

NAND3xp33_ASAP7_75t_SL g4679 ( 
.A(n_2676),
.B(n_2829),
.C(n_2728),
.Y(n_4679)
);

OR2x2_ASAP7_75t_L g4680 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_2707),
.Y(n_4681)
);

HB1xp67_ASAP7_75t_L g4682 ( 
.A(n_2381),
.Y(n_4682)
);

BUFx3_ASAP7_75t_L g4683 ( 
.A(n_2560),
.Y(n_4683)
);

HB1xp67_ASAP7_75t_L g4684 ( 
.A(n_2381),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_2282),
.Y(n_4685)
);

INVx3_ASAP7_75t_L g4686 ( 
.A(n_2707),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_2282),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_2282),
.Y(n_4688)
);

INVx3_ASAP7_75t_L g4689 ( 
.A(n_2707),
.Y(n_4689)
);

INVxp67_ASAP7_75t_SL g4690 ( 
.A(n_2299),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_2282),
.Y(n_4691)
);

INVx3_ASAP7_75t_L g4692 ( 
.A(n_2707),
.Y(n_4692)
);

INVx3_ASAP7_75t_L g4693 ( 
.A(n_2707),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_L g4694 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_2282),
.Y(n_4695)
);

AOI21xp33_ASAP7_75t_L g4696 ( 
.A1(n_2958),
.A2(n_2566),
.B(n_2428),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_L g4697 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4697)
);

NAND2xp5_ASAP7_75t_L g4698 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4700)
);

OAI22xp5_ASAP7_75t_L g4701 ( 
.A1(n_2009),
.A2(n_2410),
.B1(n_2411),
.B2(n_2407),
.Y(n_4701)
);

OR2x2_ASAP7_75t_L g4702 ( 
.A(n_2013),
.B(n_2424),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_2707),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_2010),
.B(n_2428),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_2707),
.Y(n_4705)
);

OAI22xp33_ASAP7_75t_L g4706 ( 
.A1(n_2035),
.A2(n_2036),
.B1(n_2622),
.B2(n_2586),
.Y(n_4706)
);

NOR2x2_ASAP7_75t_L g4707 ( 
.A(n_2199),
.B(n_2078),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_2707),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_SL g4709 ( 
.A(n_2543),
.B(n_2581),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_2707),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_2282),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_2282),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_2282),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_2282),
.Y(n_4715)
);

NOR2x2_ASAP7_75t_L g4716 ( 
.A(n_2199),
.B(n_2078),
.Y(n_4716)
);

AOI22xp5_ASAP7_75t_L g4717 ( 
.A1(n_2011),
.A2(n_2416),
.B1(n_2454),
.B2(n_2408),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_2414),
.B(n_2433),
.Y(n_4719)
);

O2A1O1Ixp33_ASAP7_75t_L g4720 ( 
.A1(n_2018),
.A2(n_2566),
.B(n_2599),
.C(n_2428),
.Y(n_4720)
);

NOR2xp33_ASAP7_75t_L g4721 ( 
.A(n_2036),
.B(n_2011),
.Y(n_4721)
);

NOR2xp33_ASAP7_75t_L g4722 ( 
.A(n_3275),
.B(n_4596),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_3266),
.B(n_3220),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_3575),
.B(n_3585),
.Y(n_4724)
);

INVx1_ASAP7_75t_SL g4725 ( 
.A(n_3758),
.Y(n_4725)
);

OAI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_3257),
.A2(n_4157),
.B(n_3221),
.Y(n_4726)
);

AOI21xp5_ASAP7_75t_L g4727 ( 
.A1(n_3310),
.A2(n_4247),
.B(n_4153),
.Y(n_4727)
);

NOR2xp67_ASAP7_75t_SL g4728 ( 
.A(n_3741),
.B(n_4549),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_3575),
.B(n_3585),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_3228),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_L g4731 ( 
.A1(n_3310),
.A2(n_4247),
.B(n_4153),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_3228),
.Y(n_4732)
);

INVx4_ASAP7_75t_L g4733 ( 
.A(n_4036),
.Y(n_4733)
);

INVx3_ASAP7_75t_L g4734 ( 
.A(n_3295),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_3575),
.B(n_3585),
.Y(n_4735)
);

AOI22xp5_ASAP7_75t_L g4736 ( 
.A1(n_4384),
.A2(n_4223),
.B1(n_4249),
.B2(n_3265),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_3228),
.Y(n_4737)
);

A2O1A1Ixp33_ASAP7_75t_L g4738 ( 
.A1(n_3496),
.A2(n_3221),
.B(n_4161),
.C(n_4157),
.Y(n_4738)
);

BUFx12f_ASAP7_75t_L g4739 ( 
.A(n_4251),
.Y(n_4739)
);

O2A1O1Ixp33_ASAP7_75t_L g4740 ( 
.A1(n_3257),
.A2(n_3410),
.B(n_3436),
.C(n_3265),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_3266),
.B(n_3220),
.Y(n_4741)
);

O2A1O1Ixp33_ASAP7_75t_L g4742 ( 
.A1(n_3410),
.A2(n_3436),
.B(n_4249),
.C(n_4223),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_L g4743 ( 
.A(n_3233),
.B(n_3234),
.Y(n_4743)
);

INVx2_ASAP7_75t_L g4744 ( 
.A(n_3405),
.Y(n_4744)
);

AOI22xp5_ASAP7_75t_L g4745 ( 
.A1(n_4384),
.A2(n_4673),
.B1(n_4679),
.B2(n_4636),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_3233),
.B(n_3234),
.Y(n_4746)
);

NOR2xp33_ASAP7_75t_L g4747 ( 
.A(n_3275),
.B(n_4596),
.Y(n_4747)
);

AOI21xp5_ASAP7_75t_L g4748 ( 
.A1(n_4259),
.A2(n_4562),
.B(n_4566),
.Y(n_4748)
);

OR2x6_ASAP7_75t_L g4749 ( 
.A(n_4186),
.B(n_4331),
.Y(n_4749)
);

AOI21xp5_ASAP7_75t_L g4750 ( 
.A1(n_4259),
.A2(n_4562),
.B(n_4566),
.Y(n_4750)
);

AOI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_3224),
.A2(n_4417),
.B(n_4229),
.Y(n_4751)
);

INVx2_ASAP7_75t_L g4752 ( 
.A(n_3405),
.Y(n_4752)
);

NAND2xp5_ASAP7_75t_SL g4753 ( 
.A(n_4292),
.B(n_3360),
.Y(n_4753)
);

O2A1O1Ixp33_ASAP7_75t_L g4754 ( 
.A1(n_4636),
.A2(n_4679),
.B(n_4673),
.C(n_3423),
.Y(n_4754)
);

OAI22xp5_ASAP7_75t_L g4755 ( 
.A1(n_3496),
.A2(n_3493),
.B1(n_4185),
.B2(n_3225),
.Y(n_4755)
);

INVx2_ASAP7_75t_L g4756 ( 
.A(n_3405),
.Y(n_4756)
);

AOI21xp5_ASAP7_75t_L g4757 ( 
.A1(n_3224),
.A2(n_4417),
.B(n_4229),
.Y(n_4757)
);

BUFx6f_ASAP7_75t_L g4758 ( 
.A(n_3284),
.Y(n_4758)
);

AOI21xp5_ASAP7_75t_L g4759 ( 
.A1(n_4578),
.A2(n_4604),
.B(n_3467),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4158),
.B(n_4159),
.Y(n_4760)
);

CKINVDCx8_ASAP7_75t_R g4761 ( 
.A(n_3284),
.Y(n_4761)
);

BUFx2_ASAP7_75t_L g4762 ( 
.A(n_3823),
.Y(n_4762)
);

INVx4_ASAP7_75t_L g4763 ( 
.A(n_4036),
.Y(n_4763)
);

INVxp67_ASAP7_75t_L g4764 ( 
.A(n_3909),
.Y(n_4764)
);

BUFx6f_ASAP7_75t_L g4765 ( 
.A(n_3284),
.Y(n_4765)
);

O2A1O1Ixp33_ASAP7_75t_L g4766 ( 
.A1(n_3423),
.A2(n_3438),
.B(n_3444),
.C(n_3440),
.Y(n_4766)
);

BUFx2_ASAP7_75t_L g4767 ( 
.A(n_3823),
.Y(n_4767)
);

O2A1O1Ixp33_ASAP7_75t_SL g4768 ( 
.A1(n_4369),
.A2(n_3322),
.B(n_3238),
.C(n_4587),
.Y(n_4768)
);

A2O1A1Ixp33_ASAP7_75t_L g4769 ( 
.A1(n_4161),
.A2(n_4212),
.B(n_4243),
.C(n_4232),
.Y(n_4769)
);

NOR2xp33_ASAP7_75t_L g4770 ( 
.A(n_3226),
.B(n_3236),
.Y(n_4770)
);

AND2x4_ASAP7_75t_L g4771 ( 
.A(n_3301),
.B(n_3381),
.Y(n_4771)
);

AOI21xp5_ASAP7_75t_L g4772 ( 
.A1(n_4578),
.A2(n_4604),
.B(n_3467),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4158),
.B(n_4159),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_SL g4774 ( 
.A(n_4292),
.B(n_3360),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4163),
.B(n_4166),
.Y(n_4775)
);

AOI21xp5_ASAP7_75t_L g4776 ( 
.A1(n_3278),
.A2(n_4447),
.B(n_4344),
.Y(n_4776)
);

AOI21xp5_ASAP7_75t_L g4777 ( 
.A1(n_3278),
.A2(n_4447),
.B(n_4344),
.Y(n_4777)
);

AOI21xp5_ASAP7_75t_L g4778 ( 
.A1(n_4690),
.A2(n_4451),
.B(n_4343),
.Y(n_4778)
);

NAND2xp5_ASAP7_75t_SL g4779 ( 
.A(n_3376),
.B(n_3243),
.Y(n_4779)
);

NOR2xp33_ASAP7_75t_L g4780 ( 
.A(n_3226),
.B(n_3236),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_SL g4781 ( 
.A(n_3376),
.B(n_3243),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_3405),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_3405),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4178),
.B(n_4179),
.Y(n_4784)
);

O2A1O1Ixp33_ASAP7_75t_L g4785 ( 
.A1(n_3438),
.A2(n_3440),
.B(n_3444),
.C(n_4549),
.Y(n_4785)
);

NOR3xp33_ASAP7_75t_L g4786 ( 
.A(n_3401),
.B(n_4677),
.C(n_4587),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4178),
.B(n_4179),
.Y(n_4787)
);

NOR2xp33_ASAP7_75t_L g4788 ( 
.A(n_3251),
.B(n_3252),
.Y(n_4788)
);

AOI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4690),
.A2(n_4451),
.B(n_4343),
.Y(n_4789)
);

CKINVDCx5p33_ASAP7_75t_R g4790 ( 
.A(n_3698),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_3481),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_3405),
.Y(n_4792)
);

O2A1O1Ixp33_ASAP7_75t_L g4793 ( 
.A1(n_4677),
.A2(n_4706),
.B(n_3238),
.C(n_3322),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4209),
.B(n_4211),
.Y(n_4794)
);

NOR2xp33_ASAP7_75t_L g4795 ( 
.A(n_3251),
.B(n_3252),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4209),
.B(n_4211),
.Y(n_4796)
);

OR2x6_ASAP7_75t_L g4797 ( 
.A(n_4186),
.B(n_4331),
.Y(n_4797)
);

AOI21xp5_ASAP7_75t_L g4798 ( 
.A1(n_4331),
.A2(n_4501),
.B(n_4362),
.Y(n_4798)
);

OAI21xp33_ASAP7_75t_L g4799 ( 
.A1(n_4212),
.A2(n_4243),
.B(n_4232),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_3405),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_3589),
.B(n_3634),
.Y(n_4801)
);

AOI21xp5_ASAP7_75t_L g4802 ( 
.A1(n_4331),
.A2(n_4501),
.B(n_4362),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4222),
.B(n_4226),
.Y(n_4803)
);

BUFx2_ASAP7_75t_L g4804 ( 
.A(n_3823),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4222),
.B(n_4226),
.Y(n_4805)
);

AOI221xp5_ASAP7_75t_L g4806 ( 
.A1(n_4281),
.A2(n_4334),
.B1(n_4383),
.B2(n_4338),
.C(n_4305),
.Y(n_4806)
);

O2A1O1Ixp33_ASAP7_75t_L g4807 ( 
.A1(n_4706),
.A2(n_3401),
.B(n_4369),
.C(n_3459),
.Y(n_4807)
);

INVx3_ASAP7_75t_L g4808 ( 
.A(n_3295),
.Y(n_4808)
);

OAI22xp5_ASAP7_75t_L g4809 ( 
.A1(n_3493),
.A2(n_4185),
.B1(n_4214),
.B2(n_3225),
.Y(n_4809)
);

AOI33xp33_ASAP7_75t_L g4810 ( 
.A1(n_4214),
.A2(n_4288),
.A3(n_4239),
.B1(n_4320),
.B2(n_4302),
.B3(n_4255),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_3520),
.Y(n_4811)
);

NOR2xp67_ASAP7_75t_L g4812 ( 
.A(n_3657),
.B(n_3516),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_L g4813 ( 
.A(n_4227),
.B(n_4236),
.Y(n_4813)
);

O2A1O1Ixp33_ASAP7_75t_L g4814 ( 
.A1(n_4281),
.A2(n_4334),
.B(n_4338),
.C(n_4305),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_3520),
.Y(n_4815)
);

BUFx6f_ASAP7_75t_L g4816 ( 
.A(n_3284),
.Y(n_4816)
);

NOR2x1_ASAP7_75t_L g4817 ( 
.A(n_3657),
.B(n_3516),
.Y(n_4817)
);

BUFx2_ASAP7_75t_L g4818 ( 
.A(n_3823),
.Y(n_4818)
);

OAI21xp5_ASAP7_75t_L g4819 ( 
.A1(n_4383),
.A2(n_4402),
.B(n_4401),
.Y(n_4819)
);

NAND2xp5_ASAP7_75t_L g4820 ( 
.A(n_4227),
.B(n_4236),
.Y(n_4820)
);

O2A1O1Ixp33_ASAP7_75t_L g4821 ( 
.A1(n_4401),
.A2(n_4411),
.B(n_4418),
.C(n_4402),
.Y(n_4821)
);

AOI22x1_ASAP7_75t_L g4822 ( 
.A1(n_3829),
.A2(n_3886),
.B1(n_3269),
.B2(n_3232),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_SL g4823 ( 
.A(n_3276),
.B(n_3315),
.Y(n_4823)
);

NOR2xp33_ASAP7_75t_L g4824 ( 
.A(n_3261),
.B(n_3283),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_SL g4825 ( 
.A(n_3276),
.B(n_3315),
.Y(n_4825)
);

O2A1O1Ixp33_ASAP7_75t_L g4826 ( 
.A1(n_4411),
.A2(n_4489),
.B(n_4508),
.C(n_4418),
.Y(n_4826)
);

A2O1A1Ixp33_ASAP7_75t_L g4827 ( 
.A1(n_4489),
.A2(n_4508),
.B(n_4553),
.C(n_4511),
.Y(n_4827)
);

OAI22xp5_ASAP7_75t_L g4828 ( 
.A1(n_4239),
.A2(n_4255),
.B1(n_4302),
.B2(n_4288),
.Y(n_4828)
);

NOR2x1_ASAP7_75t_L g4829 ( 
.A(n_4718),
.B(n_4719),
.Y(n_4829)
);

A2O1A1Ixp33_ASAP7_75t_L g4830 ( 
.A1(n_4511),
.A2(n_4553),
.B(n_4581),
.C(n_4564),
.Y(n_4830)
);

NOR2xp33_ASAP7_75t_L g4831 ( 
.A(n_3261),
.B(n_3283),
.Y(n_4831)
);

CKINVDCx10_ASAP7_75t_R g4832 ( 
.A(n_3904),
.Y(n_4832)
);

A2O1A1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4564),
.A2(n_4581),
.B(n_4669),
.C(n_4656),
.Y(n_4833)
);

BUFx2_ASAP7_75t_L g4834 ( 
.A(n_3823),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_3639),
.Y(n_4835)
);

O2A1O1Ixp33_ASAP7_75t_L g4836 ( 
.A1(n_4656),
.A2(n_4721),
.B(n_4669),
.C(n_3289),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4238),
.B(n_4244),
.Y(n_4837)
);

CKINVDCx5p33_ASAP7_75t_R g4838 ( 
.A(n_3723),
.Y(n_4838)
);

NOR2xp33_ASAP7_75t_SL g4839 ( 
.A(n_4668),
.B(n_3306),
.Y(n_4839)
);

AOI21x1_ASAP7_75t_L g4840 ( 
.A1(n_3223),
.A2(n_3248),
.B(n_3231),
.Y(n_4840)
);

NOR2xp33_ASAP7_75t_L g4841 ( 
.A(n_3306),
.B(n_3309),
.Y(n_4841)
);

OAI21xp5_ASAP7_75t_L g4842 ( 
.A1(n_4721),
.A2(n_3616),
.B(n_4441),
.Y(n_4842)
);

AOI21xp5_ASAP7_75t_L g4843 ( 
.A1(n_4331),
.A2(n_4501),
.B(n_4362),
.Y(n_4843)
);

OAI21xp5_ASAP7_75t_L g4844 ( 
.A1(n_3616),
.A2(n_4441),
.B(n_4181),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_3639),
.Y(n_4845)
);

BUFx6f_ASAP7_75t_L g4846 ( 
.A(n_3284),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_L g4847 ( 
.A(n_4238),
.B(n_4244),
.Y(n_4847)
);

NOR3xp33_ASAP7_75t_L g4848 ( 
.A(n_4274),
.B(n_4397),
.C(n_4497),
.Y(n_4848)
);

O2A1O1Ixp33_ASAP7_75t_L g4849 ( 
.A1(n_3287),
.A2(n_3289),
.B(n_3300),
.C(n_3293),
.Y(n_4849)
);

AOI21xp5_ASAP7_75t_L g4850 ( 
.A1(n_4331),
.A2(n_4501),
.B(n_4362),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4248),
.B(n_4250),
.Y(n_4851)
);

AO21x1_ASAP7_75t_L g4852 ( 
.A1(n_3248),
.A2(n_4187),
.B(n_4181),
.Y(n_4852)
);

CKINVDCx11_ASAP7_75t_R g4853 ( 
.A(n_4174),
.Y(n_4853)
);

NOR2xp33_ASAP7_75t_L g4854 ( 
.A(n_3309),
.B(n_3317),
.Y(n_4854)
);

AO21x1_ASAP7_75t_L g4855 ( 
.A1(n_4187),
.A2(n_4192),
.B(n_4189),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4248),
.B(n_4250),
.Y(n_4856)
);

OR2x2_ASAP7_75t_L g4857 ( 
.A(n_3229),
.B(n_4162),
.Y(n_4857)
);

OAI21xp33_ASAP7_75t_L g4858 ( 
.A1(n_4320),
.A2(n_4382),
.B(n_4348),
.Y(n_4858)
);

NAND2xp5_ASAP7_75t_L g4859 ( 
.A(n_4253),
.B(n_4254),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4253),
.B(n_4254),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4260),
.B(n_4265),
.Y(n_4861)
);

INVx2_ASAP7_75t_L g4862 ( 
.A(n_3405),
.Y(n_4862)
);

AOI22x1_ASAP7_75t_L g4863 ( 
.A1(n_3829),
.A2(n_3886),
.B1(n_3269),
.B2(n_3232),
.Y(n_4863)
);

AOI21xp5_ASAP7_75t_L g4864 ( 
.A1(n_4331),
.A2(n_4501),
.B(n_4362),
.Y(n_4864)
);

AOI21xp5_ASAP7_75t_L g4865 ( 
.A1(n_4362),
.A2(n_4506),
.B(n_4501),
.Y(n_4865)
);

CKINVDCx20_ASAP7_75t_R g4866 ( 
.A(n_4174),
.Y(n_4866)
);

AOI21xp5_ASAP7_75t_L g4867 ( 
.A1(n_4362),
.A2(n_4506),
.B(n_4501),
.Y(n_4867)
);

AOI21xp5_ASAP7_75t_L g4868 ( 
.A1(n_4506),
.A2(n_4567),
.B(n_4696),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4260),
.B(n_4265),
.Y(n_4869)
);

AOI21xp5_ASAP7_75t_L g4870 ( 
.A1(n_4506),
.A2(n_4567),
.B(n_4696),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4275),
.B(n_4278),
.Y(n_4871)
);

NOR3xp33_ASAP7_75t_L g4872 ( 
.A(n_4274),
.B(n_4397),
.C(n_4497),
.Y(n_4872)
);

AOI21x1_ASAP7_75t_L g4873 ( 
.A1(n_4189),
.A2(n_4202),
.B(n_4192),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4712),
.Y(n_4874)
);

OAI22xp5_ASAP7_75t_L g4875 ( 
.A1(n_4348),
.A2(n_4382),
.B1(n_4560),
.B2(n_4485),
.Y(n_4875)
);

NOR2xp33_ASAP7_75t_L g4876 ( 
.A(n_3317),
.B(n_3319),
.Y(n_4876)
);

O2A1O1Ixp33_ASAP7_75t_L g4877 ( 
.A1(n_3287),
.A2(n_3300),
.B(n_3352),
.C(n_3293),
.Y(n_4877)
);

OAI22xp5_ASAP7_75t_L g4878 ( 
.A1(n_4485),
.A2(n_4560),
.B1(n_4624),
.B2(n_4593),
.Y(n_4878)
);

AOI21xp5_ASAP7_75t_L g4879 ( 
.A1(n_4506),
.A2(n_4567),
.B(n_3222),
.Y(n_4879)
);

HB1xp67_ASAP7_75t_L g4880 ( 
.A(n_3311),
.Y(n_4880)
);

INVx2_ASAP7_75t_L g4881 ( 
.A(n_3418),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4275),
.B(n_4278),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4295),
.B(n_4296),
.Y(n_4883)
);

NOR2xp33_ASAP7_75t_L g4884 ( 
.A(n_3319),
.B(n_3326),
.Y(n_4884)
);

NOR3xp33_ASAP7_75t_L g4885 ( 
.A(n_3324),
.B(n_4325),
.C(n_3366),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4712),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_4295),
.B(n_4296),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_SL g4888 ( 
.A(n_3316),
.B(n_3330),
.Y(n_4888)
);

BUFx4f_ASAP7_75t_L g4889 ( 
.A(n_4186),
.Y(n_4889)
);

AOI21xp5_ASAP7_75t_L g4890 ( 
.A1(n_4506),
.A2(n_4567),
.B(n_3222),
.Y(n_4890)
);

INVx1_ASAP7_75t_L g4891 ( 
.A(n_4713),
.Y(n_4891)
);

AOI21xp5_ASAP7_75t_L g4892 ( 
.A1(n_4506),
.A2(n_4567),
.B(n_4720),
.Y(n_4892)
);

AOI21xp5_ASAP7_75t_L g4893 ( 
.A1(n_4567),
.A2(n_4720),
.B(n_4215),
.Y(n_4893)
);

AOI21xp5_ASAP7_75t_L g4894 ( 
.A1(n_4567),
.A2(n_4215),
.B(n_4206),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4300),
.B(n_4306),
.Y(n_4895)
);

NOR2xp33_ASAP7_75t_L g4896 ( 
.A(n_3326),
.B(n_3344),
.Y(n_4896)
);

AOI21xp5_ASAP7_75t_L g4897 ( 
.A1(n_4202),
.A2(n_4213),
.B(n_4206),
.Y(n_4897)
);

NOR2x1_ASAP7_75t_L g4898 ( 
.A(n_4718),
.B(n_4719),
.Y(n_4898)
);

NAND2xp33_ASAP7_75t_L g4899 ( 
.A(n_3484),
.B(n_4515),
.Y(n_4899)
);

AO21x1_ASAP7_75t_L g4900 ( 
.A1(n_4213),
.A2(n_4240),
.B(n_4219),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4300),
.B(n_4306),
.Y(n_4901)
);

NOR2xp67_ASAP7_75t_L g4902 ( 
.A(n_3760),
.B(n_3518),
.Y(n_4902)
);

NAND2xp5_ASAP7_75t_L g4903 ( 
.A(n_4309),
.B(n_4310),
.Y(n_4903)
);

NOR2xp33_ASAP7_75t_L g4904 ( 
.A(n_3344),
.B(n_3358),
.Y(n_4904)
);

AND2x2_ASAP7_75t_L g4905 ( 
.A(n_3589),
.B(n_3634),
.Y(n_4905)
);

AOI21xp5_ASAP7_75t_L g4906 ( 
.A1(n_4219),
.A2(n_4266),
.B(n_4240),
.Y(n_4906)
);

BUFx6f_ASAP7_75t_L g4907 ( 
.A(n_3284),
.Y(n_4907)
);

AOI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_4266),
.A2(n_4304),
.B(n_4279),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4309),
.B(n_4310),
.Y(n_4909)
);

AOI21xp5_ASAP7_75t_L g4910 ( 
.A1(n_4279),
.A2(n_4336),
.B(n_4304),
.Y(n_4910)
);

INVx1_ASAP7_75t_SL g4911 ( 
.A(n_3758),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_SL g4912 ( 
.A(n_3316),
.B(n_3330),
.Y(n_4912)
);

AOI21xp5_ASAP7_75t_L g4913 ( 
.A1(n_4336),
.A2(n_4353),
.B(n_4345),
.Y(n_4913)
);

AOI21xp5_ASAP7_75t_L g4914 ( 
.A1(n_4345),
.A2(n_4360),
.B(n_4353),
.Y(n_4914)
);

AOI21x1_ASAP7_75t_L g4915 ( 
.A1(n_4360),
.A2(n_4375),
.B(n_4372),
.Y(n_4915)
);

OR2x6_ASAP7_75t_SL g4916 ( 
.A(n_3246),
.B(n_3249),
.Y(n_4916)
);

AND2x2_ASAP7_75t_L g4917 ( 
.A(n_3589),
.B(n_3634),
.Y(n_4917)
);

NOR3xp33_ASAP7_75t_L g4918 ( 
.A(n_3324),
.B(n_4325),
.C(n_3366),
.Y(n_4918)
);

OAI22xp5_ASAP7_75t_L g4919 ( 
.A1(n_4593),
.A2(n_4624),
.B1(n_4654),
.B2(n_3264),
.Y(n_4919)
);

A2O1A1Ixp33_ASAP7_75t_L g4920 ( 
.A1(n_3518),
.A2(n_3368),
.B(n_3370),
.C(n_3358),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_L g4921 ( 
.A(n_4313),
.B(n_4317),
.Y(n_4921)
);

OAI21xp33_ASAP7_75t_L g4922 ( 
.A1(n_4654),
.A2(n_3264),
.B(n_3462),
.Y(n_4922)
);

O2A1O1Ixp33_ASAP7_75t_SL g4923 ( 
.A1(n_3352),
.A2(n_3384),
.B(n_3388),
.C(n_3353),
.Y(n_4923)
);

INVx6_ASAP7_75t_L g4924 ( 
.A(n_3284),
.Y(n_4924)
);

AOI22xp5_ASAP7_75t_L g4925 ( 
.A1(n_4432),
.A2(n_3462),
.B1(n_4648),
.B2(n_3695),
.Y(n_4925)
);

AOI21xp5_ASAP7_75t_L g4926 ( 
.A1(n_4372),
.A2(n_4405),
.B(n_4375),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_SL g4927 ( 
.A(n_3335),
.B(n_3341),
.Y(n_4927)
);

AND2x4_ASAP7_75t_L g4928 ( 
.A(n_3301),
.B(n_3381),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4313),
.B(n_4317),
.Y(n_4929)
);

BUFx3_ASAP7_75t_L g4930 ( 
.A(n_4036),
.Y(n_4930)
);

AOI21xp5_ASAP7_75t_L g4931 ( 
.A1(n_4405),
.A2(n_4439),
.B(n_4433),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_L g4932 ( 
.A(n_4326),
.B(n_4333),
.Y(n_4932)
);

O2A1O1Ixp33_ASAP7_75t_L g4933 ( 
.A1(n_3353),
.A2(n_3388),
.B(n_3384),
.C(n_4709),
.Y(n_4933)
);

CKINVDCx10_ASAP7_75t_R g4934 ( 
.A(n_3904),
.Y(n_4934)
);

OAI21xp5_ASAP7_75t_L g4935 ( 
.A1(n_4433),
.A2(n_4444),
.B(n_4439),
.Y(n_4935)
);

AOI21xp5_ASAP7_75t_L g4936 ( 
.A1(n_4444),
.A2(n_4450),
.B(n_4446),
.Y(n_4936)
);

AOI21x1_ASAP7_75t_L g4937 ( 
.A1(n_4446),
.A2(n_4464),
.B(n_4450),
.Y(n_4937)
);

BUFx4f_ASAP7_75t_L g4938 ( 
.A(n_4186),
.Y(n_4938)
);

INVx3_ASAP7_75t_L g4939 ( 
.A(n_3295),
.Y(n_4939)
);

AOI21xp5_ASAP7_75t_L g4940 ( 
.A1(n_4464),
.A2(n_4494),
.B(n_4465),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4713),
.Y(n_4941)
);

OAI22xp5_ASAP7_75t_SL g4942 ( 
.A1(n_3318),
.A2(n_3354),
.B1(n_3359),
.B2(n_3329),
.Y(n_4942)
);

HB1xp67_ASAP7_75t_L g4943 ( 
.A(n_3311),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4326),
.B(n_4333),
.Y(n_4944)
);

AOI21xp5_ASAP7_75t_L g4945 ( 
.A1(n_4465),
.A2(n_4534),
.B(n_4494),
.Y(n_4945)
);

OAI21xp5_ASAP7_75t_L g4946 ( 
.A1(n_4534),
.A2(n_4542),
.B(n_4537),
.Y(n_4946)
);

O2A1O1Ixp33_ASAP7_75t_L g4947 ( 
.A1(n_4709),
.A2(n_4542),
.B(n_4586),
.C(n_4537),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_SL g4948 ( 
.A(n_3335),
.B(n_3341),
.Y(n_4948)
);

HB1xp67_ASAP7_75t_L g4949 ( 
.A(n_3437),
.Y(n_4949)
);

NOR2xp33_ASAP7_75t_L g4950 ( 
.A(n_3368),
.B(n_3370),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4335),
.B(n_4354),
.Y(n_4951)
);

OAI22xp5_ASAP7_75t_L g4952 ( 
.A1(n_3318),
.A2(n_3329),
.B1(n_3359),
.B2(n_3354),
.Y(n_4952)
);

AO21x1_ASAP7_75t_L g4953 ( 
.A1(n_4586),
.A2(n_4628),
.B(n_4626),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_SL g4954 ( 
.A(n_3362),
.B(n_3391),
.Y(n_4954)
);

AOI21xp5_ASAP7_75t_L g4955 ( 
.A1(n_4626),
.A2(n_4631),
.B(n_4628),
.Y(n_4955)
);

OAI21xp5_ASAP7_75t_L g4956 ( 
.A1(n_4631),
.A2(n_3522),
.B(n_4335),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4354),
.B(n_4359),
.Y(n_4957)
);

AOI21xp5_ASAP7_75t_L g4958 ( 
.A1(n_4711),
.A2(n_4370),
.B(n_4359),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4370),
.B(n_4371),
.Y(n_4959)
);

BUFx3_ASAP7_75t_L g4960 ( 
.A(n_4036),
.Y(n_4960)
);

NOR2xp33_ASAP7_75t_L g4961 ( 
.A(n_3372),
.B(n_3382),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_3418),
.Y(n_4962)
);

AOI21xp5_ASAP7_75t_L g4963 ( 
.A1(n_4711),
.A2(n_4378),
.B(n_4371),
.Y(n_4963)
);

OAI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_3522),
.A2(n_4385),
.B(n_4378),
.Y(n_4964)
);

AOI21x1_ASAP7_75t_L g4965 ( 
.A1(n_3409),
.A2(n_3731),
.B(n_4385),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4394),
.B(n_4400),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4394),
.B(n_4400),
.Y(n_4967)
);

INVx2_ASAP7_75t_L g4968 ( 
.A(n_3418),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4426),
.B(n_4431),
.Y(n_4969)
);

AOI22xp33_ASAP7_75t_L g4970 ( 
.A1(n_3695),
.A2(n_4208),
.B1(n_4399),
.B2(n_4379),
.Y(n_4970)
);

O2A1O1Ixp33_ASAP7_75t_L g4971 ( 
.A1(n_4426),
.A2(n_4431),
.B(n_4449),
.C(n_4442),
.Y(n_4971)
);

AOI22xp5_ASAP7_75t_L g4972 ( 
.A1(n_4432),
.A2(n_3462),
.B1(n_4648),
.B2(n_3483),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4442),
.B(n_4449),
.Y(n_4973)
);

INVx3_ASAP7_75t_L g4974 ( 
.A(n_3295),
.Y(n_4974)
);

NOR2xp33_ASAP7_75t_L g4975 ( 
.A(n_3372),
.B(n_3382),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4452),
.B(n_4467),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4714),
.Y(n_4977)
);

AOI21xp5_ASAP7_75t_L g4978 ( 
.A1(n_4452),
.A2(n_4470),
.B(n_4467),
.Y(n_4978)
);

AOI21x1_ASAP7_75t_L g4979 ( 
.A1(n_3409),
.A2(n_3731),
.B(n_4470),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_SL g4980 ( 
.A(n_3362),
.B(n_3391),
.Y(n_4980)
);

INVx1_ASAP7_75t_L g4981 ( 
.A(n_4715),
.Y(n_4981)
);

OAI21xp5_ASAP7_75t_L g4982 ( 
.A1(n_4474),
.A2(n_4483),
.B(n_4475),
.Y(n_4982)
);

AOI21xp5_ASAP7_75t_L g4983 ( 
.A1(n_4474),
.A2(n_4483),
.B(n_4475),
.Y(n_4983)
);

INVx1_ASAP7_75t_L g4984 ( 
.A(n_3230),
.Y(n_4984)
);

BUFx3_ASAP7_75t_L g4985 ( 
.A(n_4036),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_3230),
.Y(n_4986)
);

AOI21xp5_ASAP7_75t_L g4987 ( 
.A1(n_4698),
.A2(n_4700),
.B(n_4699),
.Y(n_4987)
);

NOR3xp33_ASAP7_75t_L g4988 ( 
.A(n_3463),
.B(n_3857),
.C(n_3694),
.Y(n_4988)
);

NOR2xp67_ASAP7_75t_L g4989 ( 
.A(n_3760),
.B(n_3510),
.Y(n_4989)
);

AOI21x1_ASAP7_75t_L g4990 ( 
.A1(n_4488),
.A2(n_4498),
.B(n_4490),
.Y(n_4990)
);

AOI21xp5_ASAP7_75t_L g4991 ( 
.A1(n_4699),
.A2(n_4700),
.B(n_4490),
.Y(n_4991)
);

NOR3xp33_ASAP7_75t_L g4992 ( 
.A(n_3463),
.B(n_3857),
.C(n_3694),
.Y(n_4992)
);

AOI21xp5_ASAP7_75t_L g4993 ( 
.A1(n_4488),
.A2(n_4518),
.B(n_4498),
.Y(n_4993)
);

AOI21xp5_ASAP7_75t_L g4994 ( 
.A1(n_4518),
.A2(n_4533),
.B(n_4529),
.Y(n_4994)
);

AOI22xp33_ASAP7_75t_L g4995 ( 
.A1(n_4208),
.A2(n_4399),
.B1(n_4563),
.B2(n_4379),
.Y(n_4995)
);

INVx3_ASAP7_75t_L g4996 ( 
.A(n_3295),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4529),
.B(n_4533),
.Y(n_4997)
);

OAI21xp33_ASAP7_75t_L g4998 ( 
.A1(n_4152),
.A2(n_4258),
.B(n_4220),
.Y(n_4998)
);

OAI321xp33_ASAP7_75t_L g4999 ( 
.A1(n_4152),
.A2(n_4258),
.A3(n_4290),
.B1(n_4438),
.B2(n_4423),
.C(n_4220),
.Y(n_4999)
);

A2O1A1Ixp33_ASAP7_75t_L g5000 ( 
.A1(n_3414),
.A2(n_3416),
.B(n_3430),
.C(n_3419),
.Y(n_5000)
);

INVx2_ASAP7_75t_L g5001 ( 
.A(n_3418),
.Y(n_5001)
);

NOR2xp33_ASAP7_75t_L g5002 ( 
.A(n_3414),
.B(n_3416),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4545),
.B(n_4551),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4545),
.B(n_4551),
.Y(n_5004)
);

AOI21xp5_ASAP7_75t_L g5005 ( 
.A1(n_4554),
.A2(n_4580),
.B(n_4572),
.Y(n_5005)
);

INVx2_ASAP7_75t_L g5006 ( 
.A(n_3418),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_SL g5007 ( 
.A(n_4290),
.B(n_4423),
.Y(n_5007)
);

NAND2xp5_ASAP7_75t_SL g5008 ( 
.A(n_4438),
.B(n_4482),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4554),
.B(n_4572),
.Y(n_5009)
);

HB1xp67_ASAP7_75t_L g5010 ( 
.A(n_3437),
.Y(n_5010)
);

BUFx8_ASAP7_75t_SL g5011 ( 
.A(n_4361),
.Y(n_5011)
);

OAI21xp5_ASAP7_75t_L g5012 ( 
.A1(n_4580),
.A2(n_4598),
.B(n_4584),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_SL g5013 ( 
.A(n_4482),
.B(n_4521),
.Y(n_5013)
);

AOI21xp5_ASAP7_75t_L g5014 ( 
.A1(n_4584),
.A2(n_4600),
.B(n_4598),
.Y(n_5014)
);

A2O1A1Ixp33_ASAP7_75t_L g5015 ( 
.A1(n_3419),
.A2(n_3430),
.B(n_3445),
.C(n_3447),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4600),
.B(n_4602),
.Y(n_5016)
);

BUFx6f_ASAP7_75t_L g5017 ( 
.A(n_3284),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_L g5018 ( 
.A(n_4602),
.B(n_4605),
.Y(n_5018)
);

NOR2xp33_ASAP7_75t_L g5019 ( 
.A(n_3445),
.B(n_4521),
.Y(n_5019)
);

AOI21xp5_ASAP7_75t_L g5020 ( 
.A1(n_4605),
.A2(n_4611),
.B(n_4608),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_SL g5021 ( 
.A(n_4528),
.B(n_4531),
.Y(n_5021)
);

NOR2xp33_ASAP7_75t_L g5022 ( 
.A(n_4528),
.B(n_4531),
.Y(n_5022)
);

OAI21x1_ASAP7_75t_L g5023 ( 
.A1(n_3297),
.A2(n_3286),
.B(n_3227),
.Y(n_5023)
);

AOI21xp5_ASAP7_75t_L g5024 ( 
.A1(n_4608),
.A2(n_4617),
.B(n_4611),
.Y(n_5024)
);

OAI21xp5_ASAP7_75t_L g5025 ( 
.A1(n_4617),
.A2(n_4625),
.B(n_4620),
.Y(n_5025)
);

INVx2_ASAP7_75t_L g5026 ( 
.A(n_3418),
.Y(n_5026)
);

NOR2xp33_ASAP7_75t_L g5027 ( 
.A(n_4532),
.B(n_4541),
.Y(n_5027)
);

AO32x1_ASAP7_75t_L g5028 ( 
.A1(n_3235),
.A2(n_4167),
.A3(n_4183),
.B1(n_4171),
.B2(n_4165),
.Y(n_5028)
);

OAI21x1_ASAP7_75t_L g5029 ( 
.A1(n_3297),
.A2(n_3286),
.B(n_3227),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4620),
.B(n_4625),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_4627),
.A2(n_4650),
.B(n_4632),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4627),
.B(n_4632),
.Y(n_5032)
);

INVxp67_ASAP7_75t_L g5033 ( 
.A(n_3909),
.Y(n_5033)
);

OAI21xp33_ASAP7_75t_L g5034 ( 
.A1(n_4532),
.A2(n_4616),
.B(n_4541),
.Y(n_5034)
);

A2O1A1Ixp33_ASAP7_75t_L g5035 ( 
.A1(n_3447),
.A2(n_3483),
.B(n_4618),
.C(n_4616),
.Y(n_5035)
);

INVx2_ASAP7_75t_L g5036 ( 
.A(n_3418),
.Y(n_5036)
);

INVx4_ASAP7_75t_L g5037 ( 
.A(n_4036),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_4650),
.B(n_4674),
.Y(n_5038)
);

NOR2xp67_ASAP7_75t_L g5039 ( 
.A(n_3510),
.B(n_4168),
.Y(n_5039)
);

NAND2xp33_ASAP7_75t_L g5040 ( 
.A(n_3484),
.B(n_4515),
.Y(n_5040)
);

BUFx2_ASAP7_75t_L g5041 ( 
.A(n_3823),
.Y(n_5041)
);

O2A1O1Ixp33_ASAP7_75t_SL g5042 ( 
.A1(n_3953),
.A2(n_3981),
.B(n_4080),
.C(n_3624),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_4674),
.B(n_4694),
.Y(n_5043)
);

INVx2_ASAP7_75t_L g5044 ( 
.A(n_3418),
.Y(n_5044)
);

A2O1A1Ixp33_ASAP7_75t_L g5045 ( 
.A1(n_4618),
.A2(n_4641),
.B(n_4675),
.C(n_4622),
.Y(n_5045)
);

AO22x1_ASAP7_75t_L g5046 ( 
.A1(n_3692),
.A2(n_4036),
.B1(n_4047),
.B2(n_3539),
.Y(n_5046)
);

INVx3_ASAP7_75t_L g5047 ( 
.A(n_3295),
.Y(n_5047)
);

INVxp67_ASAP7_75t_L g5048 ( 
.A(n_3929),
.Y(n_5048)
);

BUFx6f_ASAP7_75t_L g5049 ( 
.A(n_4168),
.Y(n_5049)
);

CKINVDCx14_ASAP7_75t_R g5050 ( 
.A(n_4361),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4715),
.Y(n_5051)
);

AOI21x1_ASAP7_75t_L g5052 ( 
.A1(n_4694),
.A2(n_4698),
.B(n_4697),
.Y(n_5052)
);

NOR2xp33_ASAP7_75t_SL g5053 ( 
.A(n_4668),
.B(n_3741),
.Y(n_5053)
);

AOI21xp5_ASAP7_75t_L g5054 ( 
.A1(n_4697),
.A2(n_4330),
.B(n_3263),
.Y(n_5054)
);

BUFx6f_ASAP7_75t_L g5055 ( 
.A(n_4168),
.Y(n_5055)
);

NOR3xp33_ASAP7_75t_L g5056 ( 
.A(n_3598),
.B(n_4701),
.C(n_3299),
.Y(n_5056)
);

BUFx3_ASAP7_75t_L g5057 ( 
.A(n_4036),
.Y(n_5057)
);

BUFx2_ASAP7_75t_L g5058 ( 
.A(n_3823),
.Y(n_5058)
);

AOI21xp5_ASAP7_75t_L g5059 ( 
.A1(n_4330),
.A2(n_3263),
.B(n_3244),
.Y(n_5059)
);

INVx3_ASAP7_75t_L g5060 ( 
.A(n_3295),
.Y(n_5060)
);

OAI21xp5_ASAP7_75t_L g5061 ( 
.A1(n_3624),
.A2(n_3244),
.B(n_3246),
.Y(n_5061)
);

AND2x2_ASAP7_75t_L g5062 ( 
.A(n_3754),
.B(n_3229),
.Y(n_5062)
);

AND2x2_ASAP7_75t_L g5063 ( 
.A(n_3754),
.B(n_3229),
.Y(n_5063)
);

NOR2xp67_ASAP7_75t_L g5064 ( 
.A(n_4168),
.B(n_4176),
.Y(n_5064)
);

AOI21xp5_ASAP7_75t_L g5065 ( 
.A1(n_3286),
.A2(n_3232),
.B(n_4204),
.Y(n_5065)
);

AOI21xp5_ASAP7_75t_L g5066 ( 
.A1(n_4204),
.A2(n_4512),
.B(n_3279),
.Y(n_5066)
);

INVx2_ASAP7_75t_L g5067 ( 
.A(n_3428),
.Y(n_5067)
);

INVx3_ASAP7_75t_L g5068 ( 
.A(n_3295),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_SL g5069 ( 
.A(n_4622),
.B(n_4641),
.Y(n_5069)
);

AOI21xp5_ASAP7_75t_L g5070 ( 
.A1(n_4204),
.A2(n_4512),
.B(n_3279),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_3285),
.B(n_4016),
.Y(n_5071)
);

O2A1O1Ixp33_ASAP7_75t_L g5072 ( 
.A1(n_3726),
.A2(n_3691),
.B(n_3703),
.C(n_3299),
.Y(n_5072)
);

NAND2xp5_ASAP7_75t_L g5073 ( 
.A(n_3285),
.B(n_4016),
.Y(n_5073)
);

NOR2xp33_ASAP7_75t_L g5074 ( 
.A(n_4675),
.B(n_4717),
.Y(n_5074)
);

INVx1_ASAP7_75t_L g5075 ( 
.A(n_4695),
.Y(n_5075)
);

INVxp67_ASAP7_75t_L g5076 ( 
.A(n_3929),
.Y(n_5076)
);

CKINVDCx6p67_ASAP7_75t_R g5077 ( 
.A(n_4251),
.Y(n_5077)
);

OAI22xp5_ASAP7_75t_L g5078 ( 
.A1(n_4717),
.A2(n_4379),
.B1(n_4399),
.B2(n_4208),
.Y(n_5078)
);

NOR2xp33_ASAP7_75t_R g5079 ( 
.A(n_3644),
.B(n_4644),
.Y(n_5079)
);

AND2x2_ASAP7_75t_L g5080 ( 
.A(n_3754),
.B(n_4162),
.Y(n_5080)
);

AOI21x1_ASAP7_75t_L g5081 ( 
.A1(n_3804),
.A2(n_4167),
.B(n_4165),
.Y(n_5081)
);

BUFx12f_ASAP7_75t_L g5082 ( 
.A(n_4251),
.Y(n_5082)
);

AOI21x1_ASAP7_75t_L g5083 ( 
.A1(n_3804),
.A2(n_4183),
.B(n_4171),
.Y(n_5083)
);

NAND2x1p5_ASAP7_75t_L g5084 ( 
.A(n_4168),
.B(n_4176),
.Y(n_5084)
);

AOI21xp5_ASAP7_75t_L g5085 ( 
.A1(n_4204),
.A2(n_4512),
.B(n_3255),
.Y(n_5085)
);

AOI22xp5_ASAP7_75t_L g5086 ( 
.A1(n_4563),
.A2(n_3269),
.B1(n_3304),
.B2(n_3291),
.Y(n_5086)
);

AOI22xp5_ASAP7_75t_L g5087 ( 
.A1(n_4563),
.A2(n_3291),
.B1(n_3305),
.B2(n_3304),
.Y(n_5087)
);

BUFx6f_ASAP7_75t_L g5088 ( 
.A(n_4168),
.Y(n_5088)
);

OAI22xp5_ASAP7_75t_L g5089 ( 
.A1(n_3780),
.A2(n_3796),
.B1(n_3800),
.B2(n_3784),
.Y(n_5089)
);

NOR2xp33_ASAP7_75t_L g5090 ( 
.A(n_4445),
.B(n_3505),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_L g5091 ( 
.A(n_3598),
.B(n_3552),
.Y(n_5091)
);

OAI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_3249),
.A2(n_3256),
.B(n_3255),
.Y(n_5092)
);

AOI21xp5_ASAP7_75t_L g5093 ( 
.A1(n_4204),
.A2(n_4512),
.B(n_3259),
.Y(n_5093)
);

NOR2xp33_ASAP7_75t_L g5094 ( 
.A(n_4445),
.B(n_3505),
.Y(n_5094)
);

O2A1O1Ixp33_ASAP7_75t_L g5095 ( 
.A1(n_3726),
.A2(n_3691),
.B(n_3703),
.C(n_3302),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4512),
.A2(n_3259),
.B(n_3256),
.Y(n_5096)
);

OAI21xp5_ASAP7_75t_L g5097 ( 
.A1(n_3724),
.A2(n_3308),
.B(n_3305),
.Y(n_5097)
);

NAND2xp5_ASAP7_75t_L g5098 ( 
.A(n_3552),
.B(n_3564),
.Y(n_5098)
);

NAND2x1p5_ASAP7_75t_L g5099 ( 
.A(n_4168),
.B(n_4176),
.Y(n_5099)
);

INVx2_ASAP7_75t_L g5100 ( 
.A(n_3428),
.Y(n_5100)
);

CKINVDCx5p33_ASAP7_75t_R g5101 ( 
.A(n_3727),
.Y(n_5101)
);

OAI21xp5_ASAP7_75t_L g5102 ( 
.A1(n_3724),
.A2(n_3313),
.B(n_3308),
.Y(n_5102)
);

OAI22xp5_ASAP7_75t_L g5103 ( 
.A1(n_3780),
.A2(n_3796),
.B1(n_3800),
.B2(n_3784),
.Y(n_5103)
);

AND2x4_ASAP7_75t_L g5104 ( 
.A(n_3301),
.B(n_3381),
.Y(n_5104)
);

OAI21x1_ASAP7_75t_L g5105 ( 
.A1(n_3297),
.A2(n_4373),
.B(n_3227),
.Y(n_5105)
);

AOI21xp5_ASAP7_75t_L g5106 ( 
.A1(n_3550),
.A2(n_3672),
.B(n_3227),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_L g5107 ( 
.A(n_3564),
.B(n_3573),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_SL g5108 ( 
.A(n_3543),
.B(n_3560),
.Y(n_5108)
);

AOI21xp5_ASAP7_75t_L g5109 ( 
.A1(n_3550),
.A2(n_3672),
.B(n_4373),
.Y(n_5109)
);

AOI21xp5_ASAP7_75t_L g5110 ( 
.A1(n_4373),
.A2(n_4422),
.B(n_4419),
.Y(n_5110)
);

O2A1O1Ixp33_ASAP7_75t_L g5111 ( 
.A1(n_3280),
.A2(n_3302),
.B(n_4271),
.C(n_4224),
.Y(n_5111)
);

AOI21xp5_ASAP7_75t_L g5112 ( 
.A1(n_4373),
.A2(n_4422),
.B(n_4419),
.Y(n_5112)
);

OAI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_3313),
.A2(n_3325),
.B(n_3320),
.Y(n_5113)
);

BUFx6f_ASAP7_75t_L g5114 ( 
.A(n_4168),
.Y(n_5114)
);

AOI21xp5_ASAP7_75t_L g5115 ( 
.A1(n_4419),
.A2(n_4472),
.B(n_4422),
.Y(n_5115)
);

AOI21xp5_ASAP7_75t_L g5116 ( 
.A1(n_4419),
.A2(n_4472),
.B(n_4422),
.Y(n_5116)
);

NAND2xp5_ASAP7_75t_SL g5117 ( 
.A(n_3543),
.B(n_3560),
.Y(n_5117)
);

AOI21xp5_ASAP7_75t_L g5118 ( 
.A1(n_4472),
.A2(n_4591),
.B(n_4570),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_L g5119 ( 
.A(n_3573),
.B(n_3632),
.Y(n_5119)
);

AOI22xp33_ASAP7_75t_L g5120 ( 
.A1(n_3692),
.A2(n_3383),
.B1(n_3336),
.B2(n_3325),
.Y(n_5120)
);

NAND3xp33_ASAP7_75t_L g5121 ( 
.A(n_3715),
.B(n_3502),
.C(n_4210),
.Y(n_5121)
);

INVx2_ASAP7_75t_SL g5122 ( 
.A(n_3539),
.Y(n_5122)
);

BUFx6f_ASAP7_75t_L g5123 ( 
.A(n_4176),
.Y(n_5123)
);

BUFx6f_ASAP7_75t_L g5124 ( 
.A(n_4176),
.Y(n_5124)
);

AOI21xp5_ASAP7_75t_L g5125 ( 
.A1(n_4472),
.A2(n_4591),
.B(n_4570),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_L g5126 ( 
.A(n_3632),
.B(n_3652),
.Y(n_5126)
);

O2A1O1Ixp33_ASAP7_75t_L g5127 ( 
.A1(n_3280),
.A2(n_4224),
.B(n_4407),
.C(n_4271),
.Y(n_5127)
);

AOI21xp5_ASAP7_75t_L g5128 ( 
.A1(n_4570),
.A2(n_4591),
.B(n_3297),
.Y(n_5128)
);

NOR2xp33_ASAP7_75t_L g5129 ( 
.A(n_3696),
.B(n_4084),
.Y(n_5129)
);

OAI21xp5_ASAP7_75t_L g5130 ( 
.A1(n_3320),
.A2(n_3336),
.B(n_3334),
.Y(n_5130)
);

NOR2xp33_ASAP7_75t_L g5131 ( 
.A(n_4084),
.B(n_3716),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_3652),
.B(n_3676),
.Y(n_5132)
);

O2A1O1Ixp33_ASAP7_75t_L g5133 ( 
.A1(n_4407),
.A2(n_4535),
.B(n_4647),
.C(n_4573),
.Y(n_5133)
);

OR2x6_ASAP7_75t_SL g5134 ( 
.A(n_3334),
.B(n_3348),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_3676),
.B(n_4164),
.Y(n_5135)
);

NAND2x1p5_ASAP7_75t_L g5136 ( 
.A(n_4176),
.B(n_4193),
.Y(n_5136)
);

OA22x2_ASAP7_75t_L g5137 ( 
.A1(n_3903),
.A2(n_3986),
.B1(n_3970),
.B2(n_3814),
.Y(n_5137)
);

BUFx4f_ASAP7_75t_L g5138 ( 
.A(n_4186),
.Y(n_5138)
);

AOI21xp5_ASAP7_75t_L g5139 ( 
.A1(n_4570),
.A2(n_4591),
.B(n_3704),
.Y(n_5139)
);

INVx2_ASAP7_75t_L g5140 ( 
.A(n_3428),
.Y(n_5140)
);

AOI21xp5_ASAP7_75t_L g5141 ( 
.A1(n_3704),
.A2(n_3814),
.B(n_4164),
.Y(n_5141)
);

NOR2xp33_ASAP7_75t_L g5142 ( 
.A(n_3716),
.B(n_3742),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_SL g5143 ( 
.A(n_3596),
.B(n_3600),
.Y(n_5143)
);

OAI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_3801),
.A2(n_3807),
.B1(n_3811),
.B2(n_3806),
.Y(n_5144)
);

NOR2xp33_ASAP7_75t_L g5145 ( 
.A(n_3742),
.B(n_3753),
.Y(n_5145)
);

AOI22xp33_ASAP7_75t_SL g5146 ( 
.A1(n_3348),
.A2(n_3355),
.B1(n_3365),
.B2(n_3350),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_4714),
.Y(n_5147)
);

AND2x6_ASAP7_75t_L g5148 ( 
.A(n_3254),
.B(n_3274),
.Y(n_5148)
);

INVx1_ASAP7_75t_SL g5149 ( 
.A(n_3601),
.Y(n_5149)
);

NAND2xp5_ASAP7_75t_L g5150 ( 
.A(n_4164),
.B(n_4276),
.Y(n_5150)
);

BUFx2_ASAP7_75t_L g5151 ( 
.A(n_3449),
.Y(n_5151)
);

BUFx6f_ASAP7_75t_L g5152 ( 
.A(n_4176),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_4184),
.Y(n_5153)
);

NOR2xp33_ASAP7_75t_L g5154 ( 
.A(n_3753),
.B(n_3766),
.Y(n_5154)
);

NAND2xp5_ASAP7_75t_SL g5155 ( 
.A(n_3596),
.B(n_3600),
.Y(n_5155)
);

INVx1_ASAP7_75t_SL g5156 ( 
.A(n_3601),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_4276),
.B(n_4280),
.Y(n_5157)
);

AOI21xp5_ASAP7_75t_L g5158 ( 
.A1(n_4276),
.A2(n_4349),
.B(n_4280),
.Y(n_5158)
);

AOI33xp33_ASAP7_75t_L g5159 ( 
.A1(n_3791),
.A2(n_3782),
.A3(n_3838),
.B1(n_4059),
.B2(n_3235),
.B3(n_4121),
.Y(n_5159)
);

A2O1A1Ixp33_ASAP7_75t_L g5160 ( 
.A1(n_4210),
.A2(n_4216),
.B(n_4282),
.C(n_4235),
.Y(n_5160)
);

AOI22x1_ASAP7_75t_L g5161 ( 
.A1(n_4177),
.A2(n_4395),
.B1(n_4429),
.B2(n_4301),
.Y(n_5161)
);

INVx2_ASAP7_75t_L g5162 ( 
.A(n_3428),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_4280),
.B(n_4349),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_L g5164 ( 
.A(n_4349),
.B(n_4409),
.Y(n_5164)
);

AOI21xp5_ASAP7_75t_L g5165 ( 
.A1(n_4409),
.A2(n_4491),
.B(n_4478),
.Y(n_5165)
);

AOI21xp5_ASAP7_75t_L g5166 ( 
.A1(n_4409),
.A2(n_4491),
.B(n_4478),
.Y(n_5166)
);

AOI21xp5_ASAP7_75t_L g5167 ( 
.A1(n_4478),
.A2(n_4556),
.B(n_4491),
.Y(n_5167)
);

NAND2xp5_ASAP7_75t_L g5168 ( 
.A(n_4556),
.B(n_4558),
.Y(n_5168)
);

O2A1O1Ixp33_ASAP7_75t_L g5169 ( 
.A1(n_4535),
.A2(n_4647),
.B(n_4701),
.C(n_4573),
.Y(n_5169)
);

OAI22xp5_ASAP7_75t_L g5170 ( 
.A1(n_3801),
.A2(n_3807),
.B1(n_3811),
.B2(n_3806),
.Y(n_5170)
);

CKINVDCx11_ASAP7_75t_R g5171 ( 
.A(n_4644),
.Y(n_5171)
);

NOR2xp33_ASAP7_75t_L g5172 ( 
.A(n_3766),
.B(n_3771),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_SL g5173 ( 
.A(n_3635),
.B(n_3658),
.Y(n_5173)
);

AOI22xp33_ASAP7_75t_L g5174 ( 
.A1(n_3692),
.A2(n_3383),
.B1(n_3355),
.B2(n_3365),
.Y(n_5174)
);

OAI22xp5_ASAP7_75t_L g5175 ( 
.A1(n_3815),
.A2(n_3658),
.B1(n_3666),
.B2(n_3635),
.Y(n_5175)
);

NOR2x1_ASAP7_75t_R g5176 ( 
.A(n_3415),
.B(n_3457),
.Y(n_5176)
);

O2A1O1Ixp5_ASAP7_75t_L g5177 ( 
.A1(n_3776),
.A2(n_3375),
.B(n_3377),
.C(n_3350),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_SL g5178 ( 
.A(n_3666),
.B(n_3682),
.Y(n_5178)
);

OAI22xp5_ASAP7_75t_L g5179 ( 
.A1(n_3815),
.A2(n_3682),
.B1(n_3378),
.B2(n_3379),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_4184),
.Y(n_5180)
);

O2A1O1Ixp33_ASAP7_75t_L g5181 ( 
.A1(n_3375),
.A2(n_3379),
.B(n_3392),
.C(n_3377),
.Y(n_5181)
);

BUFx2_ASAP7_75t_L g5182 ( 
.A(n_3449),
.Y(n_5182)
);

NOR2xp33_ASAP7_75t_L g5183 ( 
.A(n_3771),
.B(n_4048),
.Y(n_5183)
);

AND2x2_ASAP7_75t_L g5184 ( 
.A(n_4162),
.B(n_4203),
.Y(n_5184)
);

INVx2_ASAP7_75t_L g5185 ( 
.A(n_3428),
.Y(n_5185)
);

AOI21xp5_ASAP7_75t_L g5186 ( 
.A1(n_4556),
.A2(n_4565),
.B(n_4558),
.Y(n_5186)
);

AOI21xp5_ASAP7_75t_L g5187 ( 
.A1(n_4558),
.A2(n_4589),
.B(n_4565),
.Y(n_5187)
);

NOR3xp33_ASAP7_75t_L g5188 ( 
.A(n_4042),
.B(n_3767),
.C(n_4055),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_4565),
.B(n_4589),
.Y(n_5189)
);

AOI21xp5_ASAP7_75t_L g5190 ( 
.A1(n_4589),
.A2(n_4704),
.B(n_4603),
.Y(n_5190)
);

BUFx4f_ASAP7_75t_L g5191 ( 
.A(n_4186),
.Y(n_5191)
);

AOI21xp5_ASAP7_75t_L g5192 ( 
.A1(n_4603),
.A2(n_4704),
.B(n_3919),
.Y(n_5192)
);

BUFx6f_ASAP7_75t_L g5193 ( 
.A(n_4176),
.Y(n_5193)
);

OAI21xp5_ASAP7_75t_L g5194 ( 
.A1(n_3378),
.A2(n_3393),
.B(n_3392),
.Y(n_5194)
);

AOI21xp5_ASAP7_75t_L g5195 ( 
.A1(n_4603),
.A2(n_4704),
.B(n_3919),
.Y(n_5195)
);

OAI21xp5_ASAP7_75t_L g5196 ( 
.A1(n_3393),
.A2(n_3402),
.B(n_3473),
.Y(n_5196)
);

INVx2_ASAP7_75t_L g5197 ( 
.A(n_3428),
.Y(n_5197)
);

OAI21xp5_ASAP7_75t_L g5198 ( 
.A1(n_3402),
.A2(n_3476),
.B(n_3473),
.Y(n_5198)
);

AOI21xp5_ASAP7_75t_L g5199 ( 
.A1(n_3916),
.A2(n_3943),
.B(n_4193),
.Y(n_5199)
);

INVx1_ASAP7_75t_L g5200 ( 
.A(n_4691),
.Y(n_5200)
);

NAND2xp5_ASAP7_75t_SL g5201 ( 
.A(n_3502),
.B(n_3728),
.Y(n_5201)
);

OAI21xp5_ASAP7_75t_L g5202 ( 
.A1(n_3476),
.A2(n_3528),
.B(n_3486),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_3403),
.B(n_3710),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_SL g5204 ( 
.A(n_3728),
.B(n_3976),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_4695),
.Y(n_5205)
);

AOI21xp5_ASAP7_75t_L g5206 ( 
.A1(n_3916),
.A2(n_3943),
.B(n_4193),
.Y(n_5206)
);

AOI22x1_ASAP7_75t_L g5207 ( 
.A1(n_4177),
.A2(n_4395),
.B1(n_4429),
.B2(n_4301),
.Y(n_5207)
);

O2A1O1Ixp33_ASAP7_75t_SL g5208 ( 
.A1(n_4044),
.A2(n_4042),
.B(n_4135),
.C(n_4055),
.Y(n_5208)
);

AOI21xp5_ASAP7_75t_L g5209 ( 
.A1(n_4193),
.A2(n_4261),
.B(n_4217),
.Y(n_5209)
);

AOI21xp5_ASAP7_75t_L g5210 ( 
.A1(n_4193),
.A2(n_4261),
.B(n_4217),
.Y(n_5210)
);

NOR2xp33_ASAP7_75t_L g5211 ( 
.A(n_4048),
.B(n_3946),
.Y(n_5211)
);

NAND2xp5_ASAP7_75t_L g5212 ( 
.A(n_3403),
.B(n_3710),
.Y(n_5212)
);

AOI21xp5_ASAP7_75t_L g5213 ( 
.A1(n_4193),
.A2(n_4261),
.B(n_4217),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_4687),
.Y(n_5214)
);

NOR2xp33_ASAP7_75t_SL g5215 ( 
.A(n_3741),
.B(n_4526),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_3713),
.B(n_3720),
.Y(n_5216)
);

NAND2xp5_ASAP7_75t_L g5217 ( 
.A(n_3713),
.B(n_3720),
.Y(n_5217)
);

AOI21x1_ASAP7_75t_L g5218 ( 
.A1(n_4188),
.A2(n_4191),
.B(n_4190),
.Y(n_5218)
);

BUFx2_ASAP7_75t_L g5219 ( 
.A(n_3449),
.Y(n_5219)
);

O2A1O1Ixp33_ASAP7_75t_L g5220 ( 
.A1(n_3485),
.A2(n_3554),
.B(n_3556),
.C(n_3495),
.Y(n_5220)
);

AOI21xp5_ASAP7_75t_L g5221 ( 
.A1(n_4193),
.A2(n_4261),
.B(n_4217),
.Y(n_5221)
);

INVx3_ASAP7_75t_L g5222 ( 
.A(n_3349),
.Y(n_5222)
);

OAI21xp5_ASAP7_75t_L g5223 ( 
.A1(n_3486),
.A2(n_3561),
.B(n_3528),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_SL g5224 ( 
.A(n_3976),
.B(n_3715),
.Y(n_5224)
);

AND2x4_ASAP7_75t_L g5225 ( 
.A(n_3301),
.B(n_3381),
.Y(n_5225)
);

NOR2xp33_ASAP7_75t_L g5226 ( 
.A(n_3946),
.B(n_3812),
.Y(n_5226)
);

O2A1O1Ixp33_ASAP7_75t_L g5227 ( 
.A1(n_3485),
.A2(n_3554),
.B(n_3556),
.C(n_3495),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_3733),
.B(n_3735),
.Y(n_5228)
);

O2A1O1Ixp33_ASAP7_75t_SL g5229 ( 
.A1(n_4044),
.A2(n_4135),
.B(n_3772),
.C(n_3745),
.Y(n_5229)
);

AOI21xp5_ASAP7_75t_L g5230 ( 
.A1(n_4193),
.A2(n_4261),
.B(n_4217),
.Y(n_5230)
);

AOI21xp5_ASAP7_75t_L g5231 ( 
.A1(n_4217),
.A2(n_4380),
.B(n_4261),
.Y(n_5231)
);

AOI21xp5_ASAP7_75t_L g5232 ( 
.A1(n_4217),
.A2(n_4380),
.B(n_4261),
.Y(n_5232)
);

AOI21x1_ASAP7_75t_L g5233 ( 
.A1(n_4188),
.A2(n_4191),
.B(n_4190),
.Y(n_5233)
);

AOI22xp5_ASAP7_75t_L g5234 ( 
.A1(n_4062),
.A2(n_3903),
.B1(n_3692),
.B2(n_4216),
.Y(n_5234)
);

INVx11_ASAP7_75t_L g5235 ( 
.A(n_3626),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_4194),
.Y(n_5236)
);

NOR2xp33_ASAP7_75t_L g5237 ( 
.A(n_3812),
.B(n_3699),
.Y(n_5237)
);

AOI21xp5_ASAP7_75t_L g5238 ( 
.A1(n_4217),
.A2(n_4380),
.B(n_4261),
.Y(n_5238)
);

AOI21xp5_ASAP7_75t_L g5239 ( 
.A1(n_4380),
.A2(n_4652),
.B(n_4527),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_4194),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_L g5241 ( 
.A(n_3733),
.B(n_3735),
.Y(n_5241)
);

BUFx6f_ASAP7_75t_L g5242 ( 
.A(n_4380),
.Y(n_5242)
);

BUFx2_ASAP7_75t_L g5243 ( 
.A(n_3361),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_4203),
.B(n_4273),
.Y(n_5244)
);

A2O1A1Ixp33_ASAP7_75t_L g5245 ( 
.A1(n_4235),
.A2(n_4339),
.B(n_4456),
.C(n_4282),
.Y(n_5245)
);

INVx2_ASAP7_75t_L g5246 ( 
.A(n_3428),
.Y(n_5246)
);

AOI22x1_ASAP7_75t_L g5247 ( 
.A1(n_4466),
.A2(n_3569),
.B1(n_3588),
.B2(n_4064),
.Y(n_5247)
);

NAND2xp5_ASAP7_75t_L g5248 ( 
.A(n_3744),
.B(n_3569),
.Y(n_5248)
);

OAI21xp5_ASAP7_75t_L g5249 ( 
.A1(n_3561),
.A2(n_3617),
.B(n_3567),
.Y(n_5249)
);

AO21x1_ASAP7_75t_L g5250 ( 
.A1(n_3776),
.A2(n_3763),
.B(n_3588),
.Y(n_5250)
);

OR2x6_ASAP7_75t_L g5251 ( 
.A(n_4186),
.B(n_3270),
.Y(n_5251)
);

INVx2_ASAP7_75t_L g5252 ( 
.A(n_3428),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_3744),
.B(n_3973),
.Y(n_5253)
);

INVx5_ASAP7_75t_L g5254 ( 
.A(n_4380),
.Y(n_5254)
);

BUFx6f_ASAP7_75t_L g5255 ( 
.A(n_4380),
.Y(n_5255)
);

INVx2_ASAP7_75t_L g5256 ( 
.A(n_3521),
.Y(n_5256)
);

AOI21xp5_ASAP7_75t_L g5257 ( 
.A1(n_4380),
.A2(n_4652),
.B(n_4527),
.Y(n_5257)
);

AOI21xp5_ASAP7_75t_L g5258 ( 
.A1(n_4527),
.A2(n_4658),
.B(n_4652),
.Y(n_5258)
);

BUFx8_ASAP7_75t_L g5259 ( 
.A(n_4350),
.Y(n_5259)
);

AOI21x1_ASAP7_75t_L g5260 ( 
.A1(n_4195),
.A2(n_4200),
.B(n_4198),
.Y(n_5260)
);

INVx2_ASAP7_75t_SL g5261 ( 
.A(n_3539),
.Y(n_5261)
);

AOI21xp5_ASAP7_75t_L g5262 ( 
.A1(n_4527),
.A2(n_4658),
.B(n_4652),
.Y(n_5262)
);

AOI21xp5_ASAP7_75t_L g5263 ( 
.A1(n_4527),
.A2(n_4658),
.B(n_4652),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_SL g5264 ( 
.A(n_3971),
.B(n_3709),
.Y(n_5264)
);

INVx6_ASAP7_75t_L g5265 ( 
.A(n_4527),
.Y(n_5265)
);

INVx2_ASAP7_75t_L g5266 ( 
.A(n_3521),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_SL g5267 ( 
.A(n_3971),
.B(n_3709),
.Y(n_5267)
);

OAI22xp33_ASAP7_75t_L g5268 ( 
.A1(n_3623),
.A2(n_3637),
.B1(n_3911),
.B2(n_3970),
.Y(n_5268)
);

AOI21xp5_ASAP7_75t_L g5269 ( 
.A1(n_4527),
.A2(n_4658),
.B(n_4652),
.Y(n_5269)
);

INVx8_ASAP7_75t_L g5270 ( 
.A(n_4526),
.Y(n_5270)
);

AOI21xp5_ASAP7_75t_L g5271 ( 
.A1(n_4527),
.A2(n_4658),
.B(n_4652),
.Y(n_5271)
);

OAI22xp5_ASAP7_75t_L g5272 ( 
.A1(n_3347),
.A2(n_3424),
.B1(n_3453),
.B2(n_3451),
.Y(n_5272)
);

O2A1O1Ixp33_ASAP7_75t_L g5273 ( 
.A1(n_3558),
.A2(n_3593),
.B(n_3603),
.C(n_3565),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_3973),
.B(n_3992),
.Y(n_5274)
);

NOR2xp33_ASAP7_75t_L g5275 ( 
.A(n_3699),
.B(n_3899),
.Y(n_5275)
);

AND2x4_ASAP7_75t_SL g5276 ( 
.A(n_3270),
.B(n_3314),
.Y(n_5276)
);

OAI21xp5_ASAP7_75t_L g5277 ( 
.A1(n_3567),
.A2(n_3618),
.B(n_3617),
.Y(n_5277)
);

OR2x2_ASAP7_75t_SL g5278 ( 
.A(n_4134),
.B(n_3349),
.Y(n_5278)
);

NAND2xp5_ASAP7_75t_SL g5279 ( 
.A(n_3424),
.B(n_3451),
.Y(n_5279)
);

AO21x1_ASAP7_75t_L g5280 ( 
.A1(n_3763),
.A2(n_3750),
.B(n_3896),
.Y(n_5280)
);

OAI21x1_ASAP7_75t_L g5281 ( 
.A1(n_4686),
.A2(n_4692),
.B(n_4689),
.Y(n_5281)
);

AOI21xp5_ASAP7_75t_L g5282 ( 
.A1(n_4652),
.A2(n_4658),
.B(n_3314),
.Y(n_5282)
);

AOI22xp33_ASAP7_75t_L g5283 ( 
.A1(n_3692),
.A2(n_4062),
.B1(n_3398),
.B2(n_3772),
.Y(n_5283)
);

OAI21x1_ASAP7_75t_L g5284 ( 
.A1(n_4689),
.A2(n_4693),
.B(n_4692),
.Y(n_5284)
);

AOI21xp5_ASAP7_75t_L g5285 ( 
.A1(n_4658),
.A2(n_3314),
.B(n_3270),
.Y(n_5285)
);

HB1xp67_ASAP7_75t_L g5286 ( 
.A(n_3260),
.Y(n_5286)
);

AOI21x1_ASAP7_75t_L g5287 ( 
.A1(n_4195),
.A2(n_4200),
.B(n_4198),
.Y(n_5287)
);

OAI22xp5_ASAP7_75t_L g5288 ( 
.A1(n_3347),
.A2(n_3453),
.B1(n_3469),
.B2(n_3458),
.Y(n_5288)
);

NAND2xp5_ASAP7_75t_L g5289 ( 
.A(n_3973),
.B(n_3992),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_SL g5290 ( 
.A(n_3458),
.B(n_3469),
.Y(n_5290)
);

OR2x6_ASAP7_75t_L g5291 ( 
.A(n_3270),
.B(n_3314),
.Y(n_5291)
);

INVx1_ASAP7_75t_SL g5292 ( 
.A(n_4175),
.Y(n_5292)
);

NOR2xp67_ASAP7_75t_L g5293 ( 
.A(n_4658),
.B(n_3361),
.Y(n_5293)
);

OAI21x1_ASAP7_75t_L g5294 ( 
.A1(n_4294),
.A2(n_4341),
.B(n_4340),
.Y(n_5294)
);

OA22x2_ASAP7_75t_L g5295 ( 
.A1(n_3986),
.A2(n_3730),
.B1(n_3745),
.B2(n_3759),
.Y(n_5295)
);

AOI21xp5_ASAP7_75t_L g5296 ( 
.A1(n_3270),
.A2(n_4182),
.B(n_3314),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_3992),
.B(n_3996),
.Y(n_5297)
);

AOI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_4182),
.A2(n_4314),
.B(n_4246),
.Y(n_5298)
);

NAND2xp5_ASAP7_75t_L g5299 ( 
.A(n_3996),
.B(n_4003),
.Y(n_5299)
);

INVxp67_ASAP7_75t_SL g5300 ( 
.A(n_3268),
.Y(n_5300)
);

AOI21xp5_ASAP7_75t_L g5301 ( 
.A1(n_4182),
.A2(n_4314),
.B(n_4246),
.Y(n_5301)
);

AND2x2_ASAP7_75t_L g5302 ( 
.A(n_4203),
.B(n_4273),
.Y(n_5302)
);

NAND2xp5_ASAP7_75t_L g5303 ( 
.A(n_3996),
.B(n_4003),
.Y(n_5303)
);

NOR2x1p5_ASAP7_75t_L g5304 ( 
.A(n_4134),
.B(n_3541),
.Y(n_5304)
);

AOI21xp5_ASAP7_75t_L g5305 ( 
.A1(n_4182),
.A2(n_4314),
.B(n_4246),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_SL g5306 ( 
.A(n_3477),
.B(n_3482),
.Y(n_5306)
);

BUFx6f_ASAP7_75t_L g5307 ( 
.A(n_3349),
.Y(n_5307)
);

AND2x2_ASAP7_75t_L g5308 ( 
.A(n_4273),
.B(n_4412),
.Y(n_5308)
);

NAND2xp5_ASAP7_75t_L g5309 ( 
.A(n_4003),
.B(n_4007),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_4007),
.B(n_4008),
.Y(n_5310)
);

BUFx2_ASAP7_75t_L g5311 ( 
.A(n_3361),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_4207),
.Y(n_5312)
);

AOI22xp33_ASAP7_75t_L g5313 ( 
.A1(n_3692),
.A2(n_3398),
.B1(n_3546),
.B2(n_3541),
.Y(n_5313)
);

NAND2xp5_ASAP7_75t_L g5314 ( 
.A(n_4007),
.B(n_4008),
.Y(n_5314)
);

NAND3xp33_ASAP7_75t_L g5315 ( 
.A(n_4339),
.B(n_4645),
.C(n_4456),
.Y(n_5315)
);

O2A1O1Ixp33_ASAP7_75t_SL g5316 ( 
.A1(n_3706),
.A2(n_4144),
.B(n_3565),
.C(n_3593),
.Y(n_5316)
);

NOR2xp67_ASAP7_75t_L g5317 ( 
.A(n_3539),
.B(n_4207),
.Y(n_5317)
);

AOI21x1_ASAP7_75t_L g5318 ( 
.A1(n_4230),
.A2(n_4241),
.B(n_4234),
.Y(n_5318)
);

AOI21x1_ASAP7_75t_L g5319 ( 
.A1(n_4230),
.A2(n_4241),
.B(n_4234),
.Y(n_5319)
);

O2A1O1Ixp5_ASAP7_75t_L g5320 ( 
.A1(n_4242),
.A2(n_4268),
.B(n_4269),
.C(n_4245),
.Y(n_5320)
);

INVx3_ASAP7_75t_SL g5321 ( 
.A(n_4104),
.Y(n_5321)
);

NAND2xp5_ASAP7_75t_L g5322 ( 
.A(n_4008),
.B(n_4015),
.Y(n_5322)
);

NOR2xp67_ASAP7_75t_L g5323 ( 
.A(n_3539),
.B(n_4242),
.Y(n_5323)
);

AOI21xp5_ASAP7_75t_L g5324 ( 
.A1(n_4182),
.A2(n_4314),
.B(n_4246),
.Y(n_5324)
);

OAI21xp5_ASAP7_75t_L g5325 ( 
.A1(n_3618),
.A2(n_3640),
.B(n_3853),
.Y(n_5325)
);

AOI21xp5_ASAP7_75t_L g5326 ( 
.A1(n_4246),
.A2(n_4319),
.B(n_4314),
.Y(n_5326)
);

BUFx2_ASAP7_75t_L g5327 ( 
.A(n_3272),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_4015),
.B(n_3460),
.Y(n_5328)
);

INVx2_ASAP7_75t_SL g5329 ( 
.A(n_3539),
.Y(n_5329)
);

NAND2xp5_ASAP7_75t_L g5330 ( 
.A(n_4015),
.B(n_3460),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_3460),
.B(n_3477),
.Y(n_5331)
);

AOI21xp5_ASAP7_75t_L g5332 ( 
.A1(n_4319),
.A2(n_4517),
.B(n_4461),
.Y(n_5332)
);

NAND2xp5_ASAP7_75t_SL g5333 ( 
.A(n_3482),
.B(n_3488),
.Y(n_5333)
);

NOR2xp33_ASAP7_75t_SL g5334 ( 
.A(n_4526),
.B(n_4350),
.Y(n_5334)
);

NAND2xp5_ASAP7_75t_L g5335 ( 
.A(n_3488),
.B(n_3490),
.Y(n_5335)
);

INVx6_ASAP7_75t_L g5336 ( 
.A(n_4319),
.Y(n_5336)
);

INVx4_ASAP7_75t_L g5337 ( 
.A(n_4047),
.Y(n_5337)
);

O2A1O1Ixp33_ASAP7_75t_L g5338 ( 
.A1(n_3558),
.A2(n_3621),
.B(n_3622),
.C(n_3603),
.Y(n_5338)
);

AND2x2_ASAP7_75t_L g5339 ( 
.A(n_4412),
.B(n_4471),
.Y(n_5339)
);

NAND2xp5_ASAP7_75t_L g5340 ( 
.A(n_3490),
.B(n_3498),
.Y(n_5340)
);

OA22x2_ASAP7_75t_L g5341 ( 
.A1(n_3730),
.A2(n_3759),
.B1(n_3911),
.B2(n_3840),
.Y(n_5341)
);

NOR2xp33_ASAP7_75t_L g5342 ( 
.A(n_3899),
.B(n_4091),
.Y(n_5342)
);

BUFx3_ASAP7_75t_L g5343 ( 
.A(n_4047),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_SL g5344 ( 
.A(n_3498),
.B(n_3500),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_SL g5345 ( 
.A(n_3500),
.B(n_3507),
.Y(n_5345)
);

INVx2_ASAP7_75t_L g5346 ( 
.A(n_3521),
.Y(n_5346)
);

O2A1O1Ixp33_ASAP7_75t_SL g5347 ( 
.A1(n_3706),
.A2(n_4144),
.B(n_3622),
.C(n_3625),
.Y(n_5347)
);

AOI21xp5_ASAP7_75t_L g5348 ( 
.A1(n_4319),
.A2(n_4517),
.B(n_4461),
.Y(n_5348)
);

AOI21xp5_ASAP7_75t_L g5349 ( 
.A1(n_4319),
.A2(n_4517),
.B(n_4461),
.Y(n_5349)
);

AOI21xp5_ASAP7_75t_L g5350 ( 
.A1(n_4461),
.A2(n_4568),
.B(n_4517),
.Y(n_5350)
);

A2O1A1Ixp33_ASAP7_75t_L g5351 ( 
.A1(n_4645),
.A2(n_4649),
.B(n_4661),
.C(n_4028),
.Y(n_5351)
);

NAND2xp5_ASAP7_75t_L g5352 ( 
.A(n_3507),
.B(n_3511),
.Y(n_5352)
);

OAI22xp5_ASAP7_75t_L g5353 ( 
.A1(n_3347),
.A2(n_3515),
.B1(n_3517),
.B2(n_3511),
.Y(n_5353)
);

AOI21xp5_ASAP7_75t_L g5354 ( 
.A1(n_4461),
.A2(n_4568),
.B(n_4517),
.Y(n_5354)
);

NAND3xp33_ASAP7_75t_L g5355 ( 
.A(n_4649),
.B(n_4661),
.C(n_3465),
.Y(n_5355)
);

NOR2xp33_ASAP7_75t_L g5356 ( 
.A(n_4091),
.B(n_3623),
.Y(n_5356)
);

NAND2xp5_ASAP7_75t_L g5357 ( 
.A(n_3515),
.B(n_3517),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_4688),
.Y(n_5358)
);

OR2x2_ASAP7_75t_SL g5359 ( 
.A(n_3349),
.B(n_3371),
.Y(n_5359)
);

BUFx12f_ASAP7_75t_L g5360 ( 
.A(n_4350),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_4691),
.Y(n_5361)
);

OAI22xp5_ASAP7_75t_L g5362 ( 
.A1(n_3524),
.A2(n_3533),
.B1(n_3537),
.B2(n_3530),
.Y(n_5362)
);

INVx1_ASAP7_75t_L g5363 ( 
.A(n_4245),
.Y(n_5363)
);

AOI21xp5_ASAP7_75t_L g5364 ( 
.A1(n_4568),
.A2(n_3640),
.B(n_3750),
.Y(n_5364)
);

NOR2xp33_ASAP7_75t_L g5365 ( 
.A(n_3623),
.B(n_3874),
.Y(n_5365)
);

AOI21xp5_ASAP7_75t_L g5366 ( 
.A1(n_4568),
.A2(n_3625),
.B(n_3621),
.Y(n_5366)
);

AOI21xp5_ASAP7_75t_L g5367 ( 
.A1(n_4568),
.A2(n_3651),
.B(n_3663),
.Y(n_5367)
);

AOI21xp5_ASAP7_75t_L g5368 ( 
.A1(n_3651),
.A2(n_3663),
.B(n_4021),
.Y(n_5368)
);

NOR3xp33_ASAP7_75t_L g5369 ( 
.A(n_4099),
.B(n_3530),
.C(n_3524),
.Y(n_5369)
);

INVx1_ASAP7_75t_L g5370 ( 
.A(n_4268),
.Y(n_5370)
);

NAND2xp5_ASAP7_75t_L g5371 ( 
.A(n_3533),
.B(n_3537),
.Y(n_5371)
);

BUFx2_ASAP7_75t_L g5372 ( 
.A(n_3272),
.Y(n_5372)
);

BUFx5_ASAP7_75t_L g5373 ( 
.A(n_4507),
.Y(n_5373)
);

OAI21xp5_ASAP7_75t_L g5374 ( 
.A1(n_3853),
.A2(n_3557),
.B(n_3580),
.Y(n_5374)
);

NAND2xp5_ASAP7_75t_L g5375 ( 
.A(n_3538),
.B(n_3540),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_3538),
.B(n_3540),
.Y(n_5376)
);

AOI21xp5_ASAP7_75t_L g5377 ( 
.A1(n_4021),
.A2(n_4471),
.B(n_4412),
.Y(n_5377)
);

OAI22xp5_ASAP7_75t_L g5378 ( 
.A1(n_3542),
.A2(n_3559),
.B1(n_3571),
.B2(n_3545),
.Y(n_5378)
);

AOI21xp5_ASAP7_75t_L g5379 ( 
.A1(n_4471),
.A2(n_4660),
.B(n_4585),
.Y(n_5379)
);

NOR2xp33_ASAP7_75t_L g5380 ( 
.A(n_3623),
.B(n_3874),
.Y(n_5380)
);

NAND2xp5_ASAP7_75t_L g5381 ( 
.A(n_3542),
.B(n_3545),
.Y(n_5381)
);

INVx3_ASAP7_75t_L g5382 ( 
.A(n_3349),
.Y(n_5382)
);

AOI21xp5_ASAP7_75t_L g5383 ( 
.A1(n_4585),
.A2(n_4660),
.B(n_3267),
.Y(n_5383)
);

BUFx2_ASAP7_75t_L g5384 ( 
.A(n_3272),
.Y(n_5384)
);

NAND2xp5_ASAP7_75t_L g5385 ( 
.A(n_3559),
.B(n_3571),
.Y(n_5385)
);

NOR2xp33_ASAP7_75t_L g5386 ( 
.A(n_3337),
.B(n_4201),
.Y(n_5386)
);

OAI22xp5_ASAP7_75t_L g5387 ( 
.A1(n_3574),
.A2(n_3592),
.B1(n_3607),
.B2(n_3577),
.Y(n_5387)
);

NOR2xp33_ASAP7_75t_L g5388 ( 
.A(n_3337),
.B(n_4201),
.Y(n_5388)
);

OAI22xp5_ASAP7_75t_SL g5389 ( 
.A1(n_4099),
.A2(n_3960),
.B1(n_4671),
.B2(n_4386),
.Y(n_5389)
);

INVx2_ASAP7_75t_L g5390 ( 
.A(n_3521),
.Y(n_5390)
);

OAI22xp5_ASAP7_75t_L g5391 ( 
.A1(n_3574),
.A2(n_3592),
.B1(n_3607),
.B2(n_3577),
.Y(n_5391)
);

A2O1A1Ixp33_ASAP7_75t_L g5392 ( 
.A1(n_4028),
.A2(n_4064),
.B(n_4070),
.C(n_3786),
.Y(n_5392)
);

O2A1O1Ixp33_ASAP7_75t_L g5393 ( 
.A1(n_3609),
.A2(n_3628),
.B(n_3631),
.C(n_3629),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_L g5394 ( 
.A(n_3609),
.B(n_3628),
.Y(n_5394)
);

NAND2xp5_ASAP7_75t_L g5395 ( 
.A(n_3629),
.B(n_3631),
.Y(n_5395)
);

AOI21xp5_ASAP7_75t_L g5396 ( 
.A1(n_4585),
.A2(n_4660),
.B(n_3267),
.Y(n_5396)
);

AOI21xp5_ASAP7_75t_L g5397 ( 
.A1(n_3260),
.A2(n_3267),
.B(n_3557),
.Y(n_5397)
);

A2O1A1Ixp33_ASAP7_75t_L g5398 ( 
.A1(n_4070),
.A2(n_3786),
.B(n_4065),
.C(n_3997),
.Y(n_5398)
);

AND2x2_ASAP7_75t_L g5399 ( 
.A(n_3755),
.B(n_3572),
.Y(n_5399)
);

NAND2xp5_ASAP7_75t_SL g5400 ( 
.A(n_3643),
.B(n_3659),
.Y(n_5400)
);

AOI21xp5_ASAP7_75t_L g5401 ( 
.A1(n_3260),
.A2(n_3940),
.B(n_3896),
.Y(n_5401)
);

AOI22x1_ASAP7_75t_L g5402 ( 
.A1(n_4466),
.A2(n_3995),
.B1(n_3390),
.B2(n_4022),
.Y(n_5402)
);

NOR2xp33_ASAP7_75t_L g5403 ( 
.A(n_4502),
.B(n_4582),
.Y(n_5403)
);

OR2x2_ASAP7_75t_L g5404 ( 
.A(n_3434),
.B(n_3497),
.Y(n_5404)
);

AND2x2_ASAP7_75t_L g5405 ( 
.A(n_3755),
.B(n_3572),
.Y(n_5405)
);

AOI22xp33_ASAP7_75t_L g5406 ( 
.A1(n_3692),
.A2(n_3398),
.B1(n_3546),
.B2(n_3541),
.Y(n_5406)
);

AOI21xp5_ASAP7_75t_L g5407 ( 
.A1(n_3940),
.A2(n_3708),
.B(n_3912),
.Y(n_5407)
);

NAND2xp5_ASAP7_75t_L g5408 ( 
.A(n_3643),
.B(n_3659),
.Y(n_5408)
);

BUFx2_ASAP7_75t_L g5409 ( 
.A(n_3521),
.Y(n_5409)
);

AOI21xp5_ASAP7_75t_L g5410 ( 
.A1(n_3708),
.A2(n_3921),
.B(n_3912),
.Y(n_5410)
);

AOI21xp5_ASAP7_75t_L g5411 ( 
.A1(n_3921),
.A2(n_3939),
.B(n_3926),
.Y(n_5411)
);

NAND2xp5_ASAP7_75t_SL g5412 ( 
.A(n_3661),
.B(n_3665),
.Y(n_5412)
);

NAND2xp5_ASAP7_75t_L g5413 ( 
.A(n_3661),
.B(n_3665),
.Y(n_5413)
);

NAND3xp33_ASAP7_75t_L g5414 ( 
.A(n_3465),
.B(n_3614),
.C(n_3580),
.Y(n_5414)
);

AOI21xp5_ASAP7_75t_L g5415 ( 
.A1(n_3926),
.A2(n_3944),
.B(n_3939),
.Y(n_5415)
);

AOI21xp5_ASAP7_75t_L g5416 ( 
.A1(n_3944),
.A2(n_3955),
.B(n_3954),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_3521),
.Y(n_5417)
);

AOI21xp5_ASAP7_75t_L g5418 ( 
.A1(n_3954),
.A2(n_3958),
.B(n_3955),
.Y(n_5418)
);

INVx2_ASAP7_75t_L g5419 ( 
.A(n_3521),
.Y(n_5419)
);

OAI22xp5_ASAP7_75t_L g5420 ( 
.A1(n_3668),
.A2(n_3681),
.B1(n_3687),
.B2(n_3678),
.Y(n_5420)
);

CKINVDCx10_ASAP7_75t_R g5421 ( 
.A(n_3904),
.Y(n_5421)
);

OAI22xp5_ASAP7_75t_L g5422 ( 
.A1(n_3668),
.A2(n_3681),
.B1(n_3687),
.B2(n_3678),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_3420),
.B(n_3958),
.Y(n_5423)
);

AOI21xp5_ASAP7_75t_L g5424 ( 
.A1(n_3963),
.A2(n_3975),
.B(n_3966),
.Y(n_5424)
);

NOR2xp33_ASAP7_75t_L g5425 ( 
.A(n_4502),
.B(n_4582),
.Y(n_5425)
);

AOI21xp5_ASAP7_75t_L g5426 ( 
.A1(n_3963),
.A2(n_3975),
.B(n_3966),
.Y(n_5426)
);

OAI22xp5_ASAP7_75t_L g5427 ( 
.A1(n_3863),
.A2(n_4059),
.B1(n_4671),
.B2(n_4386),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_L g5428 ( 
.A(n_3420),
.B(n_3978),
.Y(n_5428)
);

AOI22xp5_ASAP7_75t_L g5429 ( 
.A1(n_3692),
.A2(n_4066),
.B1(n_3825),
.B2(n_3840),
.Y(n_5429)
);

AOI21x1_ASAP7_75t_L g5430 ( 
.A1(n_4285),
.A2(n_4298),
.B(n_4287),
.Y(n_5430)
);

AOI21xp5_ASAP7_75t_L g5431 ( 
.A1(n_3978),
.A2(n_3984),
.B(n_3980),
.Y(n_5431)
);

INVx3_ASAP7_75t_L g5432 ( 
.A(n_3349),
.Y(n_5432)
);

OAI21xp33_ASAP7_75t_SL g5433 ( 
.A1(n_3979),
.A2(n_3764),
.B(n_3390),
.Y(n_5433)
);

NAND2xp5_ASAP7_75t_L g5434 ( 
.A(n_3980),
.B(n_3984),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_4287),
.Y(n_5435)
);

AOI21xp5_ASAP7_75t_L g5436 ( 
.A1(n_3987),
.A2(n_3998),
.B(n_3989),
.Y(n_5436)
);

NAND2xp5_ASAP7_75t_L g5437 ( 
.A(n_3987),
.B(n_3989),
.Y(n_5437)
);

XOR2xp5_ASAP7_75t_L g5438 ( 
.A(n_3644),
.B(n_3960),
.Y(n_5438)
);

INVx5_ASAP7_75t_L g5439 ( 
.A(n_3219),
.Y(n_5439)
);

BUFx2_ASAP7_75t_L g5440 ( 
.A(n_3521),
.Y(n_5440)
);

AOI221xp5_ASAP7_75t_L g5441 ( 
.A1(n_4034),
.A2(n_3683),
.B1(n_3686),
.B2(n_3660),
.C(n_3614),
.Y(n_5441)
);

NAND2xp5_ASAP7_75t_L g5442 ( 
.A(n_3998),
.B(n_4004),
.Y(n_5442)
);

AND2x2_ASAP7_75t_L g5443 ( 
.A(n_3755),
.B(n_3572),
.Y(n_5443)
);

AOI21xp5_ASAP7_75t_L g5444 ( 
.A1(n_4004),
.A2(n_4018),
.B(n_3816),
.Y(n_5444)
);

NAND2xp5_ASAP7_75t_L g5445 ( 
.A(n_4018),
.B(n_3660),
.Y(n_5445)
);

NAND2xp5_ASAP7_75t_SL g5446 ( 
.A(n_4035),
.B(n_3697),
.Y(n_5446)
);

OAI21xp33_ASAP7_75t_L g5447 ( 
.A1(n_4034),
.A2(n_3863),
.B(n_3697),
.Y(n_5447)
);

NAND2xp5_ASAP7_75t_SL g5448 ( 
.A(n_4035),
.B(n_3732),
.Y(n_5448)
);

AOI22xp5_ASAP7_75t_L g5449 ( 
.A1(n_3692),
.A2(n_4066),
.B1(n_3825),
.B2(n_3997),
.Y(n_5449)
);

NAND2xp5_ASAP7_75t_L g5450 ( 
.A(n_3683),
.B(n_3686),
.Y(n_5450)
);

BUFx6f_ASAP7_75t_L g5451 ( 
.A(n_3349),
.Y(n_5451)
);

AOI21xp5_ASAP7_75t_L g5452 ( 
.A1(n_3816),
.A2(n_4283),
.B(n_3219),
.Y(n_5452)
);

INVx2_ASAP7_75t_SL g5453 ( 
.A(n_3539),
.Y(n_5453)
);

AND2x6_ASAP7_75t_L g5454 ( 
.A(n_3254),
.B(n_3274),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_4685),
.Y(n_5455)
);

AOI21xp5_ASAP7_75t_L g5456 ( 
.A1(n_3219),
.A2(n_4284),
.B(n_4283),
.Y(n_5456)
);

NOR2xp33_ASAP7_75t_L g5457 ( 
.A(n_4592),
.B(n_3922),
.Y(n_5457)
);

NOR2xp33_ASAP7_75t_L g5458 ( 
.A(n_4592),
.B(n_3922),
.Y(n_5458)
);

AOI21xp5_ASAP7_75t_L g5459 ( 
.A1(n_3219),
.A2(n_4284),
.B(n_4283),
.Y(n_5459)
);

BUFx2_ASAP7_75t_L g5460 ( 
.A(n_3531),
.Y(n_5460)
);

NAND2xp5_ASAP7_75t_L g5461 ( 
.A(n_3719),
.B(n_3748),
.Y(n_5461)
);

NAND2xp5_ASAP7_75t_L g5462 ( 
.A(n_3719),
.B(n_3748),
.Y(n_5462)
);

INVx8_ASAP7_75t_L g5463 ( 
.A(n_4526),
.Y(n_5463)
);

A2O1A1Ixp33_ASAP7_75t_L g5464 ( 
.A1(n_4065),
.A2(n_3892),
.B(n_4081),
.C(n_3390),
.Y(n_5464)
);

NAND2xp5_ASAP7_75t_L g5465 ( 
.A(n_4702),
.B(n_3434),
.Y(n_5465)
);

AOI22xp5_ASAP7_75t_L g5466 ( 
.A1(n_3692),
.A2(n_3782),
.B1(n_3856),
.B2(n_3791),
.Y(n_5466)
);

NAND2xp5_ASAP7_75t_L g5467 ( 
.A(n_4702),
.B(n_3434),
.Y(n_5467)
);

AOI22xp33_ASAP7_75t_L g5468 ( 
.A1(n_3398),
.A2(n_3541),
.B1(n_3546),
.B2(n_3499),
.Y(n_5468)
);

A2O1A1Ixp33_ASAP7_75t_L g5469 ( 
.A1(n_4065),
.A2(n_3892),
.B(n_4081),
.C(n_3390),
.Y(n_5469)
);

AND2x2_ASAP7_75t_L g5470 ( 
.A(n_3572),
.B(n_3613),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_4298),
.Y(n_5471)
);

NAND2xp5_ASAP7_75t_L g5472 ( 
.A(n_3497),
.B(n_3570),
.Y(n_5472)
);

NAND2xp5_ASAP7_75t_L g5473 ( 
.A(n_3497),
.B(n_3570),
.Y(n_5473)
);

NAND2xp5_ASAP7_75t_L g5474 ( 
.A(n_3570),
.B(n_3717),
.Y(n_5474)
);

O2A1O1Ixp33_ASAP7_75t_L g5475 ( 
.A1(n_3869),
.A2(n_3898),
.B(n_3905),
.C(n_3894),
.Y(n_5475)
);

AOI21xp5_ASAP7_75t_L g5476 ( 
.A1(n_3219),
.A2(n_4284),
.B(n_4283),
.Y(n_5476)
);

AOI21xp5_ASAP7_75t_L g5477 ( 
.A1(n_3219),
.A2(n_4284),
.B(n_4283),
.Y(n_5477)
);

OR2x6_ASAP7_75t_SL g5478 ( 
.A(n_3717),
.B(n_4169),
.Y(n_5478)
);

AOI22x1_ASAP7_75t_L g5479 ( 
.A1(n_3995),
.A2(n_4023),
.B1(n_4032),
.B2(n_4022),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_4685),
.Y(n_5480)
);

AOI21xp5_ASAP7_75t_L g5481 ( 
.A1(n_3219),
.A2(n_4284),
.B(n_4283),
.Y(n_5481)
);

AOI21x1_ASAP7_75t_L g5482 ( 
.A1(n_4299),
.A2(n_4322),
.B(n_4315),
.Y(n_5482)
);

AND2x2_ASAP7_75t_L g5483 ( 
.A(n_3572),
.B(n_3613),
.Y(n_5483)
);

AOI21xp5_ASAP7_75t_L g5484 ( 
.A1(n_3219),
.A2(n_4284),
.B(n_4283),
.Y(n_5484)
);

NOR2xp33_ASAP7_75t_L g5485 ( 
.A(n_3798),
.B(n_3820),
.Y(n_5485)
);

NOR2xp33_ASAP7_75t_L g5486 ( 
.A(n_3798),
.B(n_3820),
.Y(n_5486)
);

O2A1O1Ixp33_ASAP7_75t_L g5487 ( 
.A1(n_3869),
.A2(n_3898),
.B(n_3905),
.C(n_3894),
.Y(n_5487)
);

O2A1O1Ixp33_ASAP7_75t_SL g5488 ( 
.A1(n_4116),
.A2(n_4126),
.B(n_4119),
.C(n_4121),
.Y(n_5488)
);

INVx2_ASAP7_75t_L g5489 ( 
.A(n_3531),
.Y(n_5489)
);

A2O1A1Ixp33_ASAP7_75t_L g5490 ( 
.A1(n_4065),
.A2(n_4095),
.B(n_4031),
.C(n_3546),
.Y(n_5490)
);

AOI21xp5_ASAP7_75t_L g5491 ( 
.A1(n_4283),
.A2(n_4311),
.B(n_4284),
.Y(n_5491)
);

A2O1A1Ixp33_ASAP7_75t_L g5492 ( 
.A1(n_4065),
.A2(n_4095),
.B(n_4031),
.C(n_3764),
.Y(n_5492)
);

NOR2xp33_ASAP7_75t_L g5493 ( 
.A(n_3677),
.B(n_3461),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_3531),
.Y(n_5494)
);

INVx2_ASAP7_75t_L g5495 ( 
.A(n_3531),
.Y(n_5495)
);

INVx2_ASAP7_75t_L g5496 ( 
.A(n_3531),
.Y(n_5496)
);

NAND2xp5_ASAP7_75t_L g5497 ( 
.A(n_3717),
.B(n_4702),
.Y(n_5497)
);

OA22x2_ASAP7_75t_L g5498 ( 
.A1(n_3499),
.A2(n_3732),
.B1(n_3774),
.B2(n_3738),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_3531),
.Y(n_5499)
);

OAI22xp5_ASAP7_75t_L g5500 ( 
.A1(n_4386),
.A2(n_4671),
.B1(n_3461),
.B2(n_4646),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_4688),
.Y(n_5501)
);

OAI22xp5_ASAP7_75t_L g5502 ( 
.A1(n_3792),
.A2(n_4646),
.B1(n_3242),
.B2(n_3774),
.Y(n_5502)
);

NAND2xp5_ASAP7_75t_L g5503 ( 
.A(n_4169),
.B(n_4180),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_4169),
.B(n_4180),
.Y(n_5504)
);

INVx2_ASAP7_75t_L g5505 ( 
.A(n_3531),
.Y(n_5505)
);

NAND2xp5_ASAP7_75t_L g5506 ( 
.A(n_4180),
.B(n_4428),
.Y(n_5506)
);

NAND2xp5_ASAP7_75t_L g5507 ( 
.A(n_4428),
.B(n_4436),
.Y(n_5507)
);

AOI21x1_ASAP7_75t_L g5508 ( 
.A1(n_4299),
.A2(n_4322),
.B(n_4315),
.Y(n_5508)
);

NAND2xp5_ASAP7_75t_L g5509 ( 
.A(n_4428),
.B(n_4436),
.Y(n_5509)
);

AND2x2_ASAP7_75t_L g5510 ( 
.A(n_3572),
.B(n_3613),
.Y(n_5510)
);

INVx2_ASAP7_75t_L g5511 ( 
.A(n_3531),
.Y(n_5511)
);

AOI21xp5_ASAP7_75t_L g5512 ( 
.A1(n_4284),
.A2(n_4342),
.B(n_4311),
.Y(n_5512)
);

AND2x4_ASAP7_75t_L g5513 ( 
.A(n_3301),
.B(n_3381),
.Y(n_5513)
);

BUFx8_ASAP7_75t_L g5514 ( 
.A(n_3415),
.Y(n_5514)
);

O2A1O1Ixp33_ASAP7_75t_SL g5515 ( 
.A1(n_4116),
.A2(n_4119),
.B(n_4126),
.C(n_4088),
.Y(n_5515)
);

NOR2xp33_ASAP7_75t_L g5516 ( 
.A(n_3677),
.B(n_3792),
.Y(n_5516)
);

OAI22xp5_ASAP7_75t_L g5517 ( 
.A1(n_3242),
.A2(n_3818),
.B1(n_3738),
.B2(n_4005),
.Y(n_5517)
);

OAI22xp5_ASAP7_75t_L g5518 ( 
.A1(n_3818),
.A2(n_4005),
.B1(n_3977),
.B2(n_3913),
.Y(n_5518)
);

OAI21x1_ASAP7_75t_L g5519 ( 
.A1(n_4294),
.A2(n_4341),
.B(n_4340),
.Y(n_5519)
);

AND2x2_ASAP7_75t_L g5520 ( 
.A(n_3572),
.B(n_3613),
.Y(n_5520)
);

AOI21xp5_ASAP7_75t_L g5521 ( 
.A1(n_4311),
.A2(n_4356),
.B(n_4342),
.Y(n_5521)
);

NAND2xp5_ASAP7_75t_L g5522 ( 
.A(n_4436),
.B(n_4495),
.Y(n_5522)
);

AOI22xp5_ASAP7_75t_L g5523 ( 
.A1(n_3856),
.A2(n_4088),
.B1(n_3979),
.B2(n_3499),
.Y(n_5523)
);

BUFx6f_ASAP7_75t_L g5524 ( 
.A(n_3349),
.Y(n_5524)
);

OR2x6_ASAP7_75t_SL g5525 ( 
.A(n_4495),
.B(n_4569),
.Y(n_5525)
);

BUFx6f_ASAP7_75t_L g5526 ( 
.A(n_3371),
.Y(n_5526)
);

NAND2xp5_ASAP7_75t_SL g5527 ( 
.A(n_3637),
.B(n_3429),
.Y(n_5527)
);

NAND3xp33_ASAP7_75t_L g5528 ( 
.A(n_3893),
.B(n_4006),
.C(n_3913),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_4687),
.Y(n_5529)
);

OAI22xp5_ASAP7_75t_L g5530 ( 
.A1(n_3977),
.A2(n_4006),
.B1(n_3893),
.B2(n_3838),
.Y(n_5530)
);

NOR3xp33_ASAP7_75t_L g5531 ( 
.A(n_4092),
.B(n_4122),
.C(n_4109),
.Y(n_5531)
);

OAI21xp5_ASAP7_75t_L g5532 ( 
.A1(n_3303),
.A2(n_3718),
.B(n_3441),
.Y(n_5532)
);

NAND2xp33_ASAP7_75t_L g5533 ( 
.A(n_4583),
.B(n_3819),
.Y(n_5533)
);

NAND2xp5_ASAP7_75t_L g5534 ( 
.A(n_4495),
.B(n_4569),
.Y(n_5534)
);

AOI21xp5_ASAP7_75t_L g5535 ( 
.A1(n_4311),
.A2(n_4356),
.B(n_4342),
.Y(n_5535)
);

O2A1O1Ixp33_ASAP7_75t_SL g5536 ( 
.A1(n_4109),
.A2(n_4092),
.B(n_4079),
.C(n_4129),
.Y(n_5536)
);

OAI22xp5_ASAP7_75t_L g5537 ( 
.A1(n_3977),
.A2(n_4297),
.B1(n_4374),
.B2(n_4175),
.Y(n_5537)
);

NOR2xp33_ASAP7_75t_SL g5538 ( 
.A(n_4526),
.B(n_3789),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_4324),
.Y(n_5539)
);

OAI21xp5_ASAP7_75t_L g5540 ( 
.A1(n_3303),
.A2(n_3718),
.B(n_3441),
.Y(n_5540)
);

OAI22xp5_ASAP7_75t_L g5541 ( 
.A1(n_4297),
.A2(n_4420),
.B1(n_4561),
.B2(n_4374),
.Y(n_5541)
);

INVxp67_ASAP7_75t_L g5542 ( 
.A(n_3839),
.Y(n_5542)
);

NAND2xp5_ASAP7_75t_L g5543 ( 
.A(n_4569),
.B(n_4680),
.Y(n_5543)
);

AO22x1_ASAP7_75t_L g5544 ( 
.A1(n_4047),
.A2(n_3539),
.B1(n_3637),
.B2(n_3626),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_L g5545 ( 
.A(n_4599),
.B(n_4680),
.Y(n_5545)
);

NAND2xp5_ASAP7_75t_SL g5546 ( 
.A(n_3637),
.B(n_3429),
.Y(n_5546)
);

AOI21x1_ASAP7_75t_L g5547 ( 
.A1(n_4346),
.A2(n_4358),
.B(n_4352),
.Y(n_5547)
);

AOI21xp5_ASAP7_75t_L g5548 ( 
.A1(n_4311),
.A2(n_4356),
.B(n_4342),
.Y(n_5548)
);

OAI22xp5_ASAP7_75t_L g5549 ( 
.A1(n_4420),
.A2(n_4613),
.B1(n_4638),
.B2(n_4561),
.Y(n_5549)
);

OAI22xp5_ASAP7_75t_L g5550 ( 
.A1(n_4613),
.A2(n_4638),
.B1(n_4060),
.B2(n_4038),
.Y(n_5550)
);

AO22x1_ASAP7_75t_L g5551 ( 
.A1(n_4047),
.A2(n_3637),
.B1(n_3707),
.B2(n_3626),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_4363),
.Y(n_5552)
);

INVx2_ASAP7_75t_L g5553 ( 
.A(n_3581),
.Y(n_5553)
);

AOI21xp5_ASAP7_75t_L g5554 ( 
.A1(n_4311),
.A2(n_4356),
.B(n_4342),
.Y(n_5554)
);

AND2x2_ASAP7_75t_L g5555 ( 
.A(n_3613),
.B(n_3581),
.Y(n_5555)
);

NAND2xp5_ASAP7_75t_L g5556 ( 
.A(n_4599),
.B(n_4680),
.Y(n_5556)
);

OAI22xp5_ASAP7_75t_L g5557 ( 
.A1(n_4060),
.A2(n_4038),
.B1(n_4093),
.B2(n_4089),
.Y(n_5557)
);

OA22x2_ASAP7_75t_L g5558 ( 
.A1(n_3398),
.A2(n_3429),
.B1(n_3367),
.B2(n_4098),
.Y(n_5558)
);

BUFx6f_ASAP7_75t_L g5559 ( 
.A(n_3371),
.Y(n_5559)
);

AOI21x1_ASAP7_75t_L g5560 ( 
.A1(n_4365),
.A2(n_4390),
.B(n_4368),
.Y(n_5560)
);

AOI21xp5_ASAP7_75t_L g5561 ( 
.A1(n_4311),
.A2(n_4356),
.B(n_4342),
.Y(n_5561)
);

NOR2xp33_ASAP7_75t_L g5562 ( 
.A(n_3787),
.B(n_3907),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_4391),
.Y(n_5563)
);

CKINVDCx10_ASAP7_75t_R g5564 ( 
.A(n_3904),
.Y(n_5564)
);

NAND2xp5_ASAP7_75t_L g5565 ( 
.A(n_4599),
.B(n_3290),
.Y(n_5565)
);

INVx2_ASAP7_75t_L g5566 ( 
.A(n_3581),
.Y(n_5566)
);

NOR2xp33_ASAP7_75t_SL g5567 ( 
.A(n_3789),
.B(n_3385),
.Y(n_5567)
);

AOI21xp5_ASAP7_75t_L g5568 ( 
.A1(n_4311),
.A2(n_4356),
.B(n_4342),
.Y(n_5568)
);

AOI21x1_ASAP7_75t_L g5569 ( 
.A1(n_4391),
.A2(n_4403),
.B(n_4398),
.Y(n_5569)
);

BUFx6f_ASAP7_75t_L g5570 ( 
.A(n_3371),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_SL g5571 ( 
.A(n_3637),
.B(n_3429),
.Y(n_5571)
);

NAND2xp5_ASAP7_75t_L g5572 ( 
.A(n_3290),
.B(n_3296),
.Y(n_5572)
);

OR2x6_ASAP7_75t_SL g5573 ( 
.A(n_3268),
.B(n_3290),
.Y(n_5573)
);

AOI21xp5_ASAP7_75t_L g5574 ( 
.A1(n_4342),
.A2(n_4389),
.B(n_4356),
.Y(n_5574)
);

NAND2xp5_ASAP7_75t_L g5575 ( 
.A(n_3296),
.B(n_3323),
.Y(n_5575)
);

BUFx4f_ASAP7_75t_L g5576 ( 
.A(n_3448),
.Y(n_5576)
);

AOI21xp5_ASAP7_75t_L g5577 ( 
.A1(n_4356),
.A2(n_4413),
.B(n_4389),
.Y(n_5577)
);

OAI21xp33_ASAP7_75t_L g5578 ( 
.A1(n_4056),
.A2(n_3908),
.B(n_3902),
.Y(n_5578)
);

NAND2xp5_ASAP7_75t_L g5579 ( 
.A(n_3296),
.B(n_3323),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_4398),
.Y(n_5580)
);

AND2x4_ASAP7_75t_L g5581 ( 
.A(n_3345),
.B(n_3351),
.Y(n_5581)
);

NAND2xp5_ASAP7_75t_L g5582 ( 
.A(n_3323),
.B(n_3328),
.Y(n_5582)
);

A2O1A1Ixp33_ASAP7_75t_L g5583 ( 
.A1(n_3605),
.A2(n_4063),
.B(n_3979),
.C(n_4113),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_3328),
.B(n_3333),
.Y(n_5584)
);

NAND2xp5_ASAP7_75t_L g5585 ( 
.A(n_3328),
.B(n_3333),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_4403),
.Y(n_5586)
);

O2A1O1Ixp33_ASAP7_75t_L g5587 ( 
.A1(n_3906),
.A2(n_3914),
.B(n_3924),
.C(n_3917),
.Y(n_5587)
);

INVx2_ASAP7_75t_L g5588 ( 
.A(n_3581),
.Y(n_5588)
);

INVxp67_ASAP7_75t_L g5589 ( 
.A(n_3839),
.Y(n_5589)
);

AOI21xp5_ASAP7_75t_L g5590 ( 
.A1(n_4389),
.A2(n_4473),
.B(n_4413),
.Y(n_5590)
);

O2A1O1Ixp33_ASAP7_75t_L g5591 ( 
.A1(n_3906),
.A2(n_3914),
.B(n_3924),
.C(n_3917),
.Y(n_5591)
);

OAI21xp5_ASAP7_75t_L g5592 ( 
.A1(n_3303),
.A2(n_3718),
.B(n_3441),
.Y(n_5592)
);

NAND2xp5_ASAP7_75t_L g5593 ( 
.A(n_3333),
.B(n_3363),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_4404),
.Y(n_5594)
);

AOI22xp5_ASAP7_75t_L g5595 ( 
.A1(n_3979),
.A2(n_3936),
.B1(n_3967),
.B2(n_4122),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_4404),
.Y(n_5596)
);

BUFx6f_ASAP7_75t_L g5597 ( 
.A(n_3371),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_4414),
.Y(n_5598)
);

NAND2xp5_ASAP7_75t_L g5599 ( 
.A(n_3363),
.B(n_3369),
.Y(n_5599)
);

BUFx2_ASAP7_75t_L g5600 ( 
.A(n_3581),
.Y(n_5600)
);

OAI21xp33_ASAP7_75t_L g5601 ( 
.A1(n_4056),
.A2(n_3908),
.B(n_3902),
.Y(n_5601)
);

INVx2_ASAP7_75t_L g5602 ( 
.A(n_3583),
.Y(n_5602)
);

OAI21x1_ASAP7_75t_L g5603 ( 
.A1(n_4294),
.A2(n_4341),
.B(n_4340),
.Y(n_5603)
);

NAND2xp5_ASAP7_75t_L g5604 ( 
.A(n_3363),
.B(n_3369),
.Y(n_5604)
);

NAND2xp5_ASAP7_75t_L g5605 ( 
.A(n_3369),
.B(n_3386),
.Y(n_5605)
);

BUFx6f_ASAP7_75t_L g5606 ( 
.A(n_3371),
.Y(n_5606)
);

NAND3xp33_ASAP7_75t_SL g5607 ( 
.A(n_3819),
.B(n_4463),
.C(n_4093),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_4414),
.Y(n_5608)
);

NAND2xp5_ASAP7_75t_L g5609 ( 
.A(n_3386),
.B(n_3389),
.Y(n_5609)
);

NOR2xp33_ASAP7_75t_L g5610 ( 
.A(n_3787),
.B(n_3907),
.Y(n_5610)
);

AOI21xp5_ASAP7_75t_L g5611 ( 
.A1(n_4389),
.A2(n_4473),
.B(n_4413),
.Y(n_5611)
);

INVx1_ASAP7_75t_L g5612 ( 
.A(n_4416),
.Y(n_5612)
);

INVx3_ASAP7_75t_L g5613 ( 
.A(n_3371),
.Y(n_5613)
);

AOI21xp5_ASAP7_75t_L g5614 ( 
.A1(n_4389),
.A2(n_4473),
.B(n_4413),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_4416),
.Y(n_5615)
);

O2A1O1Ixp33_ASAP7_75t_L g5616 ( 
.A1(n_3936),
.A2(n_3967),
.B(n_4061),
.C(n_4113),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_4425),
.Y(n_5617)
);

OAI21xp5_ASAP7_75t_L g5618 ( 
.A1(n_3303),
.A2(n_3718),
.B(n_3441),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_4425),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_L g5620 ( 
.A(n_3386),
.B(n_3389),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_L g5621 ( 
.A(n_3389),
.B(n_3396),
.Y(n_5621)
);

INVx2_ASAP7_75t_L g5622 ( 
.A(n_3583),
.Y(n_5622)
);

NAND2xp5_ASAP7_75t_L g5623 ( 
.A(n_3396),
.B(n_3397),
.Y(n_5623)
);

AOI21xp5_ASAP7_75t_L g5624 ( 
.A1(n_4389),
.A2(n_4473),
.B(n_4413),
.Y(n_5624)
);

HB1xp67_ASAP7_75t_L g5625 ( 
.A(n_4098),
.Y(n_5625)
);

INVx5_ASAP7_75t_L g5626 ( 
.A(n_4389),
.Y(n_5626)
);

AOI21xp5_ASAP7_75t_L g5627 ( 
.A1(n_4389),
.A2(n_4473),
.B(n_4413),
.Y(n_5627)
);

NOR3xp33_ASAP7_75t_L g5628 ( 
.A(n_4061),
.B(n_4076),
.C(n_4090),
.Y(n_5628)
);

NAND2xp5_ASAP7_75t_L g5629 ( 
.A(n_3396),
.B(n_3397),
.Y(n_5629)
);

AOI21xp5_ASAP7_75t_L g5630 ( 
.A1(n_4413),
.A2(n_4480),
.B(n_4473),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_4427),
.Y(n_5631)
);

AND2x2_ASAP7_75t_L g5632 ( 
.A(n_3613),
.B(n_3583),
.Y(n_5632)
);

A2O1A1Ixp33_ASAP7_75t_L g5633 ( 
.A1(n_3605),
.A2(n_4063),
.B(n_4113),
.C(n_3429),
.Y(n_5633)
);

OR2x2_ASAP7_75t_L g5634 ( 
.A(n_3613),
.B(n_3583),
.Y(n_5634)
);

NOR2x1p5_ASAP7_75t_SL g5635 ( 
.A(n_4643),
.B(n_4458),
.Y(n_5635)
);

A2O1A1Ixp33_ASAP7_75t_L g5636 ( 
.A1(n_3605),
.A2(n_4110),
.B(n_3548),
.C(n_3253),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_L g5637 ( 
.A(n_3397),
.B(n_3406),
.Y(n_5637)
);

NOR2xp33_ASAP7_75t_L g5638 ( 
.A(n_4072),
.B(n_4096),
.Y(n_5638)
);

BUFx2_ASAP7_75t_L g5639 ( 
.A(n_3583),
.Y(n_5639)
);

BUFx6f_ASAP7_75t_L g5640 ( 
.A(n_3371),
.Y(n_5640)
);

NAND2xp5_ASAP7_75t_SL g5641 ( 
.A(n_3637),
.B(n_3489),
.Y(n_5641)
);

AOI21xp5_ASAP7_75t_L g5642 ( 
.A1(n_4413),
.A2(n_4480),
.B(n_4473),
.Y(n_5642)
);

NOR2xp33_ASAP7_75t_L g5643 ( 
.A(n_4072),
.B(n_4096),
.Y(n_5643)
);

AOI21xp5_ASAP7_75t_L g5644 ( 
.A1(n_4473),
.A2(n_4493),
.B(n_4480),
.Y(n_5644)
);

O2A1O1Ixp33_ASAP7_75t_L g5645 ( 
.A1(n_4111),
.A2(n_4090),
.B(n_4107),
.C(n_3852),
.Y(n_5645)
);

OAI21xp5_ASAP7_75t_L g5646 ( 
.A1(n_3850),
.A2(n_4001),
.B(n_3988),
.Y(n_5646)
);

XOR2x2_ASAP7_75t_R g5647 ( 
.A(n_3364),
.B(n_3991),
.Y(n_5647)
);

A2O1A1Ixp33_ASAP7_75t_L g5648 ( 
.A1(n_3605),
.A2(n_4110),
.B(n_3548),
.C(n_3253),
.Y(n_5648)
);

INVx3_ASAP7_75t_L g5649 ( 
.A(n_3345),
.Y(n_5649)
);

AOI21xp5_ASAP7_75t_L g5650 ( 
.A1(n_4480),
.A2(n_4504),
.B(n_4493),
.Y(n_5650)
);

NOR2x1p5_ASAP7_75t_SL g5651 ( 
.A(n_4643),
.B(n_4462),
.Y(n_5651)
);

NOR2xp33_ASAP7_75t_L g5652 ( 
.A(n_4076),
.B(n_3925),
.Y(n_5652)
);

AOI21x1_ASAP7_75t_L g5653 ( 
.A1(n_4462),
.A2(n_4477),
.B(n_4468),
.Y(n_5653)
);

NAND2xp5_ASAP7_75t_SL g5654 ( 
.A(n_3637),
.B(n_3489),
.Y(n_5654)
);

OAI321xp33_ASAP7_75t_L g5655 ( 
.A1(n_3836),
.A2(n_3852),
.A3(n_4089),
.B1(n_4032),
.B2(n_4023),
.C(n_4001),
.Y(n_5655)
);

NAND2xp5_ASAP7_75t_L g5656 ( 
.A(n_3406),
.B(n_3426),
.Y(n_5656)
);

NAND2xp5_ASAP7_75t_L g5657 ( 
.A(n_3406),
.B(n_3426),
.Y(n_5657)
);

OAI21xp5_ASAP7_75t_L g5658 ( 
.A1(n_3850),
.A2(n_3988),
.B(n_3268),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_4468),
.Y(n_5659)
);

AOI21xp5_ASAP7_75t_L g5660 ( 
.A1(n_4480),
.A2(n_4504),
.B(n_4493),
.Y(n_5660)
);

INVx2_ASAP7_75t_L g5661 ( 
.A(n_3583),
.Y(n_5661)
);

AOI21xp5_ASAP7_75t_L g5662 ( 
.A1(n_4480),
.A2(n_4504),
.B(n_4493),
.Y(n_5662)
);

O2A1O1Ixp33_ASAP7_75t_L g5663 ( 
.A1(n_4111),
.A2(n_4107),
.B(n_3852),
.C(n_3836),
.Y(n_5663)
);

NAND2xp5_ASAP7_75t_SL g5664 ( 
.A(n_3489),
.B(n_3525),
.Y(n_5664)
);

NAND2xp5_ASAP7_75t_L g5665 ( 
.A(n_3426),
.B(n_3427),
.Y(n_5665)
);

NAND2xp5_ASAP7_75t_L g5666 ( 
.A(n_3427),
.B(n_3435),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_4477),
.Y(n_5667)
);

INVxp67_ASAP7_75t_SL g5668 ( 
.A(n_3427),
.Y(n_5668)
);

AOI21xp5_ASAP7_75t_L g5669 ( 
.A1(n_4480),
.A2(n_4504),
.B(n_4493),
.Y(n_5669)
);

AOI22xp33_ASAP7_75t_L g5670 ( 
.A1(n_3364),
.A2(n_4476),
.B1(n_4607),
.B2(n_3253),
.Y(n_5670)
);

AOI21xp5_ASAP7_75t_L g5671 ( 
.A1(n_4480),
.A2(n_4504),
.B(n_4493),
.Y(n_5671)
);

NAND2xp5_ASAP7_75t_SL g5672 ( 
.A(n_3489),
.B(n_3525),
.Y(n_5672)
);

INVx2_ASAP7_75t_L g5673 ( 
.A(n_3583),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_4479),
.Y(n_5674)
);

NOR3xp33_ASAP7_75t_L g5675 ( 
.A(n_4079),
.B(n_4130),
.C(n_4148),
.Y(n_5675)
);

O2A1O1Ixp33_ASAP7_75t_SL g5676 ( 
.A1(n_4129),
.A2(n_4133),
.B(n_4138),
.C(n_4131),
.Y(n_5676)
);

AND2x2_ASAP7_75t_L g5677 ( 
.A(n_3583),
.B(n_3641),
.Y(n_5677)
);

NAND2xp5_ASAP7_75t_L g5678 ( 
.A(n_3435),
.B(n_3464),
.Y(n_5678)
);

OR2x2_ASAP7_75t_L g5679 ( 
.A(n_3641),
.B(n_3647),
.Y(n_5679)
);

INVx2_ASAP7_75t_L g5680 ( 
.A(n_3641),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_L g5681 ( 
.A(n_3435),
.B(n_3464),
.Y(n_5681)
);

NOR2xp33_ASAP7_75t_R g5682 ( 
.A(n_3562),
.B(n_3597),
.Y(n_5682)
);

NAND2xp5_ASAP7_75t_L g5683 ( 
.A(n_3464),
.B(n_3468),
.Y(n_5683)
);

O2A1O1Ixp33_ASAP7_75t_L g5684 ( 
.A1(n_4111),
.A2(n_4107),
.B(n_3836),
.C(n_3956),
.Y(n_5684)
);

AOI21xp5_ASAP7_75t_L g5685 ( 
.A1(n_4493),
.A2(n_4520),
.B(n_4504),
.Y(n_5685)
);

OR2x6_ASAP7_75t_L g5686 ( 
.A(n_3367),
.B(n_3756),
.Y(n_5686)
);

NOR2xp67_ASAP7_75t_L g5687 ( 
.A(n_4479),
.B(n_4487),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_4487),
.Y(n_5688)
);

AOI21xp5_ASAP7_75t_L g5689 ( 
.A1(n_4493),
.A2(n_4520),
.B(n_4504),
.Y(n_5689)
);

NAND2xp5_ASAP7_75t_L g5690 ( 
.A(n_3468),
.B(n_3472),
.Y(n_5690)
);

NAND2xp5_ASAP7_75t_SL g5691 ( 
.A(n_3489),
.B(n_3525),
.Y(n_5691)
);

CKINVDCx5p33_ASAP7_75t_R g5692 ( 
.A(n_3321),
.Y(n_5692)
);

INVx2_ASAP7_75t_L g5693 ( 
.A(n_3641),
.Y(n_5693)
);

OAI22xp5_ASAP7_75t_L g5694 ( 
.A1(n_4463),
.A2(n_3667),
.B1(n_3714),
.B2(n_3579),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_L g5695 ( 
.A(n_3468),
.B(n_3472),
.Y(n_5695)
);

OAI21xp5_ASAP7_75t_L g5696 ( 
.A1(n_3472),
.A2(n_3479),
.B(n_3478),
.Y(n_5696)
);

OAI21xp5_ASAP7_75t_L g5697 ( 
.A1(n_3478),
.A2(n_3480),
.B(n_3479),
.Y(n_5697)
);

NOR2xp33_ASAP7_75t_L g5698 ( 
.A(n_3925),
.B(n_4068),
.Y(n_5698)
);

INVx1_ASAP7_75t_L g5699 ( 
.A(n_4496),
.Y(n_5699)
);

NAND2xp5_ASAP7_75t_SL g5700 ( 
.A(n_3525),
.B(n_4073),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_4496),
.Y(n_5701)
);

NAND2xp5_ASAP7_75t_L g5702 ( 
.A(n_3478),
.B(n_3479),
.Y(n_5702)
);

AOI21xp5_ASAP7_75t_L g5703 ( 
.A1(n_4504),
.A2(n_4543),
.B(n_4520),
.Y(n_5703)
);

O2A1O1Ixp33_ASAP7_75t_L g5704 ( 
.A1(n_3952),
.A2(n_3956),
.B(n_3961),
.C(n_3959),
.Y(n_5704)
);

INVx5_ASAP7_75t_L g5705 ( 
.A(n_4520),
.Y(n_5705)
);

A2O1A1Ixp33_ASAP7_75t_L g5706 ( 
.A1(n_4110),
.A2(n_3548),
.B(n_4476),
.C(n_3253),
.Y(n_5706)
);

OR2x2_ASAP7_75t_L g5707 ( 
.A(n_3641),
.B(n_3647),
.Y(n_5707)
);

AOI21xp5_ASAP7_75t_L g5708 ( 
.A1(n_4520),
.A2(n_4612),
.B(n_4543),
.Y(n_5708)
);

AOI21xp5_ASAP7_75t_L g5709 ( 
.A1(n_4520),
.A2(n_4612),
.B(n_4543),
.Y(n_5709)
);

NOR2xp33_ASAP7_75t_L g5710 ( 
.A(n_4068),
.B(n_4046),
.Y(n_5710)
);

AOI21x1_ASAP7_75t_L g5711 ( 
.A1(n_4500),
.A2(n_4524),
.B(n_4509),
.Y(n_5711)
);

NAND2xp5_ASAP7_75t_L g5712 ( 
.A(n_3480),
.B(n_3501),
.Y(n_5712)
);

A2O1A1Ixp33_ASAP7_75t_L g5713 ( 
.A1(n_4110),
.A2(n_4683),
.B(n_4634),
.C(n_4607),
.Y(n_5713)
);

NAND2xp5_ASAP7_75t_L g5714 ( 
.A(n_3480),
.B(n_3501),
.Y(n_5714)
);

INVx3_ASAP7_75t_L g5715 ( 
.A(n_3345),
.Y(n_5715)
);

AND2x2_ASAP7_75t_L g5716 ( 
.A(n_3641),
.B(n_3647),
.Y(n_5716)
);

OAI321xp33_ASAP7_75t_L g5717 ( 
.A1(n_3765),
.A2(n_3778),
.A3(n_3821),
.B1(n_3770),
.B2(n_3590),
.C(n_3512),
.Y(n_5717)
);

OAI21x1_ASAP7_75t_L g5718 ( 
.A1(n_4294),
.A2(n_4341),
.B(n_4340),
.Y(n_5718)
);

CKINVDCx5p33_ASAP7_75t_R g5719 ( 
.A(n_4252),
.Y(n_5719)
);

OAI22xp5_ASAP7_75t_L g5720 ( 
.A1(n_4463),
.A2(n_3667),
.B1(n_3714),
.B2(n_3579),
.Y(n_5720)
);

OAI22xp5_ASAP7_75t_L g5721 ( 
.A1(n_3579),
.A2(n_3714),
.B1(n_3777),
.B2(n_3667),
.Y(n_5721)
);

OR2x6_ASAP7_75t_SL g5722 ( 
.A(n_3501),
.B(n_3514),
.Y(n_5722)
);

NOR2xp33_ASAP7_75t_L g5723 ( 
.A(n_4046),
.B(n_4074),
.Y(n_5723)
);

AOI21xp5_ASAP7_75t_L g5724 ( 
.A1(n_4520),
.A2(n_4612),
.B(n_4543),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_4500),
.Y(n_5725)
);

INVx1_ASAP7_75t_L g5726 ( 
.A(n_4509),
.Y(n_5726)
);

NAND2xp5_ASAP7_75t_SL g5727 ( 
.A(n_3525),
.B(n_4073),
.Y(n_5727)
);

AOI22xp33_ASAP7_75t_L g5728 ( 
.A1(n_3364),
.A2(n_4607),
.B1(n_4621),
.B2(n_4476),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_4524),
.Y(n_5729)
);

NAND2xp5_ASAP7_75t_L g5730 ( 
.A(n_3514),
.B(n_3519),
.Y(n_5730)
);

AOI22xp5_ASAP7_75t_L g5731 ( 
.A1(n_4046),
.A2(n_4130),
.B1(n_3957),
.B2(n_3920),
.Y(n_5731)
);

INVx2_ASAP7_75t_L g5732 ( 
.A(n_3641),
.Y(n_5732)
);

NAND3xp33_ASAP7_75t_L g5733 ( 
.A(n_4085),
.B(n_3959),
.C(n_3952),
.Y(n_5733)
);

NOR2xp33_ASAP7_75t_L g5734 ( 
.A(n_4074),
.B(n_3931),
.Y(n_5734)
);

NOR2x1p5_ASAP7_75t_SL g5735 ( 
.A(n_4643),
.B(n_4530),
.Y(n_5735)
);

AOI21xp5_ASAP7_75t_L g5736 ( 
.A1(n_4520),
.A2(n_4612),
.B(n_4543),
.Y(n_5736)
);

NOR2xp33_ASAP7_75t_L g5737 ( 
.A(n_4074),
.B(n_3931),
.Y(n_5737)
);

AOI22xp5_ASAP7_75t_L g5738 ( 
.A1(n_3957),
.A2(n_3920),
.B1(n_3904),
.B2(n_4147),
.Y(n_5738)
);

OR2x2_ASAP7_75t_L g5739 ( 
.A(n_3641),
.B(n_3647),
.Y(n_5739)
);

NOR2xp33_ASAP7_75t_L g5740 ( 
.A(n_3931),
.B(n_3845),
.Y(n_5740)
);

O2A1O1Ixp33_ASAP7_75t_L g5741 ( 
.A1(n_3961),
.A2(n_3962),
.B(n_3965),
.C(n_3964),
.Y(n_5741)
);

NAND2xp5_ASAP7_75t_SL g5742 ( 
.A(n_4010),
.B(n_4085),
.Y(n_5742)
);

OAI22xp5_ASAP7_75t_L g5743 ( 
.A1(n_3777),
.A2(n_3932),
.B1(n_3835),
.B2(n_3858),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_3514),
.B(n_3519),
.Y(n_5744)
);

NOR2xp33_ASAP7_75t_L g5745 ( 
.A(n_3845),
.B(n_3866),
.Y(n_5745)
);

O2A1O1Ixp33_ASAP7_75t_L g5746 ( 
.A1(n_3962),
.A2(n_3964),
.B(n_3969),
.C(n_3965),
.Y(n_5746)
);

NOR2xp67_ASAP7_75t_L g5747 ( 
.A(n_4530),
.B(n_4536),
.Y(n_5747)
);

INVx1_ASAP7_75t_L g5748 ( 
.A(n_4536),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_4538),
.Y(n_5749)
);

AOI21xp5_ASAP7_75t_L g5750 ( 
.A1(n_4543),
.A2(n_4659),
.B(n_4612),
.Y(n_5750)
);

A2O1A1Ixp33_ASAP7_75t_L g5751 ( 
.A1(n_4110),
.A2(n_4607),
.B(n_4621),
.C(n_4476),
.Y(n_5751)
);

BUFx6f_ASAP7_75t_L g5752 ( 
.A(n_3647),
.Y(n_5752)
);

NOR2xp33_ASAP7_75t_L g5753 ( 
.A(n_3845),
.B(n_3866),
.Y(n_5753)
);

AOI21xp5_ASAP7_75t_L g5754 ( 
.A1(n_4543),
.A2(n_4659),
.B(n_4612),
.Y(n_5754)
);

OAI22xp5_ASAP7_75t_L g5755 ( 
.A1(n_3777),
.A2(n_3932),
.B1(n_3835),
.B2(n_3858),
.Y(n_5755)
);

CKINVDCx6p67_ASAP7_75t_R g5756 ( 
.A(n_3662),
.Y(n_5756)
);

INVx1_ASAP7_75t_SL g5757 ( 
.A(n_4106),
.Y(n_5757)
);

NAND2xp5_ASAP7_75t_SL g5758 ( 
.A(n_4010),
.B(n_4017),
.Y(n_5758)
);

OAI21xp5_ASAP7_75t_L g5759 ( 
.A1(n_3519),
.A2(n_3534),
.B(n_3532),
.Y(n_5759)
);

OAI21xp5_ASAP7_75t_L g5760 ( 
.A1(n_3532),
.A2(n_3549),
.B(n_3534),
.Y(n_5760)
);

AOI21xp33_ASAP7_75t_L g5761 ( 
.A1(n_3532),
.A2(n_3549),
.B(n_3534),
.Y(n_5761)
);

OAI22xp5_ASAP7_75t_L g5762 ( 
.A1(n_3835),
.A2(n_3932),
.B1(n_3974),
.B2(n_3969),
.Y(n_5762)
);

INVx2_ASAP7_75t_L g5763 ( 
.A(n_3647),
.Y(n_5763)
);

OAI21xp5_ASAP7_75t_L g5764 ( 
.A1(n_3549),
.A2(n_3584),
.B(n_3555),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_4538),
.Y(n_5765)
);

A2O1A1Ixp33_ASAP7_75t_L g5766 ( 
.A1(n_4110),
.A2(n_4634),
.B(n_4683),
.C(n_4621),
.Y(n_5766)
);

O2A1O1Ixp33_ASAP7_75t_L g5767 ( 
.A1(n_3974),
.A2(n_3982),
.B(n_3993),
.C(n_3990),
.Y(n_5767)
);

NAND2xp5_ASAP7_75t_L g5768 ( 
.A(n_3555),
.B(n_3584),
.Y(n_5768)
);

AOI21xp5_ASAP7_75t_L g5769 ( 
.A1(n_4543),
.A2(n_4659),
.B(n_4612),
.Y(n_5769)
);

NOR2xp33_ASAP7_75t_L g5770 ( 
.A(n_3845),
.B(n_3866),
.Y(n_5770)
);

AO32x1_ASAP7_75t_L g5771 ( 
.A1(n_4540),
.A2(n_4552),
.A3(n_4559),
.B1(n_4547),
.B2(n_4546),
.Y(n_5771)
);

NOR2xp33_ASAP7_75t_L g5772 ( 
.A(n_3845),
.B(n_3866),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_3647),
.Y(n_5773)
);

NOR2xp33_ASAP7_75t_L g5774 ( 
.A(n_3866),
.B(n_3568),
.Y(n_5774)
);

AO32x1_ASAP7_75t_L g5775 ( 
.A1(n_4540),
.A2(n_4552),
.A3(n_4559),
.B1(n_4547),
.B2(n_4546),
.Y(n_5775)
);

NAND2xp5_ASAP7_75t_SL g5776 ( 
.A(n_4010),
.B(n_4017),
.Y(n_5776)
);

INVx3_ASAP7_75t_L g5777 ( 
.A(n_3345),
.Y(n_5777)
);

NAND2xp5_ASAP7_75t_L g5778 ( 
.A(n_3555),
.B(n_3584),
.Y(n_5778)
);

OAI21x1_ASAP7_75t_L g5779 ( 
.A1(n_4294),
.A2(n_4689),
.B(n_4686),
.Y(n_5779)
);

A2O1A1Ixp33_ASAP7_75t_L g5780 ( 
.A1(n_4110),
.A2(n_4634),
.B(n_4683),
.C(n_4621),
.Y(n_5780)
);

NAND2xp5_ASAP7_75t_SL g5781 ( 
.A(n_4010),
.B(n_3439),
.Y(n_5781)
);

AOI21xp5_ASAP7_75t_L g5782 ( 
.A1(n_4612),
.A2(n_4665),
.B(n_4659),
.Y(n_5782)
);

AND2x2_ASAP7_75t_L g5783 ( 
.A(n_3647),
.B(n_3669),
.Y(n_5783)
);

O2A1O1Ixp33_ASAP7_75t_L g5784 ( 
.A1(n_3982),
.A2(n_3990),
.B(n_3994),
.C(n_3993),
.Y(n_5784)
);

NAND2xp5_ASAP7_75t_SL g5785 ( 
.A(n_4010),
.B(n_3439),
.Y(n_5785)
);

AOI21xp5_ASAP7_75t_L g5786 ( 
.A1(n_4659),
.A2(n_4665),
.B(n_4156),
.Y(n_5786)
);

AOI21xp5_ASAP7_75t_L g5787 ( 
.A1(n_4659),
.A2(n_4665),
.B(n_4156),
.Y(n_5787)
);

INVx2_ASAP7_75t_L g5788 ( 
.A(n_3669),
.Y(n_5788)
);

NAND2xp5_ASAP7_75t_L g5789 ( 
.A(n_3586),
.B(n_3587),
.Y(n_5789)
);

AND2x4_ASAP7_75t_L g5790 ( 
.A(n_3345),
.B(n_3351),
.Y(n_5790)
);

AOI21xp5_ASAP7_75t_L g5791 ( 
.A1(n_4659),
.A2(n_4665),
.B(n_4156),
.Y(n_5791)
);

BUFx6f_ASAP7_75t_L g5792 ( 
.A(n_3669),
.Y(n_5792)
);

NAND2xp5_ASAP7_75t_L g5793 ( 
.A(n_3586),
.B(n_3587),
.Y(n_5793)
);

AOI22xp33_ASAP7_75t_L g5794 ( 
.A1(n_3364),
.A2(n_4683),
.B1(n_4634),
.B2(n_3332),
.Y(n_5794)
);

A2O1A1Ixp33_ASAP7_75t_L g5795 ( 
.A1(n_3817),
.A2(n_3937),
.B(n_4670),
.C(n_3431),
.Y(n_5795)
);

BUFx6f_ASAP7_75t_L g5796 ( 
.A(n_3669),
.Y(n_5796)
);

AOI21xp5_ASAP7_75t_L g5797 ( 
.A1(n_4659),
.A2(n_4665),
.B(n_4170),
.Y(n_5797)
);

A2O1A1Ixp33_ASAP7_75t_L g5798 ( 
.A1(n_3817),
.A2(n_3937),
.B(n_4670),
.C(n_3431),
.Y(n_5798)
);

O2A1O1Ixp5_ASAP7_75t_L g5799 ( 
.A1(n_4575),
.A2(n_4579),
.B(n_4594),
.C(n_4576),
.Y(n_5799)
);

NOR2xp33_ASAP7_75t_L g5800 ( 
.A(n_3568),
.B(n_3619),
.Y(n_5800)
);

NAND3xp33_ASAP7_75t_L g5801 ( 
.A(n_3994),
.B(n_4029),
.C(n_4002),
.Y(n_5801)
);

AND2x2_ASAP7_75t_L g5802 ( 
.A(n_3669),
.B(n_3702),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_4575),
.Y(n_5803)
);

NOR2xp33_ASAP7_75t_L g5804 ( 
.A(n_3568),
.B(n_3619),
.Y(n_5804)
);

BUFx3_ASAP7_75t_L g5805 ( 
.A(n_4047),
.Y(n_5805)
);

CKINVDCx5p33_ASAP7_75t_R g5806 ( 
.A(n_4257),
.Y(n_5806)
);

OAI21xp5_ASAP7_75t_L g5807 ( 
.A1(n_3591),
.A2(n_3606),
.B(n_3604),
.Y(n_5807)
);

INVx5_ASAP7_75t_L g5808 ( 
.A(n_4665),
.Y(n_5808)
);

AOI21xp5_ASAP7_75t_L g5809 ( 
.A1(n_4154),
.A2(n_4173),
.B(n_4172),
.Y(n_5809)
);

AND2x2_ASAP7_75t_L g5810 ( 
.A(n_3669),
.B(n_3702),
.Y(n_5810)
);

INVx2_ASAP7_75t_L g5811 ( 
.A(n_3669),
.Y(n_5811)
);

INVx2_ASAP7_75t_L g5812 ( 
.A(n_3669),
.Y(n_5812)
);

AOI21xp5_ASAP7_75t_L g5813 ( 
.A1(n_4172),
.A2(n_4196),
.B(n_4173),
.Y(n_5813)
);

AOI21xp5_ASAP7_75t_L g5814 ( 
.A1(n_4172),
.A2(n_4196),
.B(n_4173),
.Y(n_5814)
);

INVx4_ASAP7_75t_L g5815 ( 
.A(n_4047),
.Y(n_5815)
);

OA21x2_ASAP7_75t_L g5816 ( 
.A1(n_4576),
.A2(n_4594),
.B(n_4579),
.Y(n_5816)
);

AOI22xp5_ASAP7_75t_L g5817 ( 
.A1(n_3957),
.A2(n_3920),
.B1(n_4147),
.B2(n_3512),
.Y(n_5817)
);

AOI21xp5_ASAP7_75t_L g5818 ( 
.A1(n_4196),
.A2(n_4228),
.B(n_4221),
.Y(n_5818)
);

AOI22xp5_ASAP7_75t_L g5819 ( 
.A1(n_3920),
.A2(n_4147),
.B1(n_3512),
.B2(n_3544),
.Y(n_5819)
);

NAND2xp5_ASAP7_75t_L g5820 ( 
.A(n_3591),
.B(n_3604),
.Y(n_5820)
);

AOI21xp5_ASAP7_75t_L g5821 ( 
.A1(n_4221),
.A2(n_4237),
.B(n_4228),
.Y(n_5821)
);

NOR2xp33_ASAP7_75t_L g5822 ( 
.A(n_3568),
.B(n_3619),
.Y(n_5822)
);

NOR2xp33_ASAP7_75t_L g5823 ( 
.A(n_3568),
.B(n_3619),
.Y(n_5823)
);

AOI21xp5_ASAP7_75t_L g5824 ( 
.A1(n_4221),
.A2(n_4237),
.B(n_4228),
.Y(n_5824)
);

BUFx3_ASAP7_75t_L g5825 ( 
.A(n_4047),
.Y(n_5825)
);

INVxp67_ASAP7_75t_L g5826 ( 
.A(n_3793),
.Y(n_5826)
);

INVx2_ASAP7_75t_L g5827 ( 
.A(n_3702),
.Y(n_5827)
);

NAND2xp5_ASAP7_75t_L g5828 ( 
.A(n_3606),
.B(n_3612),
.Y(n_5828)
);

A2O1A1Ixp33_ASAP7_75t_L g5829 ( 
.A1(n_3431),
.A2(n_3590),
.B(n_3650),
.C(n_3544),
.Y(n_5829)
);

OAI22xp5_ASAP7_75t_L g5830 ( 
.A1(n_4002),
.A2(n_4030),
.B1(n_4029),
.B2(n_3831),
.Y(n_5830)
);

AO22x1_ASAP7_75t_L g5831 ( 
.A1(n_3626),
.A2(n_4037),
.B1(n_3707),
.B2(n_3411),
.Y(n_5831)
);

NAND2xp5_ASAP7_75t_L g5832 ( 
.A(n_3606),
.B(n_3612),
.Y(n_5832)
);

OAI21xp5_ASAP7_75t_L g5833 ( 
.A1(n_3612),
.A2(n_3645),
.B(n_3627),
.Y(n_5833)
);

BUFx3_ASAP7_75t_L g5834 ( 
.A(n_4106),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_4597),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_4597),
.Y(n_5836)
);

A2O1A1Ixp33_ASAP7_75t_L g5837 ( 
.A1(n_3544),
.A2(n_3650),
.B(n_3654),
.C(n_3590),
.Y(n_5837)
);

NOR2xp33_ASAP7_75t_L g5838 ( 
.A(n_3619),
.B(n_3638),
.Y(n_5838)
);

INVx5_ASAP7_75t_L g5839 ( 
.A(n_3254),
.Y(n_5839)
);

INVx4_ASAP7_75t_L g5840 ( 
.A(n_3448),
.Y(n_5840)
);

O2A1O1Ixp33_ASAP7_75t_L g5841 ( 
.A1(n_4030),
.A2(n_4139),
.B(n_4150),
.C(n_4146),
.Y(n_5841)
);

NAND2xp5_ASAP7_75t_SL g5842 ( 
.A(n_3439),
.B(n_4583),
.Y(n_5842)
);

NAND2xp5_ASAP7_75t_L g5843 ( 
.A(n_3627),
.B(n_3645),
.Y(n_5843)
);

HB1xp67_ASAP7_75t_L g5844 ( 
.A(n_4106),
.Y(n_5844)
);

NAND2xp33_ASAP7_75t_L g5845 ( 
.A(n_3425),
.B(n_3452),
.Y(n_5845)
);

BUFx3_ASAP7_75t_L g5846 ( 
.A(n_3626),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_4609),
.Y(n_5847)
);

INVx3_ASAP7_75t_L g5848 ( 
.A(n_3351),
.Y(n_5848)
);

CKINVDCx10_ASAP7_75t_R g5849 ( 
.A(n_3920),
.Y(n_5849)
);

NAND2xp5_ASAP7_75t_SL g5850 ( 
.A(n_3439),
.B(n_4112),
.Y(n_5850)
);

NOR2xp33_ASAP7_75t_L g5851 ( 
.A(n_3638),
.B(n_3684),
.Y(n_5851)
);

AND2x2_ASAP7_75t_L g5852 ( 
.A(n_3702),
.B(n_3739),
.Y(n_5852)
);

INVxp67_ASAP7_75t_L g5853 ( 
.A(n_3793),
.Y(n_5853)
);

OAI22xp5_ASAP7_75t_L g5854 ( 
.A1(n_3826),
.A2(n_3833),
.B1(n_3847),
.B2(n_3831),
.Y(n_5854)
);

NOR3xp33_ASAP7_75t_L g5855 ( 
.A(n_4148),
.B(n_4146),
.C(n_4139),
.Y(n_5855)
);

NOR2xp33_ASAP7_75t_L g5856 ( 
.A(n_3638),
.B(n_3684),
.Y(n_5856)
);

AOI22xp33_ASAP7_75t_L g5857 ( 
.A1(n_3364),
.A2(n_3332),
.B1(n_3399),
.B2(n_3292),
.Y(n_5857)
);

NAND2xp5_ASAP7_75t_L g5858 ( 
.A(n_3627),
.B(n_3645),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_4609),
.Y(n_5859)
);

NAND2xp5_ASAP7_75t_L g5860 ( 
.A(n_3646),
.B(n_3649),
.Y(n_5860)
);

NAND2xp5_ASAP7_75t_L g5861 ( 
.A(n_3646),
.B(n_3649),
.Y(n_5861)
);

NAND2xp5_ASAP7_75t_L g5862 ( 
.A(n_3646),
.B(n_3649),
.Y(n_5862)
);

INVx3_ASAP7_75t_L g5863 ( 
.A(n_3351),
.Y(n_5863)
);

NOR3xp33_ASAP7_75t_L g5864 ( 
.A(n_4139),
.B(n_4150),
.C(n_4146),
.Y(n_5864)
);

BUFx12f_ASAP7_75t_L g5865 ( 
.A(n_3415),
.Y(n_5865)
);

NAND2xp5_ASAP7_75t_L g5866 ( 
.A(n_3689),
.B(n_3690),
.Y(n_5866)
);

OA22x2_ASAP7_75t_L g5867 ( 
.A1(n_3367),
.A2(n_3654),
.B1(n_3688),
.B2(n_3650),
.Y(n_5867)
);

NAND2xp5_ASAP7_75t_L g5868 ( 
.A(n_3689),
.B(n_3690),
.Y(n_5868)
);

NOR2xp33_ASAP7_75t_L g5869 ( 
.A(n_3638),
.B(n_3684),
.Y(n_5869)
);

AOI21xp5_ASAP7_75t_L g5870 ( 
.A1(n_4263),
.A2(n_4270),
.B(n_4267),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_SL g5871 ( 
.A(n_3439),
.B(n_4112),
.Y(n_5871)
);

AOI21xp5_ASAP7_75t_L g5872 ( 
.A1(n_4270),
.A2(n_4308),
.B(n_4286),
.Y(n_5872)
);

INVx1_ASAP7_75t_L g5873 ( 
.A(n_4615),
.Y(n_5873)
);

NOR2xp33_ASAP7_75t_L g5874 ( 
.A(n_3638),
.B(n_3684),
.Y(n_5874)
);

AND2x4_ASAP7_75t_L g5875 ( 
.A(n_3351),
.B(n_3373),
.Y(n_5875)
);

OR2x6_ASAP7_75t_SL g5876 ( 
.A(n_3689),
.B(n_3690),
.Y(n_5876)
);

NOR2xp33_ASAP7_75t_L g5877 ( 
.A(n_3684),
.B(n_3721),
.Y(n_5877)
);

NAND2xp5_ASAP7_75t_L g5878 ( 
.A(n_3705),
.B(n_3737),
.Y(n_5878)
);

AO32x2_ASAP7_75t_L g5879 ( 
.A1(n_3654),
.A2(n_3688),
.A3(n_3779),
.B1(n_3693),
.B2(n_3342),
.Y(n_5879)
);

OAI21xp5_ASAP7_75t_L g5880 ( 
.A1(n_3705),
.A2(n_3749),
.B(n_3737),
.Y(n_5880)
);

BUFx8_ASAP7_75t_L g5881 ( 
.A(n_3457),
.Y(n_5881)
);

NOR2x1_ASAP7_75t_L g5882 ( 
.A(n_3380),
.B(n_3411),
.Y(n_5882)
);

A2O1A1Ixp33_ASAP7_75t_L g5883 ( 
.A1(n_3688),
.A2(n_3693),
.B(n_3779),
.C(n_3602),
.Y(n_5883)
);

NAND2xp5_ASAP7_75t_L g5884 ( 
.A(n_3705),
.B(n_3737),
.Y(n_5884)
);

NOR2xp33_ASAP7_75t_L g5885 ( 
.A(n_3721),
.B(n_3762),
.Y(n_5885)
);

INVx11_ASAP7_75t_L g5886 ( 
.A(n_3707),
.Y(n_5886)
);

OAI21xp5_ASAP7_75t_L g5887 ( 
.A1(n_3749),
.A2(n_3770),
.B(n_3765),
.Y(n_5887)
);

AOI21xp5_ASAP7_75t_L g5888 ( 
.A1(n_4286),
.A2(n_4312),
.B(n_4308),
.Y(n_5888)
);

OAI21xp5_ASAP7_75t_L g5889 ( 
.A1(n_3749),
.A2(n_3821),
.B(n_3778),
.Y(n_5889)
);

OAI21xp5_ASAP7_75t_L g5890 ( 
.A1(n_4615),
.A2(n_4629),
.B(n_4623),
.Y(n_5890)
);

NAND2xp5_ASAP7_75t_L g5891 ( 
.A(n_3794),
.B(n_3693),
.Y(n_5891)
);

NAND2xp5_ASAP7_75t_SL g5892 ( 
.A(n_4112),
.B(n_3872),
.Y(n_5892)
);

NAND2xp5_ASAP7_75t_L g5893 ( 
.A(n_3794),
.B(n_3779),
.Y(n_5893)
);

INVx3_ASAP7_75t_L g5894 ( 
.A(n_3373),
.Y(n_5894)
);

BUFx2_ASAP7_75t_L g5895 ( 
.A(n_3702),
.Y(n_5895)
);

NAND2xp5_ASAP7_75t_SL g5896 ( 
.A(n_3872),
.B(n_3882),
.Y(n_5896)
);

NAND2xp5_ASAP7_75t_L g5897 ( 
.A(n_3702),
.B(n_3739),
.Y(n_5897)
);

CKINVDCx5p33_ASAP7_75t_R g5898 ( 
.A(n_4264),
.Y(n_5898)
);

NAND2xp5_ASAP7_75t_L g5899 ( 
.A(n_3739),
.B(n_4043),
.Y(n_5899)
);

OAI21xp5_ASAP7_75t_L g5900 ( 
.A1(n_4623),
.A2(n_4630),
.B(n_4629),
.Y(n_5900)
);

O2A1O1Ixp33_ASAP7_75t_SL g5901 ( 
.A1(n_4129),
.A2(n_4133),
.B(n_4138),
.C(n_4131),
.Y(n_5901)
);

A2O1A1Ixp33_ASAP7_75t_L g5902 ( 
.A1(n_3602),
.A2(n_3884),
.B(n_3876),
.C(n_3340),
.Y(n_5902)
);

NAND2xp5_ASAP7_75t_L g5903 ( 
.A(n_3739),
.B(n_4043),
.Y(n_5903)
);

HB1xp67_ASAP7_75t_L g5904 ( 
.A(n_3739),
.Y(n_5904)
);

AOI21xp5_ASAP7_75t_L g5905 ( 
.A1(n_4286),
.A2(n_4312),
.B(n_4308),
.Y(n_5905)
);

AO22x1_ASAP7_75t_L g5906 ( 
.A1(n_3707),
.A2(n_4037),
.B1(n_3411),
.B2(n_3380),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_4630),
.Y(n_5907)
);

AOI21x1_ASAP7_75t_L g5908 ( 
.A1(n_4633),
.A2(n_4651),
.B(n_4640),
.Y(n_5908)
);

BUFx3_ASAP7_75t_L g5909 ( 
.A(n_3707),
.Y(n_5909)
);

CKINVDCx10_ASAP7_75t_R g5910 ( 
.A(n_3891),
.Y(n_5910)
);

INVx3_ASAP7_75t_L g5911 ( 
.A(n_3373),
.Y(n_5911)
);

AOI21xp5_ASAP7_75t_L g5912 ( 
.A1(n_4312),
.A2(n_4332),
.B(n_4318),
.Y(n_5912)
);

NAND2xp5_ASAP7_75t_L g5913 ( 
.A(n_3739),
.B(n_4050),
.Y(n_5913)
);

INVx2_ASAP7_75t_L g5914 ( 
.A(n_3739),
.Y(n_5914)
);

AOI21x1_ASAP7_75t_L g5915 ( 
.A1(n_4633),
.A2(n_4651),
.B(n_4640),
.Y(n_5915)
);

NOR2xp33_ASAP7_75t_SL g5916 ( 
.A(n_3385),
.B(n_3380),
.Y(n_5916)
);

NAND2xp5_ASAP7_75t_SL g5917 ( 
.A(n_3872),
.B(n_3882),
.Y(n_5917)
);

NOR3xp33_ASAP7_75t_L g5918 ( 
.A(n_4150),
.B(n_4142),
.C(n_4141),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_4653),
.Y(n_5919)
);

AOI21x1_ASAP7_75t_L g5920 ( 
.A1(n_4653),
.A2(n_4678),
.B(n_4676),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_3756),
.Y(n_5921)
);

A2O1A1Ixp33_ASAP7_75t_L g5922 ( 
.A1(n_3602),
.A2(n_3884),
.B(n_3876),
.C(n_3340),
.Y(n_5922)
);

AOI21x1_ASAP7_75t_L g5923 ( 
.A1(n_4676),
.A2(n_4678),
.B(n_4332),
.Y(n_5923)
);

INVx2_ASAP7_75t_L g5924 ( 
.A(n_3756),
.Y(n_5924)
);

AND2x6_ASAP7_75t_L g5925 ( 
.A(n_3254),
.B(n_3274),
.Y(n_5925)
);

NAND2xp5_ASAP7_75t_L g5926 ( 
.A(n_4050),
.B(n_4054),
.Y(n_5926)
);

AOI22xp5_ASAP7_75t_L g5927 ( 
.A1(n_4147),
.A2(n_4136),
.B1(n_3890),
.B2(n_3941),
.Y(n_5927)
);

NAND2xp5_ASAP7_75t_L g5928 ( 
.A(n_4054),
.B(n_3756),
.Y(n_5928)
);

NAND2xp5_ASAP7_75t_L g5929 ( 
.A(n_3756),
.B(n_3761),
.Y(n_5929)
);

OAI22xp5_ASAP7_75t_L g5930 ( 
.A1(n_3826),
.A2(n_3847),
.B1(n_3854),
.B2(n_3833),
.Y(n_5930)
);

NOR2x1_ASAP7_75t_L g5931 ( 
.A(n_3380),
.B(n_3411),
.Y(n_5931)
);

AOI22xp5_ASAP7_75t_L g5932 ( 
.A1(n_4147),
.A2(n_4136),
.B1(n_3890),
.B2(n_3941),
.Y(n_5932)
);

AOI33xp33_ASAP7_75t_L g5933 ( 
.A1(n_4141),
.A2(n_4145),
.A3(n_4142),
.B1(n_4118),
.B2(n_4123),
.B3(n_4127),
.Y(n_5933)
);

BUFx6f_ASAP7_75t_L g5934 ( 
.A(n_3756),
.Y(n_5934)
);

O2A1O1Ixp33_ASAP7_75t_L g5935 ( 
.A1(n_3951),
.A2(n_4078),
.B(n_4136),
.C(n_3855),
.Y(n_5935)
);

OAI21xp5_ASAP7_75t_L g5936 ( 
.A1(n_4053),
.A2(n_4197),
.B(n_4160),
.Y(n_5936)
);

AOI21xp5_ASAP7_75t_L g5937 ( 
.A1(n_4318),
.A2(n_4351),
.B(n_4332),
.Y(n_5937)
);

NOR2xp33_ASAP7_75t_L g5938 ( 
.A(n_3721),
.B(n_3762),
.Y(n_5938)
);

AOI21xp5_ASAP7_75t_L g5939 ( 
.A1(n_4318),
.A2(n_4364),
.B(n_4351),
.Y(n_5939)
);

NAND2xp5_ASAP7_75t_SL g5940 ( 
.A(n_3872),
.B(n_3882),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_3756),
.Y(n_5941)
);

NAND2xp5_ASAP7_75t_L g5942 ( 
.A(n_3756),
.B(n_3761),
.Y(n_5942)
);

NAND2xp5_ASAP7_75t_L g5943 ( 
.A(n_3761),
.B(n_3775),
.Y(n_5943)
);

A2O1A1Ixp33_ASAP7_75t_L g5944 ( 
.A1(n_3602),
.A2(n_3884),
.B(n_3876),
.C(n_3340),
.Y(n_5944)
);

NAND2xp5_ASAP7_75t_L g5945 ( 
.A(n_3775),
.B(n_3781),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_3292),
.B(n_3399),
.Y(n_5946)
);

AOI21xp5_ASAP7_75t_L g5947 ( 
.A1(n_4351),
.A2(n_4366),
.B(n_4364),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_3775),
.Y(n_5948)
);

AOI21xp5_ASAP7_75t_L g5949 ( 
.A1(n_4364),
.A2(n_4367),
.B(n_4366),
.Y(n_5949)
);

NAND2xp5_ASAP7_75t_SL g5950 ( 
.A(n_3872),
.B(n_3882),
.Y(n_5950)
);

AND2x2_ASAP7_75t_L g5951 ( 
.A(n_3373),
.B(n_4643),
.Y(n_5951)
);

A2O1A1Ixp33_ASAP7_75t_L g5952 ( 
.A1(n_3602),
.A2(n_3876),
.B(n_3884),
.C(n_3342),
.Y(n_5952)
);

AND2x2_ASAP7_75t_L g5953 ( 
.A(n_4643),
.B(n_3781),
.Y(n_5953)
);

NOR2xp33_ASAP7_75t_L g5954 ( 
.A(n_3721),
.B(n_3762),
.Y(n_5954)
);

AOI21xp5_ASAP7_75t_L g5955 ( 
.A1(n_4366),
.A2(n_4381),
.B(n_4367),
.Y(n_5955)
);

AOI221xp5_ASAP7_75t_L g5956 ( 
.A1(n_3951),
.A2(n_4143),
.B1(n_4145),
.B2(n_3859),
.C(n_3860),
.Y(n_5956)
);

OAI22xp5_ASAP7_75t_L g5957 ( 
.A1(n_3854),
.A2(n_3859),
.B1(n_3860),
.B2(n_3855),
.Y(n_5957)
);

NAND3xp33_ASAP7_75t_L g5958 ( 
.A(n_4078),
.B(n_4037),
.C(n_3890),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_4367),
.Y(n_5959)
);

NAND2xp5_ASAP7_75t_L g5960 ( 
.A(n_3781),
.B(n_3788),
.Y(n_5960)
);

NAND2xp5_ASAP7_75t_SL g5961 ( 
.A(n_3882),
.B(n_3950),
.Y(n_5961)
);

AOI21xp5_ASAP7_75t_L g5962 ( 
.A1(n_4381),
.A2(n_4393),
.B(n_4388),
.Y(n_5962)
);

NAND2xp33_ASAP7_75t_L g5963 ( 
.A(n_3487),
.B(n_3504),
.Y(n_5963)
);

BUFx4f_ASAP7_75t_L g5964 ( 
.A(n_3448),
.Y(n_5964)
);

AND2x4_ASAP7_75t_L g5965 ( 
.A(n_3254),
.B(n_3274),
.Y(n_5965)
);

A2O1A1Ixp33_ASAP7_75t_L g5966 ( 
.A1(n_3876),
.A2(n_3884),
.B(n_3342),
.C(n_4078),
.Y(n_5966)
);

AOI22x1_ASAP7_75t_L g5967 ( 
.A1(n_3995),
.A2(n_3849),
.B1(n_3867),
.B2(n_3793),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_3788),
.Y(n_5968)
);

AND2x2_ASAP7_75t_SL g5969 ( 
.A(n_3274),
.B(n_3380),
.Y(n_5969)
);

NAND2xp5_ASAP7_75t_SL g5970 ( 
.A(n_3950),
.B(n_3983),
.Y(n_5970)
);

HB1xp67_ASAP7_75t_L g5971 ( 
.A(n_4075),
.Y(n_5971)
);

NAND2xp33_ASAP7_75t_L g5972 ( 
.A(n_3633),
.B(n_3655),
.Y(n_5972)
);

NOR2x1_ASAP7_75t_L g5973 ( 
.A(n_3411),
.B(n_3408),
.Y(n_5973)
);

NAND2xp5_ASAP7_75t_L g5974 ( 
.A(n_3788),
.B(n_3797),
.Y(n_5974)
);

BUFx6f_ASAP7_75t_L g5975 ( 
.A(n_3241),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_L g5976 ( 
.A(n_3797),
.B(n_3813),
.Y(n_5976)
);

AOI21xp5_ASAP7_75t_L g5977 ( 
.A1(n_4381),
.A2(n_4393),
.B(n_4388),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_3797),
.Y(n_5978)
);

NOR2xp33_ASAP7_75t_R g5979 ( 
.A(n_4328),
.B(n_4357),
.Y(n_5979)
);

OAI21xp5_ASAP7_75t_L g5980 ( 
.A1(n_4053),
.A2(n_4197),
.B(n_4160),
.Y(n_5980)
);

AOI21xp5_ASAP7_75t_L g5981 ( 
.A1(n_4388),
.A2(n_4408),
.B(n_4393),
.Y(n_5981)
);

OAI321xp33_ASAP7_75t_L g5982 ( 
.A1(n_4057),
.A2(n_3889),
.A3(n_3867),
.B1(n_3895),
.B2(n_3887),
.C(n_3849),
.Y(n_5982)
);

NAND2xp5_ASAP7_75t_L g5983 ( 
.A(n_3813),
.B(n_3834),
.Y(n_5983)
);

AOI21xp5_ASAP7_75t_L g5984 ( 
.A1(n_4408),
.A2(n_4434),
.B(n_4410),
.Y(n_5984)
);

AOI21x1_ASAP7_75t_L g5985 ( 
.A1(n_4408),
.A2(n_4434),
.B(n_4410),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_3813),
.Y(n_5986)
);

BUFx8_ASAP7_75t_L g5987 ( 
.A(n_3457),
.Y(n_5987)
);

NOR2xp33_ASAP7_75t_L g5988 ( 
.A(n_3721),
.B(n_3762),
.Y(n_5988)
);

NOR2xp33_ASAP7_75t_L g5989 ( 
.A(n_3762),
.B(n_3828),
.Y(n_5989)
);

BUFx6f_ASAP7_75t_L g5990 ( 
.A(n_3241),
.Y(n_5990)
);

INVx2_ASAP7_75t_L g5991 ( 
.A(n_4410),
.Y(n_5991)
);

AND2x2_ASAP7_75t_L g5992 ( 
.A(n_4643),
.B(n_3834),
.Y(n_5992)
);

INVx1_ASAP7_75t_L g5993 ( 
.A(n_3834),
.Y(n_5993)
);

NAND2xp5_ASAP7_75t_L g5994 ( 
.A(n_3837),
.B(n_3844),
.Y(n_5994)
);

NAND3xp33_ASAP7_75t_L g5995 ( 
.A(n_4037),
.B(n_3941),
.C(n_3795),
.Y(n_5995)
);

AOI21xp5_ASAP7_75t_L g5996 ( 
.A1(n_4437),
.A2(n_4484),
.B(n_4440),
.Y(n_5996)
);

OAI21xp5_ASAP7_75t_L g5997 ( 
.A1(n_4053),
.A2(n_4321),
.B(n_4262),
.Y(n_5997)
);

AND2x4_ASAP7_75t_L g5998 ( 
.A(n_4233),
.B(n_4272),
.Y(n_5998)
);

AND2x2_ASAP7_75t_L g5999 ( 
.A(n_4643),
.B(n_3837),
.Y(n_5999)
);

NAND2xp5_ASAP7_75t_SL g6000 ( 
.A(n_3950),
.B(n_3983),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_3837),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_L g6002 ( 
.A(n_3844),
.B(n_3848),
.Y(n_6002)
);

INVx1_ASAP7_75t_L g6003 ( 
.A(n_3844),
.Y(n_6003)
);

AOI21xp5_ASAP7_75t_L g6004 ( 
.A1(n_4437),
.A2(n_4484),
.B(n_4440),
.Y(n_6004)
);

INVx2_ASAP7_75t_L g6005 ( 
.A(n_4437),
.Y(n_6005)
);

AND2x2_ASAP7_75t_SL g6006 ( 
.A(n_3241),
.B(n_4009),
.Y(n_6006)
);

O2A1O1Ixp33_ASAP7_75t_L g6007 ( 
.A1(n_3864),
.A2(n_3888),
.B(n_3870),
.C(n_4143),
.Y(n_6007)
);

AO22x1_ASAP7_75t_L g6008 ( 
.A1(n_4037),
.A2(n_3968),
.B1(n_3880),
.B2(n_3877),
.Y(n_6008)
);

INVx2_ASAP7_75t_L g6009 ( 
.A(n_4440),
.Y(n_6009)
);

OA22x2_ASAP7_75t_L g6010 ( 
.A1(n_4233),
.A2(n_4272),
.B1(n_4316),
.B2(n_4289),
.Y(n_6010)
);

CKINVDCx5p33_ASAP7_75t_R g6011 ( 
.A(n_4415),
.Y(n_6011)
);

AOI21xp5_ASAP7_75t_L g6012 ( 
.A1(n_4484),
.A2(n_4492),
.B(n_4486),
.Y(n_6012)
);

NAND2xp5_ASAP7_75t_SL g6013 ( 
.A(n_3950),
.B(n_3983),
.Y(n_6013)
);

NAND2xp5_ASAP7_75t_L g6014 ( 
.A(n_3848),
.B(n_3897),
.Y(n_6014)
);

AOI21xp5_ASAP7_75t_L g6015 ( 
.A1(n_4486),
.A2(n_4499),
.B(n_4492),
.Y(n_6015)
);

NAND2xp5_ASAP7_75t_SL g6016 ( 
.A(n_3950),
.B(n_3983),
.Y(n_6016)
);

AOI21xp5_ASAP7_75t_L g6017 ( 
.A1(n_4486),
.A2(n_4499),
.B(n_4492),
.Y(n_6017)
);

INVx2_ASAP7_75t_L g6018 ( 
.A(n_4499),
.Y(n_6018)
);

AOI21xp5_ASAP7_75t_L g6019 ( 
.A1(n_4503),
.A2(n_4510),
.B(n_4505),
.Y(n_6019)
);

INVxp67_ASAP7_75t_L g6020 ( 
.A(n_3849),
.Y(n_6020)
);

AOI21xp5_ASAP7_75t_L g6021 ( 
.A1(n_4503),
.A2(n_4510),
.B(n_4505),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_3897),
.Y(n_6022)
);

NAND3xp33_ASAP7_75t_SL g6023 ( 
.A(n_3455),
.B(n_4118),
.C(n_4117),
.Y(n_6023)
);

AOI21xp5_ASAP7_75t_L g6024 ( 
.A1(n_4503),
.A2(n_4510),
.B(n_4505),
.Y(n_6024)
);

BUFx3_ASAP7_75t_L g6025 ( 
.A(n_3448),
.Y(n_6025)
);

OR2x6_ASAP7_75t_L g6026 ( 
.A(n_4513),
.B(n_4519),
.Y(n_6026)
);

OAI21x1_ASAP7_75t_L g6027 ( 
.A1(n_4340),
.A2(n_4406),
.B(n_4341),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_4643),
.B(n_4513),
.Y(n_6028)
);

AOI22x1_ASAP7_75t_L g6029 ( 
.A1(n_3995),
.A2(n_3887),
.B1(n_3889),
.B2(n_3867),
.Y(n_6029)
);

AOI21xp5_ASAP7_75t_L g6030 ( 
.A1(n_4513),
.A2(n_4522),
.B(n_4519),
.Y(n_6030)
);

AOI21xp5_ASAP7_75t_L g6031 ( 
.A1(n_4519),
.A2(n_4523),
.B(n_4522),
.Y(n_6031)
);

INVx1_ASAP7_75t_L g6032 ( 
.A(n_3736),
.Y(n_6032)
);

AOI21xp5_ASAP7_75t_L g6033 ( 
.A1(n_4522),
.A2(n_4525),
.B(n_4523),
.Y(n_6033)
);

INVx1_ASAP7_75t_L g6034 ( 
.A(n_3736),
.Y(n_6034)
);

NOR2xp33_ASAP7_75t_L g6035 ( 
.A(n_3828),
.B(n_3843),
.Y(n_6035)
);

NOR2xp33_ASAP7_75t_L g6036 ( 
.A(n_3828),
.B(n_3843),
.Y(n_6036)
);

OAI321xp33_ASAP7_75t_L g6037 ( 
.A1(n_4057),
.A2(n_3889),
.A3(n_3895),
.B1(n_3887),
.B2(n_3888),
.C(n_3870),
.Y(n_6037)
);

NAND2xp5_ASAP7_75t_SL g6038 ( 
.A(n_3983),
.B(n_3508),
.Y(n_6038)
);

NOR2xp67_ASAP7_75t_L g6039 ( 
.A(n_3277),
.B(n_3327),
.Y(n_6039)
);

A2O1A1Ixp33_ASAP7_75t_L g6040 ( 
.A1(n_4117),
.A2(n_3240),
.B(n_4155),
.C(n_3245),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_3736),
.Y(n_6041)
);

NAND3xp33_ASAP7_75t_L g6042 ( 
.A(n_3795),
.B(n_3949),
.C(n_4102),
.Y(n_6042)
);

INVxp33_ASAP7_75t_SL g6043 ( 
.A(n_4424),
.Y(n_6043)
);

OAI22xp5_ASAP7_75t_L g6044 ( 
.A1(n_3864),
.A2(n_3250),
.B1(n_3258),
.B2(n_3247),
.Y(n_6044)
);

AOI21xp5_ASAP7_75t_L g6045 ( 
.A1(n_4523),
.A2(n_4539),
.B(n_4525),
.Y(n_6045)
);

BUFx3_ASAP7_75t_L g6046 ( 
.A(n_3448),
.Y(n_6046)
);

AOI21xp5_ASAP7_75t_L g6047 ( 
.A1(n_4525),
.A2(n_4550),
.B(n_4539),
.Y(n_6047)
);

AO32x1_ASAP7_75t_L g6048 ( 
.A1(n_4539),
.A2(n_4590),
.A3(n_4606),
.B1(n_4574),
.B2(n_4550),
.Y(n_6048)
);

NAND2xp5_ASAP7_75t_L g6049 ( 
.A(n_3247),
.B(n_3250),
.Y(n_6049)
);

AOI21xp5_ASAP7_75t_L g6050 ( 
.A1(n_4550),
.A2(n_4590),
.B(n_4574),
.Y(n_6050)
);

NAND2xp5_ASAP7_75t_L g6051 ( 
.A(n_3258),
.B(n_3262),
.Y(n_6051)
);

NAND2xp5_ASAP7_75t_SL g6052 ( 
.A(n_3508),
.B(n_3523),
.Y(n_6052)
);

A2O1A1Ixp33_ASAP7_75t_L g6053 ( 
.A1(n_4117),
.A2(n_3240),
.B(n_4155),
.C(n_3245),
.Y(n_6053)
);

AOI21xp5_ASAP7_75t_L g6054 ( 
.A1(n_4574),
.A2(n_4606),
.B(n_4590),
.Y(n_6054)
);

NAND2xp5_ASAP7_75t_L g6055 ( 
.A(n_3262),
.B(n_3271),
.Y(n_6055)
);

BUFx6f_ASAP7_75t_L g6056 ( 
.A(n_3241),
.Y(n_6056)
);

AOI21xp5_ASAP7_75t_L g6057 ( 
.A1(n_4606),
.A2(n_4642),
.B(n_4614),
.Y(n_6057)
);

NAND2xp5_ASAP7_75t_L g6058 ( 
.A(n_3271),
.B(n_3273),
.Y(n_6058)
);

AOI22xp33_ASAP7_75t_L g6059 ( 
.A1(n_4643),
.A2(n_3843),
.B1(n_3828),
.B2(n_4233),
.Y(n_6059)
);

NAND2xp5_ASAP7_75t_L g6060 ( 
.A(n_3273),
.B(n_3281),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_3736),
.Y(n_6061)
);

INVx4_ASAP7_75t_L g6062 ( 
.A(n_3448),
.Y(n_6062)
);

OAI21xp33_ASAP7_75t_L g6063 ( 
.A1(n_3455),
.A2(n_3933),
.B(n_3918),
.Y(n_6063)
);

INVx3_ASAP7_75t_L g6064 ( 
.A(n_3241),
.Y(n_6064)
);

AOI21xp33_ASAP7_75t_L g6065 ( 
.A1(n_3895),
.A2(n_3282),
.B(n_3281),
.Y(n_6065)
);

A2O1A1Ixp33_ASAP7_75t_L g6066 ( 
.A1(n_3240),
.A2(n_3245),
.B(n_4218),
.C(n_4155),
.Y(n_6066)
);

AOI21xp5_ASAP7_75t_L g6067 ( 
.A1(n_4614),
.A2(n_4657),
.B(n_4642),
.Y(n_6067)
);

O2A1O1Ixp33_ASAP7_75t_L g6068 ( 
.A1(n_4262),
.A2(n_4323),
.B(n_4327),
.C(n_4321),
.Y(n_6068)
);

NOR2xp33_ASAP7_75t_L g6069 ( 
.A(n_3828),
.B(n_3843),
.Y(n_6069)
);

AND2x4_ASAP7_75t_L g6070 ( 
.A(n_4233),
.B(n_4272),
.Y(n_6070)
);

NAND2xp5_ASAP7_75t_L g6071 ( 
.A(n_3282),
.B(n_3288),
.Y(n_6071)
);

OAI22xp5_ASAP7_75t_L g6072 ( 
.A1(n_3288),
.A2(n_3298),
.B1(n_3307),
.B2(n_3294),
.Y(n_6072)
);

NAND2xp5_ASAP7_75t_L g6073 ( 
.A(n_3294),
.B(n_3298),
.Y(n_6073)
);

HB1xp67_ASAP7_75t_L g6074 ( 
.A(n_4075),
.Y(n_6074)
);

AND2x4_ASAP7_75t_L g6075 ( 
.A(n_4233),
.B(n_4272),
.Y(n_6075)
);

AND2x4_ASAP7_75t_L g6076 ( 
.A(n_4272),
.B(n_4289),
.Y(n_6076)
);

AOI21xp5_ASAP7_75t_L g6077 ( 
.A1(n_4614),
.A2(n_4657),
.B(n_4642),
.Y(n_6077)
);

INVx2_ASAP7_75t_L g6078 ( 
.A(n_4657),
.Y(n_6078)
);

INVx1_ASAP7_75t_L g6079 ( 
.A(n_4662),
.Y(n_6079)
);

A2O1A1Ixp33_ASAP7_75t_L g6080 ( 
.A1(n_4218),
.A2(n_4293),
.B(n_4595),
.C(n_4291),
.Y(n_6080)
);

NAND2xp5_ASAP7_75t_SL g6081 ( 
.A(n_3508),
.B(n_3523),
.Y(n_6081)
);

CKINVDCx5p33_ASAP7_75t_R g6082 ( 
.A(n_4443),
.Y(n_6082)
);

O2A1O1Ixp33_ASAP7_75t_L g6083 ( 
.A1(n_4323),
.A2(n_4377),
.B(n_4387),
.C(n_4327),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_4662),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_4662),
.Y(n_6085)
);

INVx1_ASAP7_75t_SL g6086 ( 
.A(n_4009),
.Y(n_6086)
);

NOR2xp33_ASAP7_75t_L g6087 ( 
.A(n_3843),
.B(n_4026),
.Y(n_6087)
);

NOR2xp33_ASAP7_75t_L g6088 ( 
.A(n_4026),
.B(n_4124),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_4663),
.Y(n_6089)
);

NAND2xp5_ASAP7_75t_SL g6090 ( 
.A(n_3508),
.B(n_3523),
.Y(n_6090)
);

NAND2xp5_ASAP7_75t_L g6091 ( 
.A(n_3307),
.B(n_3312),
.Y(n_6091)
);

OAI21x1_ASAP7_75t_L g6092 ( 
.A1(n_4406),
.A2(n_4435),
.B(n_4430),
.Y(n_6092)
);

AND2x2_ASAP7_75t_L g6093 ( 
.A(n_4643),
.B(n_4663),
.Y(n_6093)
);

AOI21xp5_ASAP7_75t_L g6094 ( 
.A1(n_4663),
.A2(n_4681),
.B(n_4667),
.Y(n_6094)
);

OAI22x1_ASAP7_75t_L g6095 ( 
.A1(n_4667),
.A2(n_4703),
.B1(n_4705),
.B2(n_4681),
.Y(n_6095)
);

NAND2xp5_ASAP7_75t_L g6096 ( 
.A(n_3312),
.B(n_3331),
.Y(n_6096)
);

AOI21xp5_ASAP7_75t_L g6097 ( 
.A1(n_4667),
.A2(n_4703),
.B(n_4681),
.Y(n_6097)
);

NAND2xp5_ASAP7_75t_L g6098 ( 
.A(n_3331),
.B(n_3338),
.Y(n_6098)
);

AOI21xp5_ASAP7_75t_L g6099 ( 
.A1(n_4703),
.A2(n_4708),
.B(n_4705),
.Y(n_6099)
);

OA22x2_ASAP7_75t_L g6100 ( 
.A1(n_4289),
.A2(n_4355),
.B1(n_4376),
.B2(n_4316),
.Y(n_6100)
);

OAI21xp5_ASAP7_75t_L g6101 ( 
.A1(n_4377),
.A2(n_4588),
.B(n_4387),
.Y(n_6101)
);

NAND2xp5_ASAP7_75t_L g6102 ( 
.A(n_3338),
.B(n_3339),
.Y(n_6102)
);

AOI21xp5_ASAP7_75t_L g6103 ( 
.A1(n_4705),
.A2(n_4710),
.B(n_4708),
.Y(n_6103)
);

NAND2xp5_ASAP7_75t_L g6104 ( 
.A(n_3339),
.B(n_3343),
.Y(n_6104)
);

OAI22x1_ASAP7_75t_L g6105 ( 
.A1(n_4708),
.A2(n_4710),
.B1(n_4430),
.B2(n_4435),
.Y(n_6105)
);

NAND2xp5_ASAP7_75t_L g6106 ( 
.A(n_3343),
.B(n_3346),
.Y(n_6106)
);

INVx2_ASAP7_75t_SL g6107 ( 
.A(n_3241),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_4710),
.Y(n_6108)
);

BUFx8_ASAP7_75t_L g6109 ( 
.A(n_3494),
.Y(n_6109)
);

NAND2xp5_ASAP7_75t_SL g6110 ( 
.A(n_3508),
.B(n_3523),
.Y(n_6110)
);

AOI22xp5_ASAP7_75t_L g6111 ( 
.A1(n_3795),
.A2(n_3949),
.B1(n_4100),
.B2(n_4151),
.Y(n_6111)
);

BUFx6f_ASAP7_75t_L g6112 ( 
.A(n_3241),
.Y(n_6112)
);

NAND2xp5_ASAP7_75t_L g6113 ( 
.A(n_3346),
.B(n_3356),
.Y(n_6113)
);

OAI21xp5_ASAP7_75t_L g6114 ( 
.A1(n_4588),
.A2(n_4682),
.B(n_4619),
.Y(n_6114)
);

HB1xp67_ASAP7_75t_L g6115 ( 
.A(n_4009),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_3356),
.Y(n_6116)
);

AOI21xp5_ASAP7_75t_L g6117 ( 
.A1(n_4406),
.A2(n_4435),
.B(n_4430),
.Y(n_6117)
);

NAND2xp5_ASAP7_75t_L g6118 ( 
.A(n_3357),
.B(n_3374),
.Y(n_6118)
);

AOI21xp5_ASAP7_75t_L g6119 ( 
.A1(n_4406),
.A2(n_4435),
.B(n_4430),
.Y(n_6119)
);

AOI21xp5_ASAP7_75t_L g6120 ( 
.A1(n_4406),
.A2(n_4435),
.B(n_4430),
.Y(n_6120)
);

NAND2xp5_ASAP7_75t_SL g6121 ( 
.A(n_3523),
.B(n_3553),
.Y(n_6121)
);

INVx2_ASAP7_75t_L g6122 ( 
.A(n_4457),
.Y(n_6122)
);

AOI21x1_ASAP7_75t_L g6123 ( 
.A1(n_4619),
.A2(n_4684),
.B(n_4682),
.Y(n_6123)
);

NOR2x1_ASAP7_75t_L g6124 ( 
.A(n_3408),
.B(n_3442),
.Y(n_6124)
);

NOR2x1_ASAP7_75t_L g6125 ( 
.A(n_3408),
.B(n_3442),
.Y(n_6125)
);

OAI22xp5_ASAP7_75t_L g6126 ( 
.A1(n_3357),
.A2(n_3387),
.B1(n_3394),
.B2(n_3374),
.Y(n_6126)
);

AO21x1_ASAP7_75t_L g6127 ( 
.A1(n_3387),
.A2(n_3395),
.B(n_3394),
.Y(n_6127)
);

OAI321xp33_ASAP7_75t_L g6128 ( 
.A1(n_3395),
.A2(n_3841),
.A3(n_3746),
.B1(n_3768),
.B2(n_3740),
.C(n_3734),
.Y(n_6128)
);

AOI33xp33_ASAP7_75t_L g6129 ( 
.A1(n_4123),
.A2(n_4125),
.A3(n_4127),
.B1(n_4102),
.B2(n_3599),
.B3(n_3901),
.Y(n_6129)
);

OR2x2_ASAP7_75t_L g6130 ( 
.A(n_4025),
.B(n_3910),
.Y(n_6130)
);

INVx2_ASAP7_75t_L g6131 ( 
.A(n_4457),
.Y(n_6131)
);

NAND2xp5_ASAP7_75t_L g6132 ( 
.A(n_3400),
.B(n_3404),
.Y(n_6132)
);

NAND2xp5_ASAP7_75t_SL g6133 ( 
.A(n_3553),
.B(n_3653),
.Y(n_6133)
);

AOI22xp5_ASAP7_75t_L g6134 ( 
.A1(n_3949),
.A2(n_4100),
.B1(n_4151),
.B2(n_4128),
.Y(n_6134)
);

BUFx6f_ASAP7_75t_L g6135 ( 
.A(n_3241),
.Y(n_6135)
);

NAND2xp5_ASAP7_75t_L g6136 ( 
.A(n_3400),
.B(n_3404),
.Y(n_6136)
);

INVx4_ASAP7_75t_L g6137 ( 
.A(n_3408),
.Y(n_6137)
);

INVx4_ASAP7_75t_L g6138 ( 
.A(n_3408),
.Y(n_6138)
);

AOI21xp5_ASAP7_75t_L g6139 ( 
.A1(n_4457),
.A2(n_4548),
.B(n_4544),
.Y(n_6139)
);

OAI21xp5_ASAP7_75t_L g6140 ( 
.A1(n_4684),
.A2(n_4049),
.B(n_4289),
.Y(n_6140)
);

NAND2xp5_ASAP7_75t_SL g6141 ( 
.A(n_3553),
.B(n_3653),
.Y(n_6141)
);

OAI22xp5_ASAP7_75t_L g6142 ( 
.A1(n_3407),
.A2(n_3413),
.B1(n_3417),
.B2(n_3412),
.Y(n_6142)
);

AND2x2_ASAP7_75t_L g6143 ( 
.A(n_4643),
.B(n_4457),
.Y(n_6143)
);

AOI21xp5_ASAP7_75t_L g6144 ( 
.A1(n_4457),
.A2(n_4548),
.B(n_4544),
.Y(n_6144)
);

OAI21xp5_ASAP7_75t_L g6145 ( 
.A1(n_4049),
.A2(n_4316),
.B(n_4289),
.Y(n_6145)
);

AOI21xp5_ASAP7_75t_L g6146 ( 
.A1(n_4544),
.A2(n_4555),
.B(n_4548),
.Y(n_6146)
);

NAND2xp5_ASAP7_75t_L g6147 ( 
.A(n_3407),
.B(n_3412),
.Y(n_6147)
);

AOI21xp5_ASAP7_75t_L g6148 ( 
.A1(n_4544),
.A2(n_4555),
.B(n_4548),
.Y(n_6148)
);

HB1xp67_ASAP7_75t_L g6149 ( 
.A(n_4058),
.Y(n_6149)
);

O2A1O1Ixp33_ASAP7_75t_L g6150 ( 
.A1(n_3918),
.A2(n_3935),
.B(n_3933),
.C(n_4102),
.Y(n_6150)
);

NAND2x1_ASAP7_75t_L g6151 ( 
.A(n_4507),
.B(n_3277),
.Y(n_6151)
);

AOI21xp5_ASAP7_75t_L g6152 ( 
.A1(n_4544),
.A2(n_4555),
.B(n_4548),
.Y(n_6152)
);

AOI21xp5_ASAP7_75t_L g6153 ( 
.A1(n_4555),
.A2(n_4577),
.B(n_4557),
.Y(n_6153)
);

AOI21xp5_ASAP7_75t_L g6154 ( 
.A1(n_4555),
.A2(n_4577),
.B(n_4557),
.Y(n_6154)
);

AOI21x1_ASAP7_75t_L g6155 ( 
.A1(n_4316),
.A2(n_4376),
.B(n_4355),
.Y(n_6155)
);

AOI21xp5_ASAP7_75t_L g6156 ( 
.A1(n_4557),
.A2(n_4610),
.B(n_4577),
.Y(n_6156)
);

INVx2_ASAP7_75t_L g6157 ( 
.A(n_4557),
.Y(n_6157)
);

AOI21xp5_ASAP7_75t_L g6158 ( 
.A1(n_4557),
.A2(n_4610),
.B(n_4577),
.Y(n_6158)
);

OAI22xp5_ASAP7_75t_L g6159 ( 
.A1(n_3417),
.A2(n_3432),
.B1(n_3433),
.B2(n_3422),
.Y(n_6159)
);

HB1xp67_ASAP7_75t_L g6160 ( 
.A(n_4058),
.Y(n_6160)
);

A2O1A1Ixp33_ASAP7_75t_L g6161 ( 
.A1(n_4218),
.A2(n_4293),
.B(n_4595),
.C(n_4291),
.Y(n_6161)
);

OAI22xp5_ASAP7_75t_L g6162 ( 
.A1(n_3433),
.A2(n_3450),
.B1(n_3466),
.B2(n_3456),
.Y(n_6162)
);

NAND2xp5_ASAP7_75t_L g6163 ( 
.A(n_3456),
.B(n_3466),
.Y(n_6163)
);

NAND2xp5_ASAP7_75t_L g6164 ( 
.A(n_3470),
.B(n_3474),
.Y(n_6164)
);

INVx2_ASAP7_75t_L g6165 ( 
.A(n_4577),
.Y(n_6165)
);

AOI21xp5_ASAP7_75t_L g6166 ( 
.A1(n_4610),
.A2(n_4686),
.B(n_4666),
.Y(n_6166)
);

O2A1O1Ixp33_ASAP7_75t_L g6167 ( 
.A1(n_3935),
.A2(n_4086),
.B(n_3470),
.C(n_3491),
.Y(n_6167)
);

NAND2xp5_ASAP7_75t_L g6168 ( 
.A(n_3491),
.B(n_3492),
.Y(n_6168)
);

INVx3_ASAP7_75t_L g6169 ( 
.A(n_4610),
.Y(n_6169)
);

NAND2xp5_ASAP7_75t_L g6170 ( 
.A(n_3492),
.B(n_3506),
.Y(n_6170)
);

AOI221xp5_ASAP7_75t_L g6171 ( 
.A1(n_3506),
.A2(n_3701),
.B1(n_3901),
.B2(n_3885),
.C(n_3883),
.Y(n_6171)
);

NAND2xp5_ASAP7_75t_L g6172 ( 
.A(n_3509),
.B(n_3513),
.Y(n_6172)
);

NAND2xp5_ASAP7_75t_SL g6173 ( 
.A(n_3553),
.B(n_3653),
.Y(n_6173)
);

NAND2xp5_ASAP7_75t_L g6174 ( 
.A(n_3509),
.B(n_3513),
.Y(n_6174)
);

BUFx6f_ASAP7_75t_L g6175 ( 
.A(n_3239),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_3529),
.Y(n_6176)
);

A2O1A1Ixp33_ASAP7_75t_L g6177 ( 
.A1(n_4291),
.A2(n_4595),
.B(n_4293),
.C(n_3875),
.Y(n_6177)
);

NOR2xp33_ASAP7_75t_L g6178 ( 
.A(n_4026),
.B(n_4124),
.Y(n_6178)
);

O2A1O1Ixp5_ASAP7_75t_L g6179 ( 
.A1(n_4610),
.A2(n_4686),
.B(n_4689),
.C(n_4666),
.Y(n_6179)
);

AOI22xp5_ASAP7_75t_L g6180 ( 
.A1(n_4100),
.A2(n_4128),
.B1(n_4026),
.B2(n_3927),
.Y(n_6180)
);

NOR2xp33_ASAP7_75t_SL g6181 ( 
.A(n_3494),
.B(n_3503),
.Y(n_6181)
);

NAND2xp5_ASAP7_75t_SL g6182 ( 
.A(n_3553),
.B(n_3653),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_3529),
.Y(n_6183)
);

NAND2xp5_ASAP7_75t_SL g6184 ( 
.A(n_3653),
.B(n_3871),
.Y(n_6184)
);

INVx2_ASAP7_75t_L g6185 ( 
.A(n_4666),
.Y(n_6185)
);

INVx2_ASAP7_75t_L g6186 ( 
.A(n_4666),
.Y(n_6186)
);

NOR3xp33_ASAP7_75t_L g6187 ( 
.A(n_4132),
.B(n_4137),
.C(n_4082),
.Y(n_6187)
);

AOI21xp5_ASAP7_75t_L g6188 ( 
.A1(n_4666),
.A2(n_4689),
.B(n_4686),
.Y(n_6188)
);

AOI21xp5_ASAP7_75t_L g6189 ( 
.A1(n_4692),
.A2(n_4693),
.B(n_3327),
.Y(n_6189)
);

NAND2xp5_ASAP7_75t_L g6190 ( 
.A(n_3535),
.B(n_3547),
.Y(n_6190)
);

AOI21xp5_ASAP7_75t_L g6191 ( 
.A1(n_4692),
.A2(n_4693),
.B(n_3327),
.Y(n_6191)
);

A2O1A1Ixp33_ASAP7_75t_L g6192 ( 
.A1(n_3871),
.A2(n_3875),
.B(n_4086),
.C(n_4132),
.Y(n_6192)
);

NAND2xp5_ASAP7_75t_L g6193 ( 
.A(n_3535),
.B(n_3547),
.Y(n_6193)
);

OAI22x1_ASAP7_75t_L g6194 ( 
.A1(n_4692),
.A2(n_4693),
.B1(n_3563),
.B2(n_3578),
.Y(n_6194)
);

AOI21xp5_ASAP7_75t_L g6195 ( 
.A1(n_4693),
.A2(n_3277),
.B(n_3910),
.Y(n_6195)
);

BUFx12f_ASAP7_75t_L g6196 ( 
.A(n_3494),
.Y(n_6196)
);

NAND2xp5_ASAP7_75t_L g6197 ( 
.A(n_3563),
.B(n_3576),
.Y(n_6197)
);

NOR2xp33_ASAP7_75t_L g6198 ( 
.A(n_4026),
.B(n_4149),
.Y(n_6198)
);

AOI21xp5_ASAP7_75t_L g6199 ( 
.A1(n_3910),
.A2(n_3934),
.B(n_3930),
.Y(n_6199)
);

AOI21xp5_ASAP7_75t_L g6200 ( 
.A1(n_3930),
.A2(n_3945),
.B(n_3934),
.Y(n_6200)
);

INVx5_ASAP7_75t_L g6201 ( 
.A(n_4507),
.Y(n_6201)
);

AND2x2_ASAP7_75t_L g6202 ( 
.A(n_4643),
.B(n_4025),
.Y(n_6202)
);

NAND2xp5_ASAP7_75t_L g6203 ( 
.A(n_3576),
.B(n_3578),
.Y(n_6203)
);

AOI21xp5_ASAP7_75t_L g6204 ( 
.A1(n_3930),
.A2(n_3945),
.B(n_3934),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_3582),
.Y(n_6205)
);

NOR2x1_ASAP7_75t_L g6206 ( 
.A(n_3442),
.B(n_3446),
.Y(n_6206)
);

A2O1A1Ixp33_ASAP7_75t_L g6207 ( 
.A1(n_3871),
.A2(n_3875),
.B(n_4137),
.C(n_4132),
.Y(n_6207)
);

NAND2xp5_ASAP7_75t_L g6208 ( 
.A(n_3582),
.B(n_3594),
.Y(n_6208)
);

OAI21xp5_ASAP7_75t_L g6209 ( 
.A1(n_4316),
.A2(n_4376),
.B(n_4355),
.Y(n_6209)
);

OAI321xp33_ASAP7_75t_L g6210 ( 
.A1(n_3594),
.A2(n_3746),
.A3(n_3740),
.B1(n_3885),
.B2(n_3883),
.C(n_3881),
.Y(n_6210)
);

NAND2xp5_ASAP7_75t_L g6211 ( 
.A(n_3595),
.B(n_3599),
.Y(n_6211)
);

INVx2_ASAP7_75t_SL g6212 ( 
.A(n_3239),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_3595),
.Y(n_6213)
);

INVx3_ASAP7_75t_SL g6214 ( 
.A(n_4104),
.Y(n_6214)
);

AOI21xp5_ASAP7_75t_L g6215 ( 
.A1(n_3945),
.A2(n_3948),
.B(n_4025),
.Y(n_6215)
);

NAND2xp5_ASAP7_75t_L g6216 ( 
.A(n_3610),
.B(n_3611),
.Y(n_6216)
);

NAND2xp5_ASAP7_75t_L g6217 ( 
.A(n_3610),
.B(n_3611),
.Y(n_6217)
);

BUFx2_ASAP7_75t_L g6218 ( 
.A(n_4507),
.Y(n_6218)
);

AOI21xp5_ASAP7_75t_L g6219 ( 
.A1(n_3948),
.A2(n_3620),
.B(n_3615),
.Y(n_6219)
);

INVx1_ASAP7_75t_L g6220 ( 
.A(n_3615),
.Y(n_6220)
);

NOR2xp33_ASAP7_75t_L g6221 ( 
.A(n_4082),
.B(n_4455),
.Y(n_6221)
);

HB1xp67_ASAP7_75t_L g6222 ( 
.A(n_4058),
.Y(n_6222)
);

BUFx8_ASAP7_75t_L g6223 ( 
.A(n_3503),
.Y(n_6223)
);

OAI22xp5_ASAP7_75t_SL g6224 ( 
.A1(n_3832),
.A2(n_4114),
.B1(n_3503),
.B2(n_4094),
.Y(n_6224)
);

AOI21xp5_ASAP7_75t_L g6225 ( 
.A1(n_3948),
.A2(n_3630),
.B(n_3620),
.Y(n_6225)
);

AOI22xp33_ASAP7_75t_L g6226 ( 
.A1(n_4355),
.A2(n_4571),
.B1(n_4459),
.B2(n_4448),
.Y(n_6226)
);

BUFx6f_ASAP7_75t_L g6227 ( 
.A(n_3239),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_SL g6228 ( 
.A(n_3968),
.B(n_3972),
.Y(n_6228)
);

AOI22xp5_ASAP7_75t_L g6229 ( 
.A1(n_4128),
.A2(n_3927),
.B1(n_4132),
.B2(n_4137),
.Y(n_6229)
);

O2A1O1Ixp33_ASAP7_75t_L g6230 ( 
.A1(n_3636),
.A2(n_3881),
.B(n_3873),
.C(n_3865),
.Y(n_6230)
);

BUFx2_ASAP7_75t_L g6231 ( 
.A(n_4507),
.Y(n_6231)
);

BUFx2_ASAP7_75t_L g6232 ( 
.A(n_4507),
.Y(n_6232)
);

NOR2xp33_ASAP7_75t_L g6233 ( 
.A(n_4469),
.B(n_4655),
.Y(n_6233)
);

INVxp67_ASAP7_75t_L g6234 ( 
.A(n_3636),
.Y(n_6234)
);

CKINVDCx14_ASAP7_75t_R g6235 ( 
.A(n_3832),
.Y(n_6235)
);

INVx1_ASAP7_75t_SL g6236 ( 
.A(n_3608),
.Y(n_6236)
);

NOR2xp33_ASAP7_75t_L g6237 ( 
.A(n_4664),
.B(n_3802),
.Y(n_6237)
);

INVx1_ASAP7_75t_L g6238 ( 
.A(n_3642),
.Y(n_6238)
);

AOI21xp5_ASAP7_75t_L g6239 ( 
.A1(n_3642),
.A2(n_3656),
.B(n_3648),
.Y(n_6239)
);

NAND2xp5_ASAP7_75t_L g6240 ( 
.A(n_3648),
.B(n_3656),
.Y(n_6240)
);

NOR2xp33_ASAP7_75t_L g6241 ( 
.A(n_4125),
.B(n_4132),
.Y(n_6241)
);

NAND2xp5_ASAP7_75t_SL g6242 ( 
.A(n_3968),
.B(n_3972),
.Y(n_6242)
);

OAI21xp5_ASAP7_75t_L g6243 ( 
.A1(n_4355),
.A2(n_4448),
.B(n_4376),
.Y(n_6243)
);

AOI21xp5_ASAP7_75t_L g6244 ( 
.A1(n_3664),
.A2(n_3671),
.B(n_3670),
.Y(n_6244)
);

NAND2xp5_ASAP7_75t_L g6245 ( 
.A(n_3664),
.B(n_3670),
.Y(n_6245)
);

NAND2xp5_ASAP7_75t_L g6246 ( 
.A(n_3671),
.B(n_3674),
.Y(n_6246)
);

NOR2xp33_ASAP7_75t_L g6247 ( 
.A(n_4137),
.B(n_4128),
.Y(n_6247)
);

A2O1A1Ixp33_ASAP7_75t_L g6248 ( 
.A1(n_4137),
.A2(n_3679),
.B(n_3773),
.C(n_3769),
.Y(n_6248)
);

O2A1O1Ixp33_ASAP7_75t_L g6249 ( 
.A1(n_3674),
.A2(n_3842),
.B(n_3722),
.C(n_3729),
.Y(n_6249)
);

NAND2xp5_ASAP7_75t_L g6250 ( 
.A(n_3675),
.B(n_3679),
.Y(n_6250)
);

AOI221xp5_ASAP7_75t_L g6251 ( 
.A1(n_3675),
.A2(n_3808),
.B1(n_3722),
.B2(n_3729),
.C(n_3873),
.Y(n_6251)
);

NAND2xp5_ASAP7_75t_L g6252 ( 
.A(n_3680),
.B(n_3700),
.Y(n_6252)
);

NAND2xp5_ASAP7_75t_L g6253 ( 
.A(n_3700),
.B(n_3701),
.Y(n_6253)
);

AOI21x1_ASAP7_75t_L g6254 ( 
.A1(n_5218),
.A2(n_3769),
.B(n_3757),
.Y(n_6254)
);

HB1xp67_ASAP7_75t_L g6255 ( 
.A(n_5687),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_6127),
.Y(n_6256)
);

AOI21xp5_ASAP7_75t_L g6257 ( 
.A1(n_4727),
.A2(n_3773),
.B(n_3757),
.Y(n_6257)
);

AND2x4_ASAP7_75t_L g6258 ( 
.A(n_4749),
.B(n_4797),
.Y(n_6258)
);

BUFx6f_ASAP7_75t_L g6259 ( 
.A(n_4758),
.Y(n_6259)
);

OAI21x1_ASAP7_75t_L g6260 ( 
.A1(n_4727),
.A2(n_3799),
.B(n_3824),
.Y(n_6260)
);

OAI21x1_ASAP7_75t_L g6261 ( 
.A1(n_4731),
.A2(n_3799),
.B(n_3790),
.Y(n_6261)
);

AO31x2_ASAP7_75t_L g6262 ( 
.A1(n_5280),
.A2(n_3808),
.A3(n_3803),
.B(n_3809),
.Y(n_6262)
);

NAND2xp5_ASAP7_75t_L g6263 ( 
.A(n_4958),
.B(n_3803),
.Y(n_6263)
);

NAND2xp5_ASAP7_75t_L g6264 ( 
.A(n_4958),
.B(n_3809),
.Y(n_6264)
);

AOI21x1_ASAP7_75t_L g6265 ( 
.A1(n_5218),
.A2(n_5260),
.B(n_5233),
.Y(n_6265)
);

BUFx2_ASAP7_75t_L g6266 ( 
.A(n_5478),
.Y(n_6266)
);

AOI21xp5_ASAP7_75t_L g6267 ( 
.A1(n_4731),
.A2(n_3810),
.B(n_4303),
.Y(n_6267)
);

AOI21xp5_ASAP7_75t_L g6268 ( 
.A1(n_4748),
.A2(n_3810),
.B(n_4303),
.Y(n_6268)
);

CKINVDCx5p33_ASAP7_75t_R g6269 ( 
.A(n_5011),
.Y(n_6269)
);

AO21x1_ASAP7_75t_L g6270 ( 
.A1(n_5272),
.A2(n_4453),
.B(n_4454),
.Y(n_6270)
);

AOI221xp5_ASAP7_75t_SL g6271 ( 
.A1(n_4785),
.A2(n_3239),
.B1(n_4040),
.B2(n_4027),
.C(n_4069),
.Y(n_6271)
);

AO31x2_ASAP7_75t_L g6272 ( 
.A1(n_5280),
.A2(n_4027),
.A3(n_4040),
.B(n_4069),
.Y(n_6272)
);

NOR2x1_ASAP7_75t_SL g6273 ( 
.A(n_5291),
.B(n_3239),
.Y(n_6273)
);

INVx3_ASAP7_75t_L g6274 ( 
.A(n_5975),
.Y(n_6274)
);

A2O1A1Ixp33_ASAP7_75t_L g6275 ( 
.A1(n_4793),
.A2(n_3446),
.B(n_3442),
.C(n_4133),
.Y(n_6275)
);

O2A1O1Ixp5_ASAP7_75t_L g6276 ( 
.A1(n_4852),
.A2(n_4855),
.B(n_4953),
.C(n_4900),
.Y(n_6276)
);

O2A1O1Ixp33_ASAP7_75t_L g6277 ( 
.A1(n_4738),
.A2(n_4115),
.B(n_4347),
.C(n_4637),
.Y(n_6277)
);

OAI21x1_ASAP7_75t_L g6278 ( 
.A1(n_4750),
.A2(n_4011),
.B(n_4039),
.Y(n_6278)
);

NAND2xp5_ASAP7_75t_L g6279 ( 
.A(n_4963),
.B(n_3239),
.Y(n_6279)
);

NAND2xp5_ASAP7_75t_L g6280 ( 
.A(n_4963),
.B(n_3239),
.Y(n_6280)
);

OAI21xp5_ASAP7_75t_L g6281 ( 
.A1(n_4807),
.A2(n_4453),
.B(n_4639),
.Y(n_6281)
);

INVx1_ASAP7_75t_L g6282 ( 
.A(n_6127),
.Y(n_6282)
);

CKINVDCx5p33_ASAP7_75t_R g6283 ( 
.A(n_4853),
.Y(n_6283)
);

AND2x4_ASAP7_75t_L g6284 ( 
.A(n_4749),
.B(n_4376),
.Y(n_6284)
);

A2O1A1Ixp33_ASAP7_75t_L g6285 ( 
.A1(n_4793),
.A2(n_3446),
.B(n_3442),
.C(n_3743),
.Y(n_6285)
);

NAND3xp33_ASAP7_75t_SL g6286 ( 
.A(n_4766),
.B(n_3923),
.C(n_4114),
.Y(n_6286)
);

INVx2_ASAP7_75t_SL g6287 ( 
.A(n_5439),
.Y(n_6287)
);

BUFx10_ASAP7_75t_L g6288 ( 
.A(n_5276),
.Y(n_6288)
);

O2A1O1Ixp5_ASAP7_75t_L g6289 ( 
.A1(n_4852),
.A2(n_4448),
.B(n_4460),
.C(n_4459),
.Y(n_6289)
);

INVx1_ASAP7_75t_L g6290 ( 
.A(n_5816),
.Y(n_6290)
);

INVx4_ASAP7_75t_L g6291 ( 
.A(n_5254),
.Y(n_6291)
);

BUFx6f_ASAP7_75t_SL g6292 ( 
.A(n_4758),
.Y(n_6292)
);

OAI21x1_ASAP7_75t_L g6293 ( 
.A1(n_5106),
.A2(n_4011),
.B(n_4039),
.Y(n_6293)
);

NAND2xp5_ASAP7_75t_L g6294 ( 
.A(n_4978),
.B(n_3239),
.Y(n_6294)
);

AO31x2_ASAP7_75t_L g6295 ( 
.A1(n_6194),
.A2(n_4027),
.A3(n_4040),
.B(n_3972),
.Y(n_6295)
);

OAI21x1_ASAP7_75t_L g6296 ( 
.A1(n_5109),
.A2(n_4011),
.B(n_4039),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_5816),
.Y(n_6297)
);

OAI21xp5_ASAP7_75t_L g6298 ( 
.A1(n_4807),
.A2(n_4459),
.B(n_4639),
.Y(n_6298)
);

OAI21x1_ASAP7_75t_L g6299 ( 
.A1(n_5109),
.A2(n_4011),
.B(n_4039),
.Y(n_6299)
);

AND2x2_ASAP7_75t_L g6300 ( 
.A(n_5677),
.B(n_5716),
.Y(n_6300)
);

AND3x2_ASAP7_75t_L g6301 ( 
.A(n_4786),
.B(n_4128),
.C(n_4460),
.Y(n_6301)
);

HB1xp67_ASAP7_75t_L g6302 ( 
.A(n_5687),
.Y(n_6302)
);

AO21x2_ASAP7_75t_L g6303 ( 
.A1(n_4868),
.A2(n_4459),
.B(n_4448),
.Y(n_6303)
);

OAI21xp5_ASAP7_75t_L g6304 ( 
.A1(n_4786),
.A2(n_4827),
.B(n_4769),
.Y(n_6304)
);

AOI21xp5_ASAP7_75t_L g6305 ( 
.A1(n_4778),
.A2(n_3237),
.B(n_4337),
.Y(n_6305)
);

AOI21xp5_ASAP7_75t_L g6306 ( 
.A1(n_4778),
.A2(n_3237),
.B(n_4337),
.Y(n_6306)
);

INVx1_ASAP7_75t_L g6307 ( 
.A(n_5816),
.Y(n_6307)
);

NAND2xp5_ASAP7_75t_SL g6308 ( 
.A(n_4806),
.B(n_4011),
.Y(n_6308)
);

BUFx3_ASAP7_75t_L g6309 ( 
.A(n_5359),
.Y(n_6309)
);

BUFx3_ASAP7_75t_L g6310 ( 
.A(n_5359),
.Y(n_6310)
);

AOI21xp5_ASAP7_75t_L g6311 ( 
.A1(n_4789),
.A2(n_4347),
.B(n_4337),
.Y(n_6311)
);

INVx4_ASAP7_75t_L g6312 ( 
.A(n_5254),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_5816),
.Y(n_6313)
);

NAND2xp5_ASAP7_75t_L g6314 ( 
.A(n_4978),
.B(n_4507),
.Y(n_6314)
);

AOI221x1_ASAP7_75t_L g6315 ( 
.A1(n_4988),
.A2(n_4639),
.B1(n_4571),
.B2(n_4448),
.C(n_4514),
.Y(n_6315)
);

NAND2xp5_ASAP7_75t_L g6316 ( 
.A(n_4983),
.B(n_4507),
.Y(n_6316)
);

BUFx10_ASAP7_75t_L g6317 ( 
.A(n_5276),
.Y(n_6317)
);

AOI21xp5_ASAP7_75t_L g6318 ( 
.A1(n_4789),
.A2(n_4329),
.B(n_4307),
.Y(n_6318)
);

AOI21xp5_ASAP7_75t_L g6319 ( 
.A1(n_4759),
.A2(n_4329),
.B(n_4307),
.Y(n_6319)
);

INVx2_ASAP7_75t_L g6320 ( 
.A(n_5233),
.Y(n_6320)
);

OAI22x1_ASAP7_75t_L g6321 ( 
.A1(n_4925),
.A2(n_4639),
.B1(n_4453),
.B2(n_4454),
.Y(n_6321)
);

INVx2_ASAP7_75t_L g6322 ( 
.A(n_5260),
.Y(n_6322)
);

NAND2xp5_ASAP7_75t_L g6323 ( 
.A(n_4983),
.B(n_4507),
.Y(n_6323)
);

INVx4_ASAP7_75t_L g6324 ( 
.A(n_5254),
.Y(n_6324)
);

OAI21x1_ASAP7_75t_L g6325 ( 
.A1(n_5209),
.A2(n_4041),
.B(n_4052),
.Y(n_6325)
);

INVx1_ASAP7_75t_L g6326 ( 
.A(n_5287),
.Y(n_6326)
);

NAND3xp33_ASAP7_75t_L g6327 ( 
.A(n_4766),
.B(n_4454),
.C(n_4571),
.Y(n_6327)
);

AOI21xp5_ASAP7_75t_L g6328 ( 
.A1(n_4759),
.A2(n_4329),
.B(n_4307),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_5287),
.Y(n_6329)
);

NOR2x1_ASAP7_75t_L g6330 ( 
.A(n_4817),
.B(n_3446),
.Y(n_6330)
);

NAND2xp5_ASAP7_75t_L g6331 ( 
.A(n_4987),
.B(n_4507),
.Y(n_6331)
);

AOI21xp5_ASAP7_75t_L g6332 ( 
.A1(n_4772),
.A2(n_4277),
.B(n_4303),
.Y(n_6332)
);

AOI21xp5_ASAP7_75t_L g6333 ( 
.A1(n_4772),
.A2(n_4277),
.B(n_4231),
.Y(n_6333)
);

AOI21xp5_ASAP7_75t_L g6334 ( 
.A1(n_4893),
.A2(n_4277),
.B(n_4231),
.Y(n_6334)
);

INVxp67_ASAP7_75t_L g6335 ( 
.A(n_5625),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_SL g6336 ( 
.A(n_4806),
.B(n_4453),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_5318),
.Y(n_6337)
);

AND2x2_ASAP7_75t_L g6338 ( 
.A(n_5677),
.B(n_4453),
.Y(n_6338)
);

NAND2xp5_ASAP7_75t_L g6339 ( 
.A(n_4987),
.B(n_4454),
.Y(n_6339)
);

INVx1_ASAP7_75t_SL g6340 ( 
.A(n_4725),
.Y(n_6340)
);

OAI21x1_ASAP7_75t_L g6341 ( 
.A1(n_5210),
.A2(n_4041),
.B(n_4052),
.Y(n_6341)
);

NOR2xp33_ASAP7_75t_L g6342 ( 
.A(n_4799),
.B(n_4454),
.Y(n_6342)
);

OAI21x1_ASAP7_75t_L g6343 ( 
.A1(n_5213),
.A2(n_4041),
.B(n_4052),
.Y(n_6343)
);

AOI21x1_ASAP7_75t_SL g6344 ( 
.A1(n_5091),
.A2(n_4639),
.B(n_4571),
.Y(n_6344)
);

AOI21x1_ASAP7_75t_L g6345 ( 
.A1(n_5318),
.A2(n_4459),
.B(n_4460),
.Y(n_6345)
);

AOI21xp5_ASAP7_75t_L g6346 ( 
.A1(n_4893),
.A2(n_4199),
.B(n_4205),
.Y(n_6346)
);

NOR2xp33_ASAP7_75t_L g6347 ( 
.A(n_4799),
.B(n_4460),
.Y(n_6347)
);

INVx2_ASAP7_75t_L g6348 ( 
.A(n_5319),
.Y(n_6348)
);

AOI22xp5_ASAP7_75t_L g6349 ( 
.A1(n_4925),
.A2(n_4571),
.B1(n_4514),
.B2(n_4460),
.Y(n_6349)
);

OAI21x1_ASAP7_75t_L g6350 ( 
.A1(n_5213),
.A2(n_5230),
.B(n_5221),
.Y(n_6350)
);

AOI21xp5_ASAP7_75t_L g6351 ( 
.A1(n_4776),
.A2(n_4777),
.B(n_4879),
.Y(n_6351)
);

NAND2xp5_ASAP7_75t_L g6352 ( 
.A(n_4991),
.B(n_4993),
.Y(n_6352)
);

OAI21x1_ASAP7_75t_L g6353 ( 
.A1(n_5221),
.A2(n_4052),
.B(n_3446),
.Y(n_6353)
);

NAND2xp5_ASAP7_75t_L g6354 ( 
.A(n_4991),
.B(n_4514),
.Y(n_6354)
);

CKINVDCx8_ASAP7_75t_R g6355 ( 
.A(n_6201),
.Y(n_6355)
);

INVx1_ASAP7_75t_SL g6356 ( 
.A(n_4725),
.Y(n_6356)
);

AO21x2_ASAP7_75t_L g6357 ( 
.A1(n_4868),
.A2(n_4514),
.B(n_4067),
.Y(n_6357)
);

AOI21xp5_ASAP7_75t_L g6358 ( 
.A1(n_4776),
.A2(n_4396),
.B(n_4516),
.Y(n_6358)
);

OAI21x1_ASAP7_75t_L g6359 ( 
.A1(n_5230),
.A2(n_5232),
.B(n_5231),
.Y(n_6359)
);

A2O1A1Ixp33_ASAP7_75t_L g6360 ( 
.A1(n_4740),
.A2(n_3673),
.B(n_3443),
.C(n_3454),
.Y(n_6360)
);

AOI21xp5_ASAP7_75t_L g6361 ( 
.A1(n_4777),
.A2(n_4396),
.B(n_4516),
.Y(n_6361)
);

A2O1A1Ixp33_ASAP7_75t_L g6362 ( 
.A1(n_4740),
.A2(n_3673),
.B(n_3443),
.C(n_3454),
.Y(n_6362)
);

AOI21xp5_ASAP7_75t_L g6363 ( 
.A1(n_4879),
.A2(n_4396),
.B(n_4516),
.Y(n_6363)
);

OAI21xp5_ASAP7_75t_L g6364 ( 
.A1(n_4830),
.A2(n_4833),
.B(n_4754),
.Y(n_6364)
);

OAI21x1_ASAP7_75t_L g6365 ( 
.A1(n_5231),
.A2(n_3923),
.B(n_4071),
.Y(n_6365)
);

INVx2_ASAP7_75t_L g6366 ( 
.A(n_5319),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_5430),
.Y(n_6367)
);

NAND2xp33_ASAP7_75t_L g6368 ( 
.A(n_4988),
.B(n_3877),
.Y(n_6368)
);

AOI21xp33_ASAP7_75t_L g6369 ( 
.A1(n_4742),
.A2(n_4225),
.B(n_4637),
.Y(n_6369)
);

NOR2xp33_ASAP7_75t_L g6370 ( 
.A(n_4785),
.B(n_4514),
.Y(n_6370)
);

AOI21xp5_ASAP7_75t_L g6371 ( 
.A1(n_4890),
.A2(n_4225),
.B(n_4635),
.Y(n_6371)
);

AND2x4_ASAP7_75t_L g6372 ( 
.A(n_4749),
.B(n_4199),
.Y(n_6372)
);

AOI21xp5_ASAP7_75t_L g6373 ( 
.A1(n_4890),
.A2(n_4225),
.B(n_4635),
.Y(n_6373)
);

OAI21xp5_ASAP7_75t_L g6374 ( 
.A1(n_4754),
.A2(n_4637),
.B(n_4347),
.Y(n_6374)
);

NAND2xp5_ASAP7_75t_L g6375 ( 
.A(n_4993),
.B(n_4199),
.Y(n_6375)
);

AOI21x1_ASAP7_75t_L g6376 ( 
.A1(n_5430),
.A2(n_4392),
.B(n_4635),
.Y(n_6376)
);

OAI21x1_ASAP7_75t_L g6377 ( 
.A1(n_5232),
.A2(n_3923),
.B(n_4071),
.Y(n_6377)
);

NAND2xp5_ASAP7_75t_L g6378 ( 
.A(n_4994),
.B(n_4205),
.Y(n_6378)
);

INVx1_ASAP7_75t_L g6379 ( 
.A(n_5482),
.Y(n_6379)
);

AO21x1_ASAP7_75t_L g6380 ( 
.A1(n_5272),
.A2(n_3972),
.B(n_3923),
.Y(n_6380)
);

NAND2xp5_ASAP7_75t_L g6381 ( 
.A(n_4994),
.B(n_4205),
.Y(n_6381)
);

AOI21x1_ASAP7_75t_L g6382 ( 
.A1(n_5482),
.A2(n_4392),
.B(n_4601),
.Y(n_6382)
);

AOI22xp5_ASAP7_75t_L g6383 ( 
.A1(n_4755),
.A2(n_3942),
.B1(n_4421),
.B2(n_4392),
.Y(n_6383)
);

INVx2_ASAP7_75t_SL g6384 ( 
.A(n_5439),
.Y(n_6384)
);

AO21x1_ASAP7_75t_L g6385 ( 
.A1(n_5288),
.A2(n_3972),
.B(n_4067),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_L g6386 ( 
.A(n_5005),
.B(n_4231),
.Y(n_6386)
);

AND2x4_ASAP7_75t_L g6387 ( 
.A(n_4749),
.B(n_4421),
.Y(n_6387)
);

BUFx6f_ASAP7_75t_L g6388 ( 
.A(n_4758),
.Y(n_6388)
);

AOI21xp33_ASAP7_75t_L g6389 ( 
.A1(n_4742),
.A2(n_4601),
.B(n_4421),
.Y(n_6389)
);

A2O1A1Ixp33_ASAP7_75t_L g6390 ( 
.A1(n_4751),
.A2(n_3846),
.B(n_3443),
.C(n_3454),
.Y(n_6390)
);

NAND2xp5_ASAP7_75t_L g6391 ( 
.A(n_5005),
.B(n_5014),
.Y(n_6391)
);

NOR2x1_ASAP7_75t_L g6392 ( 
.A(n_4817),
.B(n_4108),
.Y(n_6392)
);

INVx1_ASAP7_75t_L g6393 ( 
.A(n_5508),
.Y(n_6393)
);

AOI21xp5_ASAP7_75t_L g6394 ( 
.A1(n_4892),
.A2(n_4601),
.B(n_3942),
.Y(n_6394)
);

AOI21xp5_ASAP7_75t_L g6395 ( 
.A1(n_4892),
.A2(n_3942),
.B(n_4019),
.Y(n_6395)
);

INVx1_ASAP7_75t_SL g6396 ( 
.A(n_4911),
.Y(n_6396)
);

OR2x2_ASAP7_75t_L g6397 ( 
.A(n_4857),
.B(n_4083),
.Y(n_6397)
);

OAI21x1_ASAP7_75t_L g6398 ( 
.A1(n_5238),
.A2(n_4071),
.B(n_3725),
.Y(n_6398)
);

INVx3_ASAP7_75t_L g6399 ( 
.A(n_5975),
.Y(n_6399)
);

AOI21xp5_ASAP7_75t_L g6400 ( 
.A1(n_4798),
.A2(n_3942),
.B(n_4019),
.Y(n_6400)
);

NAND2xp5_ASAP7_75t_L g6401 ( 
.A(n_5014),
.B(n_5020),
.Y(n_6401)
);

OAI21xp33_ASAP7_75t_SL g6402 ( 
.A1(n_4995),
.A2(n_3942),
.B(n_3891),
.Y(n_6402)
);

OAI21xp5_ASAP7_75t_L g6403 ( 
.A1(n_4814),
.A2(n_4083),
.B(n_4115),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_5508),
.Y(n_6404)
);

OR2x2_ASAP7_75t_L g6405 ( 
.A(n_4857),
.B(n_4083),
.Y(n_6405)
);

NAND2xp5_ASAP7_75t_L g6406 ( 
.A(n_5020),
.B(n_4019),
.Y(n_6406)
);

INVxp67_ASAP7_75t_L g6407 ( 
.A(n_5971),
.Y(n_6407)
);

AO21x2_ASAP7_75t_L g6408 ( 
.A1(n_4870),
.A2(n_4097),
.B(n_4716),
.Y(n_6408)
);

AOI21xp5_ASAP7_75t_L g6409 ( 
.A1(n_4798),
.A2(n_3942),
.B(n_4019),
.Y(n_6409)
);

BUFx2_ASAP7_75t_L g6410 ( 
.A(n_5478),
.Y(n_6410)
);

AO31x2_ASAP7_75t_L g6411 ( 
.A1(n_6194),
.A2(n_4870),
.A3(n_4900),
.B(n_4855),
.Y(n_6411)
);

OAI21x1_ASAP7_75t_L g6412 ( 
.A1(n_5238),
.A2(n_4071),
.B(n_3685),
.Y(n_6412)
);

OAI21x1_ASAP7_75t_L g6413 ( 
.A1(n_5239),
.A2(n_4071),
.B(n_3685),
.Y(n_6413)
);

OAI21x1_ASAP7_75t_L g6414 ( 
.A1(n_5239),
.A2(n_3827),
.B(n_3711),
.Y(n_6414)
);

NAND2xp5_ASAP7_75t_L g6415 ( 
.A(n_5024),
.B(n_4019),
.Y(n_6415)
);

INVxp67_ASAP7_75t_SL g6416 ( 
.A(n_5923),
.Y(n_6416)
);

NOR2xp67_ASAP7_75t_SL g6417 ( 
.A(n_5121),
.B(n_3968),
.Y(n_6417)
);

NOR2xp33_ASAP7_75t_L g6418 ( 
.A(n_4726),
.B(n_3526),
.Y(n_6418)
);

INVx4_ASAP7_75t_L g6419 ( 
.A(n_5254),
.Y(n_6419)
);

OAI21x1_ASAP7_75t_L g6420 ( 
.A1(n_5257),
.A2(n_3827),
.B(n_3711),
.Y(n_6420)
);

OAI22xp5_ASAP7_75t_L g6421 ( 
.A1(n_4972),
.A2(n_4077),
.B1(n_3868),
.B2(n_3862),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_5547),
.Y(n_6422)
);

NAND2xp5_ASAP7_75t_L g6423 ( 
.A(n_5024),
.B(n_4019),
.Y(n_6423)
);

AOI21x1_ASAP7_75t_L g6424 ( 
.A1(n_5547),
.A2(n_3942),
.B(n_3891),
.Y(n_6424)
);

NOR2xp67_ASAP7_75t_L g6425 ( 
.A(n_5065),
.B(n_3968),
.Y(n_6425)
);

INVx4_ASAP7_75t_L g6426 ( 
.A(n_5254),
.Y(n_6426)
);

OAI21xp5_ASAP7_75t_L g6427 ( 
.A1(n_4814),
.A2(n_3968),
.B(n_4087),
.Y(n_6427)
);

NAND2xp5_ASAP7_75t_L g6428 ( 
.A(n_5031),
.B(n_4019),
.Y(n_6428)
);

INVxp67_ASAP7_75t_L g6429 ( 
.A(n_6074),
.Y(n_6429)
);

INVx2_ASAP7_75t_L g6430 ( 
.A(n_5560),
.Y(n_6430)
);

NAND2xp5_ASAP7_75t_SL g6431 ( 
.A(n_4992),
.B(n_3968),
.Y(n_6431)
);

OAI21x1_ASAP7_75t_L g6432 ( 
.A1(n_5257),
.A2(n_3827),
.B(n_3711),
.Y(n_6432)
);

HB1xp67_ASAP7_75t_L g6433 ( 
.A(n_5747),
.Y(n_6433)
);

AO21x1_ASAP7_75t_L g6434 ( 
.A1(n_5288),
.A2(n_3900),
.B(n_3747),
.Y(n_6434)
);

AOI21x1_ASAP7_75t_L g6435 ( 
.A1(n_5560),
.A2(n_3891),
.B(n_4108),
.Y(n_6435)
);

NAND2xp5_ASAP7_75t_L g6436 ( 
.A(n_5031),
.B(n_5071),
.Y(n_6436)
);

OAI21x1_ASAP7_75t_L g6437 ( 
.A1(n_5258),
.A2(n_5263),
.B(n_5262),
.Y(n_6437)
);

OR2x2_ASAP7_75t_L g6438 ( 
.A(n_5379),
.B(n_5404),
.Y(n_6438)
);

AND3x4_ASAP7_75t_L g6439 ( 
.A(n_4992),
.B(n_3868),
.C(n_3862),
.Y(n_6439)
);

AO31x2_ASAP7_75t_L g6440 ( 
.A1(n_6194),
.A2(n_3900),
.A3(n_3747),
.B(n_3526),
.Y(n_6440)
);

OAI22xp5_ASAP7_75t_L g6441 ( 
.A1(n_4972),
.A2(n_4077),
.B1(n_3862),
.B2(n_3868),
.Y(n_6441)
);

OAI22xp5_ASAP7_75t_L g6442 ( 
.A1(n_4970),
.A2(n_4077),
.B1(n_3891),
.B2(n_4108),
.Y(n_6442)
);

OAI21xp5_ASAP7_75t_L g6443 ( 
.A1(n_4821),
.A2(n_3968),
.B(n_4087),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_5569),
.Y(n_6444)
);

INVx1_ASAP7_75t_L g6445 ( 
.A(n_5569),
.Y(n_6445)
);

OAI21x1_ASAP7_75t_L g6446 ( 
.A1(n_5258),
.A2(n_3827),
.B(n_3711),
.Y(n_6446)
);

OAI21x1_ASAP7_75t_SL g6447 ( 
.A1(n_5066),
.A2(n_3900),
.B(n_3526),
.Y(n_6447)
);

O2A1O1Ixp5_ASAP7_75t_L g6448 ( 
.A1(n_4953),
.A2(n_3879),
.B(n_3805),
.C(n_3725),
.Y(n_6448)
);

OAI21xp5_ASAP7_75t_L g6449 ( 
.A1(n_4821),
.A2(n_4087),
.B(n_4108),
.Y(n_6449)
);

NAND2xp5_ASAP7_75t_L g6450 ( 
.A(n_5073),
.B(n_4723),
.Y(n_6450)
);

OAI21xp5_ASAP7_75t_L g6451 ( 
.A1(n_4826),
.A2(n_4108),
.B(n_3725),
.Y(n_6451)
);

OAI21xp5_ASAP7_75t_L g6452 ( 
.A1(n_4826),
.A2(n_4108),
.B(n_3725),
.Y(n_6452)
);

BUFx4f_ASAP7_75t_L g6453 ( 
.A(n_5756),
.Y(n_6453)
);

A2O1A1Ixp33_ASAP7_75t_L g6454 ( 
.A1(n_4751),
.A2(n_3846),
.B(n_3471),
.C(n_3475),
.Y(n_6454)
);

OAI22xp5_ASAP7_75t_L g6455 ( 
.A1(n_4736),
.A2(n_3891),
.B1(n_4108),
.B2(n_3662),
.Y(n_6455)
);

AOI21x1_ASAP7_75t_L g6456 ( 
.A1(n_5653),
.A2(n_3891),
.B(n_4097),
.Y(n_6456)
);

OAI21x1_ASAP7_75t_L g6457 ( 
.A1(n_5262),
.A2(n_3879),
.B(n_3685),
.Y(n_6457)
);

AOI22xp33_ASAP7_75t_L g6458 ( 
.A1(n_4922),
.A2(n_4094),
.B1(n_4672),
.B2(n_3877),
.Y(n_6458)
);

NAND3xp33_ASAP7_75t_L g6459 ( 
.A(n_4836),
.B(n_4745),
.C(n_4736),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_5653),
.Y(n_6460)
);

INVx4_ASAP7_75t_L g6461 ( 
.A(n_5254),
.Y(n_6461)
);

NAND2xp5_ASAP7_75t_L g6462 ( 
.A(n_4741),
.B(n_4051),
.Y(n_6462)
);

AND2x4_ASAP7_75t_L g6463 ( 
.A(n_4749),
.B(n_4797),
.Y(n_6463)
);

BUFx2_ASAP7_75t_L g6464 ( 
.A(n_5478),
.Y(n_6464)
);

AND2x2_ASAP7_75t_L g6465 ( 
.A(n_5677),
.B(n_4051),
.Y(n_6465)
);

AOI21xp5_ASAP7_75t_L g6466 ( 
.A1(n_4802),
.A2(n_4051),
.B(n_3751),
.Y(n_6466)
);

O2A1O1Ixp5_ASAP7_75t_L g6467 ( 
.A1(n_4842),
.A2(n_4844),
.B(n_4753),
.C(n_4774),
.Y(n_6467)
);

OAI21xp33_ASAP7_75t_SL g6468 ( 
.A1(n_4844),
.A2(n_3900),
.B(n_3747),
.Y(n_6468)
);

OA21x2_ASAP7_75t_L g6469 ( 
.A1(n_5325),
.A2(n_3421),
.B(n_4707),
.Y(n_6469)
);

A2O1A1Ixp33_ASAP7_75t_L g6470 ( 
.A1(n_4757),
.A2(n_3471),
.B(n_3475),
.C(n_3846),
.Y(n_6470)
);

OAI21x1_ASAP7_75t_L g6471 ( 
.A1(n_5263),
.A2(n_3879),
.B(n_3685),
.Y(n_6471)
);

NAND2xp5_ASAP7_75t_L g6472 ( 
.A(n_5410),
.B(n_5444),
.Y(n_6472)
);

OAI21x1_ASAP7_75t_L g6473 ( 
.A1(n_5269),
.A2(n_3879),
.B(n_3685),
.Y(n_6473)
);

OAI21x1_ASAP7_75t_L g6474 ( 
.A1(n_5269),
.A2(n_3805),
.B(n_3879),
.Y(n_6474)
);

AOI21xp5_ASAP7_75t_SL g6475 ( 
.A1(n_5035),
.A2(n_4120),
.B(n_3471),
.Y(n_6475)
);

INVx2_ASAP7_75t_L g6476 ( 
.A(n_5711),
.Y(n_6476)
);

INVx4_ASAP7_75t_L g6477 ( 
.A(n_5254),
.Y(n_6477)
);

AO22x2_ASAP7_75t_L g6478 ( 
.A1(n_5078),
.A2(n_3421),
.B1(n_4707),
.B2(n_4481),
.Y(n_6478)
);

AOI221x1_ASAP7_75t_L g6479 ( 
.A1(n_4848),
.A2(n_4872),
.B1(n_5056),
.B2(n_4842),
.C(n_4906),
.Y(n_6479)
);

AND3x2_ASAP7_75t_L g6480 ( 
.A(n_5334),
.B(n_4120),
.C(n_4716),
.Y(n_6480)
);

OAI21x1_ASAP7_75t_L g6481 ( 
.A1(n_5271),
.A2(n_3752),
.B(n_3725),
.Y(n_6481)
);

O2A1O1Ixp5_ASAP7_75t_L g6482 ( 
.A1(n_4726),
.A2(n_3827),
.B(n_3805),
.C(n_3752),
.Y(n_6482)
);

INVx2_ASAP7_75t_SL g6483 ( 
.A(n_5439),
.Y(n_6483)
);

OAI21xp5_ASAP7_75t_L g6484 ( 
.A1(n_4836),
.A2(n_3805),
.B(n_3752),
.Y(n_6484)
);

AOI21x1_ASAP7_75t_L g6485 ( 
.A1(n_5711),
.A2(n_4120),
.B(n_4105),
.Y(n_6485)
);

HB1xp67_ASAP7_75t_L g6486 ( 
.A(n_5747),
.Y(n_6486)
);

NOR2xp33_ASAP7_75t_L g6487 ( 
.A(n_4819),
.B(n_3900),
.Y(n_6487)
);

AOI22xp5_ASAP7_75t_L g6488 ( 
.A1(n_4755),
.A2(n_3880),
.B1(n_3877),
.B2(n_3527),
.Y(n_6488)
);

AOI21x1_ASAP7_75t_L g6489 ( 
.A1(n_5908),
.A2(n_4120),
.B(n_4105),
.Y(n_6489)
);

AOI21xp5_ASAP7_75t_L g6490 ( 
.A1(n_4843),
.A2(n_3751),
.B(n_3915),
.Y(n_6490)
);

AOI21xp5_ASAP7_75t_L g6491 ( 
.A1(n_4850),
.A2(n_3751),
.B(n_3915),
.Y(n_6491)
);

AOI21x1_ASAP7_75t_L g6492 ( 
.A1(n_5908),
.A2(n_4120),
.B(n_4105),
.Y(n_6492)
);

BUFx10_ASAP7_75t_L g6493 ( 
.A(n_5276),
.Y(n_6493)
);

AOI21x1_ASAP7_75t_L g6494 ( 
.A1(n_5915),
.A2(n_4256),
.B(n_4481),
.Y(n_6494)
);

NOR2xp67_ASAP7_75t_L g6495 ( 
.A(n_5065),
.B(n_3861),
.Y(n_6495)
);

INVx2_ASAP7_75t_L g6496 ( 
.A(n_5915),
.Y(n_6496)
);

AOI21xp5_ASAP7_75t_L g6497 ( 
.A1(n_4864),
.A2(n_3915),
.B(n_3751),
.Y(n_6497)
);

OAI21x1_ASAP7_75t_L g6498 ( 
.A1(n_5271),
.A2(n_4865),
.B(n_4864),
.Y(n_6498)
);

CKINVDCx11_ASAP7_75t_R g6499 ( 
.A(n_5171),
.Y(n_6499)
);

NAND2xp5_ASAP7_75t_L g6500 ( 
.A(n_5054),
.B(n_3822),
.Y(n_6500)
);

A2O1A1Ixp33_ASAP7_75t_L g6501 ( 
.A1(n_4757),
.A2(n_3475),
.B(n_3743),
.C(n_3673),
.Y(n_6501)
);

AOI21x1_ASAP7_75t_L g6502 ( 
.A1(n_5920),
.A2(n_5923),
.B(n_5052),
.Y(n_6502)
);

AOI21xp5_ASAP7_75t_L g6503 ( 
.A1(n_4865),
.A2(n_3751),
.B(n_3915),
.Y(n_6503)
);

OAI21xp5_ASAP7_75t_L g6504 ( 
.A1(n_4768),
.A2(n_3805),
.B(n_3711),
.Y(n_6504)
);

AOI21x1_ASAP7_75t_L g6505 ( 
.A1(n_5920),
.A2(n_4256),
.B(n_3551),
.Y(n_6505)
);

AOI21xp33_ASAP7_75t_L g6506 ( 
.A1(n_4849),
.A2(n_3938),
.B(n_3785),
.Y(n_6506)
);

AND2x2_ASAP7_75t_L g6507 ( 
.A(n_5716),
.B(n_4045),
.Y(n_6507)
);

OAI21x1_ASAP7_75t_L g6508 ( 
.A1(n_4867),
.A2(n_3861),
.B(n_3752),
.Y(n_6508)
);

AND2x2_ASAP7_75t_L g6509 ( 
.A(n_5716),
.B(n_5783),
.Y(n_6509)
);

NOR2xp67_ASAP7_75t_L g6510 ( 
.A(n_4874),
.B(n_3861),
.Y(n_6510)
);

AOI22xp5_ASAP7_75t_L g6511 ( 
.A1(n_4745),
.A2(n_3880),
.B1(n_3877),
.B2(n_3536),
.Y(n_6511)
);

AND2x2_ASAP7_75t_L g6512 ( 
.A(n_5783),
.B(n_4045),
.Y(n_6512)
);

OA21x2_ASAP7_75t_L g6513 ( 
.A1(n_5325),
.A2(n_3551),
.B(n_3999),
.Y(n_6513)
);

A2O1A1Ixp33_ASAP7_75t_L g6514 ( 
.A1(n_5111),
.A2(n_3743),
.B(n_3566),
.C(n_3991),
.Y(n_6514)
);

NAND2xp5_ASAP7_75t_L g6515 ( 
.A(n_5059),
.B(n_3783),
.Y(n_6515)
);

BUFx6f_ASAP7_75t_L g6516 ( 
.A(n_4758),
.Y(n_6516)
);

OAI21x1_ASAP7_75t_L g6517 ( 
.A1(n_4867),
.A2(n_3861),
.B(n_3752),
.Y(n_6517)
);

OAI22xp5_ASAP7_75t_L g6518 ( 
.A1(n_4922),
.A2(n_3915),
.B1(n_3751),
.B2(n_3662),
.Y(n_6518)
);

AOI21xp5_ASAP7_75t_L g6519 ( 
.A1(n_4894),
.A2(n_3915),
.B(n_3751),
.Y(n_6519)
);

BUFx3_ASAP7_75t_L g6520 ( 
.A(n_5573),
.Y(n_6520)
);

OAI21x1_ASAP7_75t_L g6521 ( 
.A1(n_5202),
.A2(n_5249),
.B(n_5223),
.Y(n_6521)
);

NAND2xp5_ASAP7_75t_L g6522 ( 
.A(n_4982),
.B(n_3785),
.Y(n_6522)
);

CKINVDCx5p33_ASAP7_75t_R g6523 ( 
.A(n_5079),
.Y(n_6523)
);

NOR2xp33_ASAP7_75t_L g6524 ( 
.A(n_4819),
.B(n_3526),
.Y(n_6524)
);

AND2x2_ASAP7_75t_L g6525 ( 
.A(n_5783),
.B(n_4045),
.Y(n_6525)
);

INVx1_ASAP7_75t_L g6526 ( 
.A(n_5771),
.Y(n_6526)
);

NAND3xp33_ASAP7_75t_SL g6527 ( 
.A(n_4848),
.B(n_4872),
.C(n_5015),
.Y(n_6527)
);

AND2x2_ASAP7_75t_SL g6528 ( 
.A(n_5056),
.B(n_3947),
.Y(n_6528)
);

INVx1_ASAP7_75t_L g6529 ( 
.A(n_5771),
.Y(n_6529)
);

NAND2xp5_ASAP7_75t_L g6530 ( 
.A(n_4982),
.B(n_3785),
.Y(n_6530)
);

NAND2x1p5_ASAP7_75t_L g6531 ( 
.A(n_6201),
.B(n_3915),
.Y(n_6531)
);

CKINVDCx5p33_ASAP7_75t_R g6532 ( 
.A(n_5979),
.Y(n_6532)
);

AO21x1_ASAP7_75t_L g6533 ( 
.A1(n_5353),
.A2(n_3526),
.B(n_3527),
.Y(n_6533)
);

NAND2xp5_ASAP7_75t_L g6534 ( 
.A(n_5012),
.B(n_5025),
.Y(n_6534)
);

AO31x2_ASAP7_75t_L g6535 ( 
.A1(n_6095),
.A2(n_3527),
.A3(n_3536),
.B(n_3747),
.Y(n_6535)
);

NAND2xp5_ASAP7_75t_L g6536 ( 
.A(n_5012),
.B(n_3928),
.Y(n_6536)
);

NOR2xp33_ASAP7_75t_L g6537 ( 
.A(n_5091),
.B(n_4999),
.Y(n_6537)
);

INVx3_ASAP7_75t_L g6538 ( 
.A(n_5975),
.Y(n_6538)
);

OAI21xp5_ASAP7_75t_L g6539 ( 
.A1(n_5121),
.A2(n_3861),
.B(n_3751),
.Y(n_6539)
);

OAI21x1_ASAP7_75t_L g6540 ( 
.A1(n_5202),
.A2(n_4101),
.B(n_3999),
.Y(n_6540)
);

AND2x2_ASAP7_75t_L g6541 ( 
.A(n_5802),
.B(n_5810),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_5775),
.Y(n_6542)
);

A2O1A1Ixp33_ASAP7_75t_L g6543 ( 
.A1(n_5111),
.A2(n_3566),
.B(n_3915),
.C(n_3662),
.Y(n_6543)
);

AND2x4_ASAP7_75t_L g6544 ( 
.A(n_4749),
.B(n_4797),
.Y(n_6544)
);

A2O1A1Ixp33_ASAP7_75t_L g6545 ( 
.A1(n_5127),
.A2(n_3566),
.B(n_3662),
.C(n_3830),
.Y(n_6545)
);

OAI21xp5_ASAP7_75t_L g6546 ( 
.A1(n_4897),
.A2(n_3662),
.B(n_3877),
.Y(n_6546)
);

OAI21xp5_ASAP7_75t_L g6547 ( 
.A1(n_4897),
.A2(n_3662),
.B(n_3877),
.Y(n_6547)
);

OAI21xp5_ASAP7_75t_L g6548 ( 
.A1(n_4906),
.A2(n_3662),
.B(n_3877),
.Y(n_6548)
);

NAND2xp5_ASAP7_75t_L g6549 ( 
.A(n_5025),
.B(n_3947),
.Y(n_6549)
);

AOI21xp5_ASAP7_75t_L g6550 ( 
.A1(n_4894),
.A2(n_3947),
.B(n_3928),
.Y(n_6550)
);

AND2x4_ASAP7_75t_L g6551 ( 
.A(n_4797),
.B(n_3527),
.Y(n_6551)
);

NAND2xp5_ASAP7_75t_L g6552 ( 
.A(n_4743),
.B(n_3947),
.Y(n_6552)
);

OAI21x1_ASAP7_75t_L g6553 ( 
.A1(n_5223),
.A2(n_5277),
.B(n_5249),
.Y(n_6553)
);

OAI21x1_ASAP7_75t_L g6554 ( 
.A1(n_5277),
.A2(n_4101),
.B(n_3608),
.Y(n_6554)
);

OAI21x1_ASAP7_75t_L g6555 ( 
.A1(n_5282),
.A2(n_5459),
.B(n_5456),
.Y(n_6555)
);

BUFx6f_ASAP7_75t_L g6556 ( 
.A(n_4758),
.Y(n_6556)
);

NAND2xp5_ASAP7_75t_L g6557 ( 
.A(n_4743),
.B(n_3947),
.Y(n_6557)
);

INVx8_ASAP7_75t_L g6558 ( 
.A(n_5270),
.Y(n_6558)
);

A2O1A1Ixp33_ASAP7_75t_L g6559 ( 
.A1(n_5127),
.A2(n_3830),
.B(n_3938),
.C(n_3928),
.Y(n_6559)
);

NAND2xp5_ASAP7_75t_L g6560 ( 
.A(n_4746),
.B(n_3947),
.Y(n_6560)
);

OAI21xp5_ASAP7_75t_L g6561 ( 
.A1(n_4908),
.A2(n_3877),
.B(n_3880),
.Y(n_6561)
);

AOI21xp5_ASAP7_75t_L g6562 ( 
.A1(n_5199),
.A2(n_3822),
.B(n_3928),
.Y(n_6562)
);

NAND2xp5_ASAP7_75t_L g6563 ( 
.A(n_4746),
.B(n_3947),
.Y(n_6563)
);

OAI21x1_ASAP7_75t_L g6564 ( 
.A1(n_5282),
.A2(n_4101),
.B(n_3880),
.Y(n_6564)
);

OAI21x1_ASAP7_75t_L g6565 ( 
.A1(n_5456),
.A2(n_4101),
.B(n_3880),
.Y(n_6565)
);

NAND2xp5_ASAP7_75t_L g6566 ( 
.A(n_4760),
.B(n_3947),
.Y(n_6566)
);

NAND2xp5_ASAP7_75t_L g6567 ( 
.A(n_4760),
.B(n_3938),
.Y(n_6567)
);

NAND2xp5_ASAP7_75t_L g6568 ( 
.A(n_4773),
.B(n_3938),
.Y(n_6568)
);

AOI21xp5_ASAP7_75t_L g6569 ( 
.A1(n_5199),
.A2(n_3822),
.B(n_3938),
.Y(n_6569)
);

AND2x2_ASAP7_75t_L g6570 ( 
.A(n_5802),
.B(n_4045),
.Y(n_6570)
);

OAI21xp5_ASAP7_75t_L g6571 ( 
.A1(n_4908),
.A2(n_3880),
.B(n_3536),
.Y(n_6571)
);

AOI21xp5_ASAP7_75t_L g6572 ( 
.A1(n_5206),
.A2(n_3785),
.B(n_3938),
.Y(n_6572)
);

INVx2_ASAP7_75t_SL g6573 ( 
.A(n_5439),
.Y(n_6573)
);

AND2x2_ASAP7_75t_L g6574 ( 
.A(n_5802),
.B(n_3785),
.Y(n_6574)
);

AOI21x1_ASAP7_75t_L g6575 ( 
.A1(n_4990),
.A2(n_3785),
.B(n_3928),
.Y(n_6575)
);

AOI21xp5_ASAP7_75t_L g6576 ( 
.A1(n_5206),
.A2(n_3785),
.B(n_3851),
.Y(n_6576)
);

CKINVDCx5p33_ASAP7_75t_R g6577 ( 
.A(n_4866),
.Y(n_6577)
);

OAI21x1_ASAP7_75t_L g6578 ( 
.A1(n_5459),
.A2(n_5477),
.B(n_5476),
.Y(n_6578)
);

INVx1_ASAP7_75t_SL g6579 ( 
.A(n_4911),
.Y(n_6579)
);

INVx4_ASAP7_75t_L g6580 ( 
.A(n_6201),
.Y(n_6580)
);

BUFx12f_ASAP7_75t_L g6581 ( 
.A(n_5259),
.Y(n_6581)
);

NAND2xp5_ASAP7_75t_L g6582 ( 
.A(n_4775),
.B(n_3783),
.Y(n_6582)
);

AOI21xp5_ASAP7_75t_L g6583 ( 
.A1(n_5072),
.A2(n_3783),
.B(n_3851),
.Y(n_6583)
);

AOI21xp5_ASAP7_75t_SL g6584 ( 
.A1(n_5095),
.A2(n_4103),
.B(n_3536),
.Y(n_6584)
);

INVx3_ASAP7_75t_L g6585 ( 
.A(n_5975),
.Y(n_6585)
);

NAND2xp5_ASAP7_75t_L g6586 ( 
.A(n_4775),
.B(n_3783),
.Y(n_6586)
);

OAI22xp5_ASAP7_75t_L g6587 ( 
.A1(n_5078),
.A2(n_3851),
.B1(n_3928),
.B2(n_3783),
.Y(n_6587)
);

A2O1A1Ixp33_ASAP7_75t_L g6588 ( 
.A1(n_5133),
.A2(n_3830),
.B(n_3928),
.C(n_3851),
.Y(n_6588)
);

NAND2xp5_ASAP7_75t_L g6589 ( 
.A(n_4784),
.B(n_4787),
.Y(n_6589)
);

OAI21xp5_ASAP7_75t_L g6590 ( 
.A1(n_4910),
.A2(n_3880),
.B(n_3536),
.Y(n_6590)
);

NAND2xp5_ASAP7_75t_L g6591 ( 
.A(n_4784),
.B(n_3822),
.Y(n_6591)
);

AOI21xp5_ASAP7_75t_L g6592 ( 
.A1(n_5476),
.A2(n_3822),
.B(n_3851),
.Y(n_6592)
);

OAI22xp5_ASAP7_75t_L g6593 ( 
.A1(n_5000),
.A2(n_3851),
.B1(n_3928),
.B2(n_3783),
.Y(n_6593)
);

AOI21x1_ASAP7_75t_L g6594 ( 
.A1(n_4990),
.A2(n_3783),
.B(n_3880),
.Y(n_6594)
);

CKINVDCx11_ASAP7_75t_R g6595 ( 
.A(n_5865),
.Y(n_6595)
);

AOI21xp5_ASAP7_75t_L g6596 ( 
.A1(n_5477),
.A2(n_4013),
.B(n_4033),
.Y(n_6596)
);

INVx3_ASAP7_75t_L g6597 ( 
.A(n_5975),
.Y(n_6597)
);

NOR2xp33_ASAP7_75t_L g6598 ( 
.A(n_4999),
.B(n_3527),
.Y(n_6598)
);

OAI21x1_ASAP7_75t_L g6599 ( 
.A1(n_5481),
.A2(n_4101),
.B(n_3880),
.Y(n_6599)
);

OAI22x1_ASAP7_75t_L g6600 ( 
.A1(n_4822),
.A2(n_3747),
.B1(n_4103),
.B2(n_4014),
.Y(n_6600)
);

AOI21xp5_ASAP7_75t_L g6601 ( 
.A1(n_5481),
.A2(n_4020),
.B(n_4033),
.Y(n_6601)
);

OR2x6_ASAP7_75t_L g6602 ( 
.A(n_4797),
.B(n_5285),
.Y(n_6602)
);

OAI21xp5_ASAP7_75t_L g6603 ( 
.A1(n_4910),
.A2(n_4020),
.B(n_4033),
.Y(n_6603)
);

AOI21xp5_ASAP7_75t_L g6604 ( 
.A1(n_5484),
.A2(n_4013),
.B(n_3985),
.Y(n_6604)
);

AOI22xp33_ASAP7_75t_SL g6605 ( 
.A1(n_4942),
.A2(n_4094),
.B1(n_4672),
.B2(n_4024),
.Y(n_6605)
);

AOI21xp5_ASAP7_75t_L g6606 ( 
.A1(n_5484),
.A2(n_4012),
.B(n_4013),
.Y(n_6606)
);

INVx4_ASAP7_75t_L g6607 ( 
.A(n_6201),
.Y(n_6607)
);

OAI22xp5_ASAP7_75t_L g6608 ( 
.A1(n_4920),
.A2(n_3830),
.B1(n_3985),
.B2(n_4012),
.Y(n_6608)
);

OAI21x1_ASAP7_75t_SL g6609 ( 
.A1(n_5066),
.A2(n_4103),
.B(n_4012),
.Y(n_6609)
);

OAI21x1_ASAP7_75t_L g6610 ( 
.A1(n_5491),
.A2(n_4103),
.B(n_3985),
.Y(n_6610)
);

OR2x2_ASAP7_75t_L g6611 ( 
.A(n_5379),
.B(n_4020),
.Y(n_6611)
);

CKINVDCx5p33_ASAP7_75t_R g6612 ( 
.A(n_5682),
.Y(n_6612)
);

OAI22xp5_ASAP7_75t_L g6613 ( 
.A1(n_4916),
.A2(n_4000),
.B1(n_4103),
.B2(n_3878),
.Y(n_6613)
);

NAND2xp5_ASAP7_75t_L g6614 ( 
.A(n_4787),
.B(n_4794),
.Y(n_6614)
);

OR2x2_ASAP7_75t_L g6615 ( 
.A(n_5404),
.B(n_4140),
.Y(n_6615)
);

OAI21xp5_ASAP7_75t_L g6616 ( 
.A1(n_4913),
.A2(n_4140),
.B(n_3712),
.Y(n_6616)
);

AND2x2_ASAP7_75t_L g6617 ( 
.A(n_5810),
.B(n_3712),
.Y(n_6617)
);

AO31x2_ASAP7_75t_L g6618 ( 
.A1(n_6095),
.A2(n_6105),
.A3(n_5250),
.B(n_5192),
.Y(n_6618)
);

NAND2xp5_ASAP7_75t_L g6619 ( 
.A(n_4794),
.B(n_4796),
.Y(n_6619)
);

AOI21xp5_ASAP7_75t_SL g6620 ( 
.A1(n_4947),
.A2(n_5469),
.B(n_5464),
.Y(n_6620)
);

AOI21xp5_ASAP7_75t_L g6621 ( 
.A1(n_5491),
.A2(n_5521),
.B(n_5512),
.Y(n_6621)
);

AND2x2_ASAP7_75t_L g6622 ( 
.A(n_5810),
.B(n_5852),
.Y(n_6622)
);

OR2x6_ASAP7_75t_L g6623 ( 
.A(n_5285),
.B(n_5270),
.Y(n_6623)
);

AOI21xp5_ASAP7_75t_L g6624 ( 
.A1(n_5512),
.A2(n_5535),
.B(n_5521),
.Y(n_6624)
);

OAI21x1_ASAP7_75t_L g6625 ( 
.A1(n_5535),
.A2(n_5554),
.B(n_5548),
.Y(n_6625)
);

AOI21x1_ASAP7_75t_SL g6626 ( 
.A1(n_5450),
.A2(n_5462),
.B(n_5461),
.Y(n_6626)
);

INVx1_ASAP7_75t_SL g6627 ( 
.A(n_5149),
.Y(n_6627)
);

OAI21x1_ASAP7_75t_L g6628 ( 
.A1(n_5548),
.A2(n_5561),
.B(n_5554),
.Y(n_6628)
);

CKINVDCx5p33_ASAP7_75t_R g6629 ( 
.A(n_4790),
.Y(n_6629)
);

O2A1O1Ixp5_ASAP7_75t_L g6630 ( 
.A1(n_4956),
.A2(n_4946),
.B(n_4935),
.C(n_5201),
.Y(n_6630)
);

OAI21x1_ASAP7_75t_L g6631 ( 
.A1(n_5561),
.A2(n_5574),
.B(n_5568),
.Y(n_6631)
);

NAND2xp5_ASAP7_75t_SL g6632 ( 
.A(n_4989),
.B(n_4902),
.Y(n_6632)
);

INVxp67_ASAP7_75t_L g6633 ( 
.A(n_5243),
.Y(n_6633)
);

NOR2x1_ASAP7_75t_L g6634 ( 
.A(n_5414),
.B(n_4829),
.Y(n_6634)
);

OAI21x1_ASAP7_75t_L g6635 ( 
.A1(n_5568),
.A2(n_5577),
.B(n_5574),
.Y(n_6635)
);

NAND2xp5_ASAP7_75t_L g6636 ( 
.A(n_4796),
.B(n_4803),
.Y(n_6636)
);

AO31x2_ASAP7_75t_L g6637 ( 
.A1(n_6095),
.A2(n_6105),
.A3(n_5250),
.B(n_5192),
.Y(n_6637)
);

OAI21x1_ASAP7_75t_L g6638 ( 
.A1(n_5577),
.A2(n_5611),
.B(n_5590),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_5775),
.Y(n_6639)
);

BUFx6f_ASAP7_75t_L g6640 ( 
.A(n_4758),
.Y(n_6640)
);

BUFx12f_ASAP7_75t_L g6641 ( 
.A(n_5259),
.Y(n_6641)
);

OAI21xp33_ASAP7_75t_L g6642 ( 
.A1(n_4998),
.A2(n_5034),
.B(n_4858),
.Y(n_6642)
);

OAI21xp5_ASAP7_75t_L g6643 ( 
.A1(n_4913),
.A2(n_4926),
.B(n_4914),
.Y(n_6643)
);

INVx4_ASAP7_75t_L g6644 ( 
.A(n_6201),
.Y(n_6644)
);

OAI21x1_ASAP7_75t_L g6645 ( 
.A1(n_5590),
.A2(n_5614),
.B(n_5611),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_5775),
.Y(n_6646)
);

AOI21x1_ASAP7_75t_L g6647 ( 
.A1(n_5052),
.A2(n_5624),
.B(n_5614),
.Y(n_6647)
);

BUFx8_ASAP7_75t_SL g6648 ( 
.A(n_5865),
.Y(n_6648)
);

NAND2xp5_ASAP7_75t_L g6649 ( 
.A(n_4803),
.B(n_4805),
.Y(n_6649)
);

OAI21x1_ASAP7_75t_L g6650 ( 
.A1(n_5627),
.A2(n_5642),
.B(n_5630),
.Y(n_6650)
);

OAI21x1_ASAP7_75t_L g6651 ( 
.A1(n_5642),
.A2(n_5650),
.B(n_5644),
.Y(n_6651)
);

AND2x4_ASAP7_75t_L g6652 ( 
.A(n_5921),
.B(n_5924),
.Y(n_6652)
);

INVx1_ASAP7_75t_L g6653 ( 
.A(n_5775),
.Y(n_6653)
);

NAND2xp5_ASAP7_75t_SL g6654 ( 
.A(n_4989),
.B(n_4902),
.Y(n_6654)
);

NAND3x1_ASAP7_75t_L g6655 ( 
.A(n_4885),
.B(n_4918),
.C(n_5356),
.Y(n_6655)
);

OAI21x1_ASAP7_75t_L g6656 ( 
.A1(n_5660),
.A2(n_5669),
.B(n_5662),
.Y(n_6656)
);

AOI21x1_ASAP7_75t_L g6657 ( 
.A1(n_5662),
.A2(n_5671),
.B(n_5669),
.Y(n_6657)
);

A2O1A1Ixp33_ASAP7_75t_L g6658 ( 
.A1(n_5133),
.A2(n_5169),
.B(n_4947),
.C(n_5433),
.Y(n_6658)
);

OAI21x1_ASAP7_75t_L g6659 ( 
.A1(n_5671),
.A2(n_5689),
.B(n_5685),
.Y(n_6659)
);

INVx1_ASAP7_75t_SL g6660 ( 
.A(n_5149),
.Y(n_6660)
);

AND2x2_ASAP7_75t_L g6661 ( 
.A(n_5852),
.B(n_5399),
.Y(n_6661)
);

OAI21x1_ASAP7_75t_L g6662 ( 
.A1(n_5685),
.A2(n_5703),
.B(n_5689),
.Y(n_6662)
);

AOI21xp33_ASAP7_75t_L g6663 ( 
.A1(n_4849),
.A2(n_4877),
.B(n_4933),
.Y(n_6663)
);

AND2x2_ASAP7_75t_L g6664 ( 
.A(n_5852),
.B(n_5399),
.Y(n_6664)
);

AOI21xp5_ASAP7_75t_L g6665 ( 
.A1(n_5703),
.A2(n_5709),
.B(n_5708),
.Y(n_6665)
);

NOR2xp33_ASAP7_75t_L g6666 ( 
.A(n_4779),
.B(n_4781),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_4874),
.Y(n_6667)
);

AOI21xp5_ASAP7_75t_L g6668 ( 
.A1(n_5708),
.A2(n_5724),
.B(n_5709),
.Y(n_6668)
);

NAND3x1_ASAP7_75t_L g6669 ( 
.A(n_4885),
.B(n_4918),
.C(n_5449),
.Y(n_6669)
);

OAI22x1_ASAP7_75t_L g6670 ( 
.A1(n_4822),
.A2(n_4863),
.B1(n_5402),
.B2(n_5449),
.Y(n_6670)
);

NAND2xp5_ASAP7_75t_L g6671 ( 
.A(n_4805),
.B(n_4813),
.Y(n_6671)
);

AOI21xp5_ASAP7_75t_L g6672 ( 
.A1(n_5724),
.A2(n_5750),
.B(n_5736),
.Y(n_6672)
);

O2A1O1Ixp5_ASAP7_75t_L g6673 ( 
.A1(n_4956),
.A2(n_4935),
.B(n_4946),
.C(n_5374),
.Y(n_6673)
);

AOI21xp5_ASAP7_75t_L g6674 ( 
.A1(n_5736),
.A2(n_5754),
.B(n_5750),
.Y(n_6674)
);

AOI21xp33_ASAP7_75t_L g6675 ( 
.A1(n_4877),
.A2(n_4933),
.B(n_5169),
.Y(n_6675)
);

NAND2xp5_ASAP7_75t_L g6676 ( 
.A(n_4813),
.B(n_4820),
.Y(n_6676)
);

BUFx6f_ASAP7_75t_L g6677 ( 
.A(n_4758),
.Y(n_6677)
);

A2O1A1Ixp33_ASAP7_75t_L g6678 ( 
.A1(n_5433),
.A2(n_4914),
.B(n_4931),
.C(n_4926),
.Y(n_6678)
);

AOI21xp5_ASAP7_75t_SL g6679 ( 
.A1(n_5392),
.A2(n_5176),
.B(n_5045),
.Y(n_6679)
);

BUFx2_ASAP7_75t_L g6680 ( 
.A(n_5525),
.Y(n_6680)
);

AOI21xp5_ASAP7_75t_L g6681 ( 
.A1(n_5754),
.A2(n_5782),
.B(n_5769),
.Y(n_6681)
);

O2A1O1Ixp5_ASAP7_75t_L g6682 ( 
.A1(n_5374),
.A2(n_4936),
.B(n_4940),
.C(n_4931),
.Y(n_6682)
);

INVx8_ASAP7_75t_L g6683 ( 
.A(n_5270),
.Y(n_6683)
);

INVx1_ASAP7_75t_SL g6684 ( 
.A(n_5156),
.Y(n_6684)
);

AOI21x1_ASAP7_75t_L g6685 ( 
.A1(n_5769),
.A2(n_5782),
.B(n_5083),
.Y(n_6685)
);

OAI22xp5_ASAP7_75t_L g6686 ( 
.A1(n_4916),
.A2(n_4780),
.B1(n_4788),
.B2(n_4770),
.Y(n_6686)
);

NOR2xp33_ASAP7_75t_SL g6687 ( 
.A(n_4728),
.B(n_5538),
.Y(n_6687)
);

AND2x4_ASAP7_75t_L g6688 ( 
.A(n_5921),
.B(n_5924),
.Y(n_6688)
);

OAI21xp5_ASAP7_75t_L g6689 ( 
.A1(n_4936),
.A2(n_4945),
.B(n_4940),
.Y(n_6689)
);

AND2x4_ASAP7_75t_L g6690 ( 
.A(n_5924),
.B(n_4744),
.Y(n_6690)
);

AND2x4_ASAP7_75t_L g6691 ( 
.A(n_4744),
.B(n_4752),
.Y(n_6691)
);

AND2x4_ASAP7_75t_L g6692 ( 
.A(n_4744),
.B(n_4752),
.Y(n_6692)
);

NAND2xp5_ASAP7_75t_SL g6693 ( 
.A(n_4998),
.B(n_5034),
.Y(n_6693)
);

OAI21xp5_ASAP7_75t_L g6694 ( 
.A1(n_4945),
.A2(n_4955),
.B(n_4812),
.Y(n_6694)
);

AOI21xp5_ASAP7_75t_L g6695 ( 
.A1(n_4923),
.A2(n_5415),
.B(n_5411),
.Y(n_6695)
);

NAND2xp33_ASAP7_75t_L g6696 ( 
.A(n_4858),
.B(n_5389),
.Y(n_6696)
);

OAI21x1_ASAP7_75t_L g6697 ( 
.A1(n_5081),
.A2(n_5083),
.B(n_5786),
.Y(n_6697)
);

OAI21x1_ASAP7_75t_L g6698 ( 
.A1(n_5081),
.A2(n_5787),
.B(n_5786),
.Y(n_6698)
);

NAND2xp5_ASAP7_75t_L g6699 ( 
.A(n_4820),
.B(n_4837),
.Y(n_6699)
);

BUFx6f_ASAP7_75t_L g6700 ( 
.A(n_4765),
.Y(n_6700)
);

AND2x2_ASAP7_75t_L g6701 ( 
.A(n_5399),
.B(n_5405),
.Y(n_6701)
);

INVx1_ASAP7_75t_L g6702 ( 
.A(n_4886),
.Y(n_6702)
);

INVxp67_ASAP7_75t_L g6703 ( 
.A(n_5243),
.Y(n_6703)
);

OAI21xp5_ASAP7_75t_L g6704 ( 
.A1(n_4955),
.A2(n_4812),
.B(n_4964),
.Y(n_6704)
);

OAI21x1_ASAP7_75t_L g6705 ( 
.A1(n_5787),
.A2(n_5797),
.B(n_5791),
.Y(n_6705)
);

AND3x2_ASAP7_75t_L g6706 ( 
.A(n_5334),
.B(n_5916),
.C(n_5538),
.Y(n_6706)
);

INVx2_ASAP7_75t_SL g6707 ( 
.A(n_5439),
.Y(n_6707)
);

AOI21xp5_ASAP7_75t_L g6708 ( 
.A1(n_5411),
.A2(n_5416),
.B(n_5415),
.Y(n_6708)
);

OAI21xp5_ASAP7_75t_L g6709 ( 
.A1(n_4964),
.A2(n_5224),
.B(n_4809),
.Y(n_6709)
);

OAI21x1_ASAP7_75t_L g6710 ( 
.A1(n_5791),
.A2(n_5797),
.B(n_4979),
.Y(n_6710)
);

OAI21xp33_ASAP7_75t_L g6711 ( 
.A1(n_4810),
.A2(n_4809),
.B(n_5022),
.Y(n_6711)
);

OAI21x1_ASAP7_75t_L g6712 ( 
.A1(n_4965),
.A2(n_4979),
.B(n_5364),
.Y(n_6712)
);

INVx4_ASAP7_75t_L g6713 ( 
.A(n_6201),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_4886),
.Y(n_6714)
);

INVx1_ASAP7_75t_L g6715 ( 
.A(n_4891),
.Y(n_6715)
);

INVx2_ASAP7_75t_L g6716 ( 
.A(n_5959),
.Y(n_6716)
);

OAI21x1_ASAP7_75t_L g6717 ( 
.A1(n_4965),
.A2(n_5364),
.B(n_5320),
.Y(n_6717)
);

OAI21xp5_ASAP7_75t_L g6718 ( 
.A1(n_5108),
.A2(n_5117),
.B(n_5414),
.Y(n_6718)
);

NAND2xp5_ASAP7_75t_L g6719 ( 
.A(n_4837),
.B(n_4847),
.Y(n_6719)
);

NAND2xp5_ASAP7_75t_L g6720 ( 
.A(n_4847),
.B(n_4851),
.Y(n_6720)
);

AND2x2_ASAP7_75t_L g6721 ( 
.A(n_5405),
.B(n_5443),
.Y(n_6721)
);

INVx1_ASAP7_75t_SL g6722 ( 
.A(n_5156),
.Y(n_6722)
);

NOR2x1_ASAP7_75t_L g6723 ( 
.A(n_4829),
.B(n_4898),
.Y(n_6723)
);

INVx1_ASAP7_75t_L g6724 ( 
.A(n_4891),
.Y(n_6724)
);

INVx1_ASAP7_75t_L g6725 ( 
.A(n_4941),
.Y(n_6725)
);

OA22x2_ASAP7_75t_L g6726 ( 
.A1(n_5234),
.A2(n_5389),
.B1(n_5466),
.B2(n_6229),
.Y(n_6726)
);

AND2x4_ASAP7_75t_L g6727 ( 
.A(n_4752),
.B(n_4756),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_L g6728 ( 
.A(n_4851),
.B(n_4856),
.Y(n_6728)
);

A2O1A1Ixp33_ASAP7_75t_L g6729 ( 
.A1(n_5234),
.A2(n_5074),
.B(n_5027),
.C(n_5141),
.Y(n_6729)
);

NOR2x1_ASAP7_75t_SL g6730 ( 
.A(n_5291),
.B(n_5251),
.Y(n_6730)
);

BUFx6f_ASAP7_75t_L g6731 ( 
.A(n_4765),
.Y(n_6731)
);

INVx6_ASAP7_75t_L g6732 ( 
.A(n_6201),
.Y(n_6732)
);

AOI21xp5_ASAP7_75t_L g6733 ( 
.A1(n_5416),
.A2(n_5424),
.B(n_5418),
.Y(n_6733)
);

NAND2xp5_ASAP7_75t_L g6734 ( 
.A(n_4856),
.B(n_4859),
.Y(n_6734)
);

AO31x2_ASAP7_75t_L g6735 ( 
.A1(n_6105),
.A2(n_5195),
.A3(n_5396),
.B(n_5383),
.Y(n_6735)
);

A2O1A1Ixp33_ASAP7_75t_L g6736 ( 
.A1(n_5141),
.A2(n_4747),
.B(n_4722),
.C(n_4728),
.Y(n_6736)
);

AOI21xp5_ASAP7_75t_L g6737 ( 
.A1(n_5418),
.A2(n_5426),
.B(n_5424),
.Y(n_6737)
);

OAI21xp5_ASAP7_75t_L g6738 ( 
.A1(n_4828),
.A2(n_4878),
.B(n_4875),
.Y(n_6738)
);

AOI21xp5_ASAP7_75t_L g6739 ( 
.A1(n_5426),
.A2(n_5436),
.B(n_5431),
.Y(n_6739)
);

AOI21xp33_ASAP7_75t_L g6740 ( 
.A1(n_5137),
.A2(n_5341),
.B(n_4863),
.Y(n_6740)
);

OAI21xp5_ASAP7_75t_L g6741 ( 
.A1(n_4828),
.A2(n_4878),
.B(n_4875),
.Y(n_6741)
);

INVx1_ASAP7_75t_L g6742 ( 
.A(n_4941),
.Y(n_6742)
);

NAND2xp5_ASAP7_75t_L g6743 ( 
.A(n_4859),
.B(n_4860),
.Y(n_6743)
);

AO31x2_ASAP7_75t_L g6744 ( 
.A1(n_5195),
.A2(n_5396),
.A3(n_5383),
.B(n_5401),
.Y(n_6744)
);

A2O1A1Ixp33_ASAP7_75t_L g6745 ( 
.A1(n_5143),
.A2(n_5155),
.B(n_5178),
.C(n_5173),
.Y(n_6745)
);

OAI21x1_ASAP7_75t_SL g6746 ( 
.A1(n_5070),
.A2(n_5093),
.B(n_5085),
.Y(n_6746)
);

OAI21x1_ASAP7_75t_L g6747 ( 
.A1(n_5799),
.A2(n_6179),
.B(n_6119),
.Y(n_6747)
);

NAND3xp33_ASAP7_75t_L g6748 ( 
.A(n_4919),
.B(n_4952),
.C(n_5204),
.Y(n_6748)
);

OAI21x1_ASAP7_75t_L g6749 ( 
.A1(n_6117),
.A2(n_6120),
.B(n_6119),
.Y(n_6749)
);

INVx2_ASAP7_75t_L g6750 ( 
.A(n_5959),
.Y(n_6750)
);

AOI21xp5_ASAP7_75t_L g6751 ( 
.A1(n_5431),
.A2(n_5436),
.B(n_5042),
.Y(n_6751)
);

BUFx3_ASAP7_75t_L g6752 ( 
.A(n_5573),
.Y(n_6752)
);

AOI21xp5_ASAP7_75t_L g6753 ( 
.A1(n_4971),
.A2(n_5070),
.B(n_5039),
.Y(n_6753)
);

OAI21x1_ASAP7_75t_L g6754 ( 
.A1(n_6117),
.A2(n_6139),
.B(n_6120),
.Y(n_6754)
);

O2A1O1Ixp33_ASAP7_75t_L g6755 ( 
.A1(n_4823),
.A2(n_4948),
.B(n_4825),
.C(n_4912),
.Y(n_6755)
);

BUFx6f_ASAP7_75t_SL g6756 ( 
.A(n_4765),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_L g6757 ( 
.A(n_4860),
.B(n_4861),
.Y(n_6757)
);

OAI21x1_ASAP7_75t_L g6758 ( 
.A1(n_6139),
.A2(n_6146),
.B(n_6144),
.Y(n_6758)
);

INVx2_ASAP7_75t_L g6759 ( 
.A(n_5959),
.Y(n_6759)
);

OAI22x1_ASAP7_75t_L g6760 ( 
.A1(n_5402),
.A2(n_6032),
.B1(n_6041),
.B2(n_6034),
.Y(n_6760)
);

NAND2xp5_ASAP7_75t_L g6761 ( 
.A(n_4861),
.B(n_4869),
.Y(n_6761)
);

AO31x2_ASAP7_75t_L g6762 ( 
.A1(n_5401),
.A2(n_5377),
.A3(n_5353),
.B(n_5368),
.Y(n_6762)
);

NAND2xp5_ASAP7_75t_L g6763 ( 
.A(n_4869),
.B(n_4871),
.Y(n_6763)
);

OAI21x1_ASAP7_75t_L g6764 ( 
.A1(n_6144),
.A2(n_6148),
.B(n_6146),
.Y(n_6764)
);

INVx2_ASAP7_75t_L g6765 ( 
.A(n_5991),
.Y(n_6765)
);

A2O1A1Ixp33_ASAP7_75t_L g6766 ( 
.A1(n_5429),
.A2(n_5019),
.B(n_5039),
.C(n_5342),
.Y(n_6766)
);

AND2x4_ASAP7_75t_L g6767 ( 
.A(n_4756),
.B(n_4782),
.Y(n_6767)
);

NAND2xp5_ASAP7_75t_L g6768 ( 
.A(n_4871),
.B(n_4882),
.Y(n_6768)
);

INVx2_ASAP7_75t_L g6769 ( 
.A(n_5991),
.Y(n_6769)
);

AOI21xp5_ASAP7_75t_L g6770 ( 
.A1(n_4971),
.A2(n_5046),
.B(n_5139),
.Y(n_6770)
);

OAI21xp5_ASAP7_75t_L g6771 ( 
.A1(n_4919),
.A2(n_4952),
.B(n_5355),
.Y(n_6771)
);

NAND2x1_ASAP7_75t_L g6772 ( 
.A(n_4924),
.B(n_5265),
.Y(n_6772)
);

OAI21x1_ASAP7_75t_L g6773 ( 
.A1(n_6148),
.A2(n_6153),
.B(n_6152),
.Y(n_6773)
);

AOI21x1_ASAP7_75t_L g6774 ( 
.A1(n_5985),
.A2(n_6153),
.B(n_6152),
.Y(n_6774)
);

INVx2_ASAP7_75t_L g6775 ( 
.A(n_5991),
.Y(n_6775)
);

BUFx6f_ASAP7_75t_L g6776 ( 
.A(n_4765),
.Y(n_6776)
);

NAND2xp33_ASAP7_75t_L g6777 ( 
.A(n_4942),
.B(n_5188),
.Y(n_6777)
);

AND2x2_ASAP7_75t_L g6778 ( 
.A(n_5405),
.B(n_5443),
.Y(n_6778)
);

NAND2xp5_ASAP7_75t_SL g6779 ( 
.A(n_5188),
.B(n_5268),
.Y(n_6779)
);

AOI21xp5_ASAP7_75t_L g6780 ( 
.A1(n_5046),
.A2(n_5139),
.B(n_5452),
.Y(n_6780)
);

NAND2xp5_ASAP7_75t_SL g6781 ( 
.A(n_5175),
.B(n_6007),
.Y(n_6781)
);

OAI21x1_ASAP7_75t_L g6782 ( 
.A1(n_6154),
.A2(n_6158),
.B(n_6156),
.Y(n_6782)
);

AND2x2_ASAP7_75t_L g6783 ( 
.A(n_5443),
.B(n_5555),
.Y(n_6783)
);

NAND2x1p5_ASAP7_75t_L g6784 ( 
.A(n_4765),
.B(n_4816),
.Y(n_6784)
);

AOI221xp5_ASAP7_75t_SL g6785 ( 
.A1(n_5061),
.A2(n_5441),
.B1(n_5427),
.B2(n_4954),
.C(n_4980),
.Y(n_6785)
);

INVx1_ASAP7_75t_L g6786 ( 
.A(n_4977),
.Y(n_6786)
);

A2O1A1Ixp33_ASAP7_75t_L g6787 ( 
.A1(n_5429),
.A2(n_5365),
.B(n_5380),
.C(n_5096),
.Y(n_6787)
);

AOI21xp5_ASAP7_75t_L g6788 ( 
.A1(n_5452),
.A2(n_5407),
.B(n_4898),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_4977),
.Y(n_6789)
);

OAI21x1_ASAP7_75t_L g6790 ( 
.A1(n_6154),
.A2(n_6158),
.B(n_6156),
.Y(n_6790)
);

OAI21x1_ASAP7_75t_L g6791 ( 
.A1(n_6166),
.A2(n_6188),
.B(n_5029),
.Y(n_6791)
);

AOI21xp5_ASAP7_75t_L g6792 ( 
.A1(n_5407),
.A2(n_6195),
.B(n_5096),
.Y(n_6792)
);

OAI21xp5_ASAP7_75t_L g6793 ( 
.A1(n_5355),
.A2(n_5351),
.B(n_4927),
.Y(n_6793)
);

OAI21xp5_ASAP7_75t_L g6794 ( 
.A1(n_4888),
.A2(n_5008),
.B(n_5007),
.Y(n_6794)
);

OAI21xp5_ASAP7_75t_L g6795 ( 
.A1(n_5013),
.A2(n_5069),
.B(n_5021),
.Y(n_6795)
);

A2O1A1Ixp33_ASAP7_75t_L g6796 ( 
.A1(n_5441),
.A2(n_5466),
.B(n_5388),
.C(n_5403),
.Y(n_6796)
);

OAI21x1_ASAP7_75t_L g6797 ( 
.A1(n_6166),
.A2(n_6188),
.B(n_5029),
.Y(n_6797)
);

NOR2xp33_ASAP7_75t_L g6798 ( 
.A(n_5447),
.B(n_5264),
.Y(n_6798)
);

INVx1_ASAP7_75t_L g6799 ( 
.A(n_4981),
.Y(n_6799)
);

AOI21xp5_ASAP7_75t_L g6800 ( 
.A1(n_6195),
.A2(n_5301),
.B(n_5298),
.Y(n_6800)
);

AOI21xp5_ASAP7_75t_L g6801 ( 
.A1(n_5301),
.A2(n_5348),
.B(n_5298),
.Y(n_6801)
);

OAI22xp5_ASAP7_75t_L g6802 ( 
.A1(n_4916),
.A2(n_4824),
.B1(n_4831),
.B2(n_4795),
.Y(n_6802)
);

NAND2xp5_ASAP7_75t_L g6803 ( 
.A(n_4882),
.B(n_4883),
.Y(n_6803)
);

AOI221xp5_ASAP7_75t_SL g6804 ( 
.A1(n_5427),
.A2(n_5500),
.B1(n_5092),
.B2(n_5179),
.C(n_5102),
.Y(n_6804)
);

OAI21xp5_ASAP7_75t_L g6805 ( 
.A1(n_5129),
.A2(n_5177),
.B(n_4873),
.Y(n_6805)
);

BUFx2_ASAP7_75t_L g6806 ( 
.A(n_5525),
.Y(n_6806)
);

AOI21xp5_ASAP7_75t_L g6807 ( 
.A1(n_5296),
.A2(n_5348),
.B(n_5324),
.Y(n_6807)
);

NAND2x1p5_ASAP7_75t_L g6808 ( 
.A(n_4765),
.B(n_4816),
.Y(n_6808)
);

AOI21xp5_ASAP7_75t_L g6809 ( 
.A1(n_5296),
.A2(n_5349),
.B(n_5324),
.Y(n_6809)
);

OAI21x1_ASAP7_75t_L g6810 ( 
.A1(n_5023),
.A2(n_5029),
.B(n_5110),
.Y(n_6810)
);

OAI21x1_ASAP7_75t_SL g6811 ( 
.A1(n_5085),
.A2(n_5093),
.B(n_5220),
.Y(n_6811)
);

OAI21xp33_ASAP7_75t_SL g6812 ( 
.A1(n_5341),
.A2(n_6100),
.B(n_6010),
.Y(n_6812)
);

OAI21xp5_ASAP7_75t_L g6813 ( 
.A1(n_5177),
.A2(n_4873),
.B(n_4840),
.Y(n_6813)
);

OAI21x1_ASAP7_75t_L g6814 ( 
.A1(n_5023),
.A2(n_5112),
.B(n_5110),
.Y(n_6814)
);

OAI21x1_ASAP7_75t_L g6815 ( 
.A1(n_5023),
.A2(n_5115),
.B(n_5112),
.Y(n_6815)
);

AND2x2_ASAP7_75t_L g6816 ( 
.A(n_5555),
.B(n_5632),
.Y(n_6816)
);

AOI21xp5_ASAP7_75t_L g6817 ( 
.A1(n_5350),
.A2(n_5326),
.B(n_5305),
.Y(n_6817)
);

AOI21xp5_ASAP7_75t_L g6818 ( 
.A1(n_5350),
.A2(n_5326),
.B(n_5305),
.Y(n_6818)
);

OAI21xp5_ASAP7_75t_L g6819 ( 
.A1(n_4840),
.A2(n_4937),
.B(n_4915),
.Y(n_6819)
);

OAI21xp5_ASAP7_75t_L g6820 ( 
.A1(n_4915),
.A2(n_4937),
.B(n_5137),
.Y(n_6820)
);

AOI21xp5_ASAP7_75t_L g6821 ( 
.A1(n_5332),
.A2(n_5354),
.B(n_5349),
.Y(n_6821)
);

NAND2xp5_ASAP7_75t_SL g6822 ( 
.A(n_6007),
.B(n_5393),
.Y(n_6822)
);

NAND2xp5_ASAP7_75t_L g6823 ( 
.A(n_4883),
.B(n_4887),
.Y(n_6823)
);

AOI21x1_ASAP7_75t_L g6824 ( 
.A1(n_5985),
.A2(n_5544),
.B(n_6189),
.Y(n_6824)
);

OR2x6_ASAP7_75t_L g6825 ( 
.A(n_5270),
.B(n_5463),
.Y(n_6825)
);

OR2x6_ASAP7_75t_L g6826 ( 
.A(n_5270),
.B(n_5463),
.Y(n_6826)
);

NAND2xp5_ASAP7_75t_L g6827 ( 
.A(n_4887),
.B(n_4895),
.Y(n_6827)
);

BUFx6f_ASAP7_75t_L g6828 ( 
.A(n_4765),
.Y(n_6828)
);

BUFx12f_ASAP7_75t_L g6829 ( 
.A(n_5259),
.Y(n_6829)
);

A2O1A1Ixp33_ASAP7_75t_L g6830 ( 
.A1(n_5386),
.A2(n_5425),
.B(n_5398),
.C(n_5655),
.Y(n_6830)
);

INVx2_ASAP7_75t_L g6831 ( 
.A(n_6005),
.Y(n_6831)
);

INVx4_ASAP7_75t_SL g6832 ( 
.A(n_5148),
.Y(n_6832)
);

NOR2xp33_ASAP7_75t_L g6833 ( 
.A(n_5447),
.B(n_5267),
.Y(n_6833)
);

NAND2xp5_ASAP7_75t_L g6834 ( 
.A(n_4895),
.B(n_4901),
.Y(n_6834)
);

OAI22x1_ASAP7_75t_L g6835 ( 
.A1(n_6032),
.A2(n_6041),
.B1(n_6061),
.B2(n_6034),
.Y(n_6835)
);

OAI21xp5_ASAP7_75t_L g6836 ( 
.A1(n_5137),
.A2(n_5211),
.B(n_5366),
.Y(n_6836)
);

AO31x2_ASAP7_75t_L g6837 ( 
.A1(n_5397),
.A2(n_5813),
.A3(n_5814),
.B(n_5809),
.Y(n_6837)
);

CKINVDCx5p33_ASAP7_75t_R g6838 ( 
.A(n_4838),
.Y(n_6838)
);

OAI21x1_ASAP7_75t_L g6839 ( 
.A1(n_5115),
.A2(n_5118),
.B(n_5116),
.Y(n_6839)
);

CKINVDCx5p33_ASAP7_75t_R g6840 ( 
.A(n_5101),
.Y(n_6840)
);

NAND2xp5_ASAP7_75t_L g6841 ( 
.A(n_4901),
.B(n_4903),
.Y(n_6841)
);

AND3x2_ASAP7_75t_L g6842 ( 
.A(n_5916),
.B(n_5215),
.C(n_5567),
.Y(n_6842)
);

INVx2_ASAP7_75t_L g6843 ( 
.A(n_6005),
.Y(n_6843)
);

NOR3xp33_ASAP7_75t_L g6844 ( 
.A(n_5457),
.B(n_5458),
.C(n_5500),
.Y(n_6844)
);

OAI21xp5_ASAP7_75t_L g6845 ( 
.A1(n_5137),
.A2(n_5367),
.B(n_5366),
.Y(n_6845)
);

OAI21xp5_ASAP7_75t_L g6846 ( 
.A1(n_5367),
.A2(n_5315),
.B(n_5245),
.Y(n_6846)
);

OAI21x1_ASAP7_75t_L g6847 ( 
.A1(n_5116),
.A2(n_5125),
.B(n_5118),
.Y(n_6847)
);

INVx1_ASAP7_75t_SL g6848 ( 
.A(n_5292),
.Y(n_6848)
);

A2O1A1Ixp33_ASAP7_75t_L g6849 ( 
.A1(n_5655),
.A2(n_5159),
.B(n_5393),
.C(n_5492),
.Y(n_6849)
);

NAND2x1p5_ASAP7_75t_L g6850 ( 
.A(n_4816),
.B(n_4846),
.Y(n_6850)
);

A2O1A1Ixp33_ASAP7_75t_L g6851 ( 
.A1(n_5583),
.A2(n_6063),
.B(n_5131),
.C(n_4841),
.Y(n_6851)
);

NAND2x1p5_ASAP7_75t_L g6852 ( 
.A(n_4816),
.B(n_4846),
.Y(n_6852)
);

OAI21x1_ASAP7_75t_L g6853 ( 
.A1(n_5128),
.A2(n_5284),
.B(n_5281),
.Y(n_6853)
);

OAI21x1_ASAP7_75t_L g6854 ( 
.A1(n_5281),
.A2(n_5294),
.B(n_5284),
.Y(n_6854)
);

AOI21xp33_ASAP7_75t_L g6855 ( 
.A1(n_5341),
.A2(n_5295),
.B(n_5227),
.Y(n_6855)
);

NAND3xp33_ASAP7_75t_SL g6856 ( 
.A(n_5369),
.B(n_5675),
.C(n_4839),
.Y(n_6856)
);

OAI21xp5_ASAP7_75t_L g6857 ( 
.A1(n_5315),
.A2(n_5160),
.B(n_5341),
.Y(n_6857)
);

AOI21x1_ASAP7_75t_L g6858 ( 
.A1(n_5544),
.A2(n_6191),
.B(n_6189),
.Y(n_6858)
);

CKINVDCx5p33_ASAP7_75t_R g6859 ( 
.A(n_4739),
.Y(n_6859)
);

AND2x2_ASAP7_75t_L g6860 ( 
.A(n_5555),
.B(n_5632),
.Y(n_6860)
);

OAI22x1_ASAP7_75t_L g6861 ( 
.A1(n_6061),
.A2(n_5247),
.B1(n_5086),
.B2(n_5523),
.Y(n_6861)
);

NAND3x1_ASAP7_75t_L g6862 ( 
.A(n_5086),
.B(n_5523),
.C(n_5738),
.Y(n_6862)
);

NAND2xp5_ASAP7_75t_L g6863 ( 
.A(n_4903),
.B(n_4909),
.Y(n_6863)
);

AND2x2_ASAP7_75t_L g6864 ( 
.A(n_5632),
.B(n_5470),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_4981),
.Y(n_6865)
);

OAI21x1_ASAP7_75t_L g6866 ( 
.A1(n_5281),
.A2(n_5294),
.B(n_5284),
.Y(n_6866)
);

BUFx4f_ASAP7_75t_SL g6867 ( 
.A(n_4739),
.Y(n_6867)
);

INVx2_ASAP7_75t_L g6868 ( 
.A(n_6005),
.Y(n_6868)
);

NAND2xp5_ASAP7_75t_L g6869 ( 
.A(n_4909),
.B(n_4921),
.Y(n_6869)
);

OAI21x1_ASAP7_75t_L g6870 ( 
.A1(n_5294),
.A2(n_5603),
.B(n_5519),
.Y(n_6870)
);

OAI21xp5_ASAP7_75t_L g6871 ( 
.A1(n_5220),
.A2(n_5273),
.B(n_5227),
.Y(n_6871)
);

AOI211x1_ASAP7_75t_L g6872 ( 
.A1(n_5092),
.A2(n_5130),
.B(n_5194),
.C(n_5113),
.Y(n_6872)
);

OAI22xp33_ASAP7_75t_L g6873 ( 
.A1(n_4839),
.A2(n_5295),
.B1(n_5107),
.B2(n_5119),
.Y(n_6873)
);

AOI21xp5_ASAP7_75t_L g6874 ( 
.A1(n_6219),
.A2(n_6225),
.B(n_5479),
.Y(n_6874)
);

AOI21x1_ASAP7_75t_L g6875 ( 
.A1(n_6191),
.A2(n_5813),
.B(n_5809),
.Y(n_6875)
);

NAND2xp5_ASAP7_75t_L g6876 ( 
.A(n_4921),
.B(n_4929),
.Y(n_6876)
);

AOI21xp5_ASAP7_75t_L g6877 ( 
.A1(n_6219),
.A2(n_6225),
.B(n_5479),
.Y(n_6877)
);

NAND2xp5_ASAP7_75t_L g6878 ( 
.A(n_4929),
.B(n_4932),
.Y(n_6878)
);

AOI21xp5_ASAP7_75t_SL g6879 ( 
.A1(n_5176),
.A2(n_5490),
.B(n_5902),
.Y(n_6879)
);

NAND2xp5_ASAP7_75t_L g6880 ( 
.A(n_4932),
.B(n_4944),
.Y(n_6880)
);

AOI21xp33_ASAP7_75t_L g6881 ( 
.A1(n_5295),
.A2(n_5338),
.B(n_5273),
.Y(n_6881)
);

HB1xp67_ASAP7_75t_L g6882 ( 
.A(n_6026),
.Y(n_6882)
);

OAI21xp5_ASAP7_75t_L g6883 ( 
.A1(n_5338),
.A2(n_4876),
.B(n_4854),
.Y(n_6883)
);

AOI21xp5_ASAP7_75t_SL g6884 ( 
.A1(n_5922),
.A2(n_5952),
.B(n_5944),
.Y(n_6884)
);

OAI21x1_ASAP7_75t_L g6885 ( 
.A1(n_5519),
.A2(n_5718),
.B(n_5603),
.Y(n_6885)
);

AOI21xp33_ASAP7_75t_L g6886 ( 
.A1(n_5295),
.A2(n_5181),
.B(n_5198),
.Y(n_6886)
);

INVx2_ASAP7_75t_SL g6887 ( 
.A(n_5439),
.Y(n_6887)
);

AOI22xp5_ASAP7_75t_L g6888 ( 
.A1(n_5369),
.A2(n_4884),
.B1(n_4904),
.B2(n_4896),
.Y(n_6888)
);

O2A1O1Ixp5_ASAP7_75t_L g6889 ( 
.A1(n_5198),
.A2(n_5102),
.B(n_5097),
.C(n_5532),
.Y(n_6889)
);

NAND2xp5_ASAP7_75t_L g6890 ( 
.A(n_4944),
.B(n_4951),
.Y(n_6890)
);

A2O1A1Ixp33_ASAP7_75t_L g6891 ( 
.A1(n_6063),
.A2(n_4950),
.B(n_4975),
.C(n_4961),
.Y(n_6891)
);

BUFx2_ASAP7_75t_L g6892 ( 
.A(n_5525),
.Y(n_6892)
);

OAI21x1_ASAP7_75t_L g6893 ( 
.A1(n_5519),
.A2(n_5718),
.B(n_5603),
.Y(n_6893)
);

OAI21xp5_ASAP7_75t_L g6894 ( 
.A1(n_5002),
.A2(n_5097),
.B(n_5196),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_4984),
.Y(n_6895)
);

A2O1A1Ixp33_ASAP7_75t_L g6896 ( 
.A1(n_5158),
.A2(n_5165),
.B(n_5167),
.C(n_5166),
.Y(n_6896)
);

AO31x2_ASAP7_75t_L g6897 ( 
.A1(n_5397),
.A2(n_5818),
.A3(n_5821),
.B(n_5814),
.Y(n_6897)
);

OAI21x1_ASAP7_75t_L g6898 ( 
.A1(n_5718),
.A2(n_6027),
.B(n_5779),
.Y(n_6898)
);

OR2x6_ASAP7_75t_L g6899 ( 
.A(n_5270),
.B(n_5463),
.Y(n_6899)
);

INVx2_ASAP7_75t_L g6900 ( 
.A(n_6009),
.Y(n_6900)
);

NAND2xp5_ASAP7_75t_L g6901 ( 
.A(n_4951),
.B(n_4957),
.Y(n_6901)
);

AND2x2_ASAP7_75t_L g6902 ( 
.A(n_5470),
.B(n_5483),
.Y(n_6902)
);

OAI21x1_ASAP7_75t_L g6903 ( 
.A1(n_5779),
.A2(n_6092),
.B(n_6027),
.Y(n_6903)
);

NAND2xp5_ASAP7_75t_L g6904 ( 
.A(n_4957),
.B(n_4959),
.Y(n_6904)
);

INVx2_ASAP7_75t_L g6905 ( 
.A(n_6009),
.Y(n_6905)
);

INVx1_ASAP7_75t_L g6906 ( 
.A(n_4984),
.Y(n_6906)
);

NAND2xp5_ASAP7_75t_L g6907 ( 
.A(n_4959),
.B(n_4966),
.Y(n_6907)
);

A2O1A1Ixp33_ASAP7_75t_L g6908 ( 
.A1(n_5158),
.A2(n_5165),
.B(n_5167),
.C(n_5166),
.Y(n_6908)
);

BUFx12f_ASAP7_75t_L g6909 ( 
.A(n_5259),
.Y(n_6909)
);

OAI21xp5_ASAP7_75t_L g6910 ( 
.A1(n_5196),
.A2(n_5646),
.B(n_5146),
.Y(n_6910)
);

AOI21xp5_ASAP7_75t_L g6911 ( 
.A1(n_6215),
.A2(n_6039),
.B(n_6150),
.Y(n_6911)
);

AOI21xp5_ASAP7_75t_L g6912 ( 
.A1(n_6215),
.A2(n_6039),
.B(n_6150),
.Y(n_6912)
);

NAND2xp5_ASAP7_75t_SL g6913 ( 
.A(n_5247),
.B(n_5362),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_4986),
.Y(n_6914)
);

AOI21xp5_ASAP7_75t_L g6915 ( 
.A1(n_5439),
.A2(n_5705),
.B(n_5626),
.Y(n_6915)
);

INVx2_ASAP7_75t_SL g6916 ( 
.A(n_5626),
.Y(n_6916)
);

OR2x2_ASAP7_75t_L g6917 ( 
.A(n_5465),
.B(n_5467),
.Y(n_6917)
);

AOI21xp5_ASAP7_75t_L g6918 ( 
.A1(n_5626),
.A2(n_5808),
.B(n_5705),
.Y(n_6918)
);

NAND2x1p5_ASAP7_75t_L g6919 ( 
.A(n_4816),
.B(n_4846),
.Y(n_6919)
);

INVx1_ASAP7_75t_SL g6920 ( 
.A(n_5292),
.Y(n_6920)
);

INVx1_ASAP7_75t_L g6921 ( 
.A(n_4986),
.Y(n_6921)
);

AOI21xp5_ASAP7_75t_L g6922 ( 
.A1(n_5626),
.A2(n_5808),
.B(n_5705),
.Y(n_6922)
);

NOR2xp67_ASAP7_75t_L g6923 ( 
.A(n_5051),
.B(n_5075),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_5051),
.Y(n_6924)
);

OAI21xp5_ASAP7_75t_L g6925 ( 
.A1(n_5646),
.A2(n_5146),
.B(n_5181),
.Y(n_6925)
);

OAI22x1_ASAP7_75t_L g6926 ( 
.A1(n_5087),
.A2(n_5161),
.B1(n_5207),
.B2(n_5819),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_5075),
.Y(n_6927)
);

NOR2xp33_ASAP7_75t_R g6928 ( 
.A(n_5050),
.B(n_5607),
.Y(n_6928)
);

AND3x4_ASAP7_75t_L g6929 ( 
.A(n_5846),
.B(n_5909),
.C(n_5531),
.Y(n_6929)
);

INVx2_ASAP7_75t_L g6930 ( 
.A(n_6009),
.Y(n_6930)
);

OAI21x1_ASAP7_75t_L g6931 ( 
.A1(n_5779),
.A2(n_6092),
.B(n_6027),
.Y(n_6931)
);

AOI21xp5_ASAP7_75t_L g6932 ( 
.A1(n_5626),
.A2(n_5808),
.B(n_5705),
.Y(n_6932)
);

OAI21x1_ASAP7_75t_L g6933 ( 
.A1(n_6092),
.A2(n_5105),
.B(n_5824),
.Y(n_6933)
);

BUFx2_ASAP7_75t_L g6934 ( 
.A(n_5879),
.Y(n_6934)
);

HB1xp67_ASAP7_75t_SL g6935 ( 
.A(n_5514),
.Y(n_6935)
);

OAI22x1_ASAP7_75t_L g6936 ( 
.A1(n_5087),
.A2(n_5161),
.B1(n_5207),
.B2(n_5819),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_5147),
.Y(n_6937)
);

BUFx6f_ASAP7_75t_L g6938 ( 
.A(n_4816),
.Y(n_6938)
);

AOI21xp33_ASAP7_75t_L g6939 ( 
.A1(n_5179),
.A2(n_5645),
.B(n_5461),
.Y(n_6939)
);

AOI21xp5_ASAP7_75t_L g6940 ( 
.A1(n_5626),
.A2(n_5808),
.B(n_5705),
.Y(n_6940)
);

AND2x2_ASAP7_75t_L g6941 ( 
.A(n_5470),
.B(n_5483),
.Y(n_6941)
);

INVxp67_ASAP7_75t_L g6942 ( 
.A(n_5311),
.Y(n_6942)
);

NAND2xp5_ASAP7_75t_L g6943 ( 
.A(n_4966),
.B(n_4967),
.Y(n_6943)
);

AOI21xp5_ASAP7_75t_L g6944 ( 
.A1(n_5626),
.A2(n_5808),
.B(n_5705),
.Y(n_6944)
);

AOI21xp5_ASAP7_75t_L g6945 ( 
.A1(n_5705),
.A2(n_5808),
.B(n_6199),
.Y(n_6945)
);

NAND2xp5_ASAP7_75t_L g6946 ( 
.A(n_4967),
.B(n_4969),
.Y(n_6946)
);

NAND2xp5_ASAP7_75t_L g6947 ( 
.A(n_4969),
.B(n_4973),
.Y(n_6947)
);

NAND2xp5_ASAP7_75t_SL g6948 ( 
.A(n_5362),
.B(n_5378),
.Y(n_6948)
);

OAI22xp5_ASAP7_75t_L g6949 ( 
.A1(n_5098),
.A2(n_5119),
.B1(n_5126),
.B2(n_5107),
.Y(n_6949)
);

OAI21x1_ASAP7_75t_L g6950 ( 
.A1(n_5105),
.A2(n_5872),
.B(n_5870),
.Y(n_6950)
);

O2A1O1Ixp5_ASAP7_75t_L g6951 ( 
.A1(n_5532),
.A2(n_5540),
.B(n_5618),
.C(n_5592),
.Y(n_6951)
);

NAND2x2_ASAP7_75t_L g6952 ( 
.A(n_5846),
.B(n_5909),
.Y(n_6952)
);

INVx1_ASAP7_75t_L g6953 ( 
.A(n_5147),
.Y(n_6953)
);

OAI21x1_ASAP7_75t_L g6954 ( 
.A1(n_5105),
.A2(n_5905),
.B(n_5888),
.Y(n_6954)
);

AO31x2_ASAP7_75t_L g6955 ( 
.A1(n_5905),
.A2(n_5937),
.A3(n_5939),
.B(n_5912),
.Y(n_6955)
);

NAND2xp5_ASAP7_75t_SL g6956 ( 
.A(n_5378),
.B(n_5387),
.Y(n_6956)
);

OAI21x1_ASAP7_75t_L g6957 ( 
.A1(n_5912),
.A2(n_5939),
.B(n_5937),
.Y(n_6957)
);

OAI21xp5_ASAP7_75t_L g6958 ( 
.A1(n_5733),
.A2(n_5516),
.B(n_5493),
.Y(n_6958)
);

OAI21x1_ASAP7_75t_L g6959 ( 
.A1(n_5947),
.A2(n_5955),
.B(n_5949),
.Y(n_6959)
);

BUFx6f_ASAP7_75t_L g6960 ( 
.A(n_4816),
.Y(n_6960)
);

OAI21x1_ASAP7_75t_L g6961 ( 
.A1(n_5947),
.A2(n_5955),
.B(n_5949),
.Y(n_6961)
);

AOI221xp5_ASAP7_75t_L g6962 ( 
.A1(n_5530),
.A2(n_5183),
.B1(n_5391),
.B2(n_5420),
.C(n_5387),
.Y(n_6962)
);

INVx1_ASAP7_75t_L g6963 ( 
.A(n_5153),
.Y(n_6963)
);

INVx2_ASAP7_75t_L g6964 ( 
.A(n_6018),
.Y(n_6964)
);

OAI22xp33_ASAP7_75t_L g6965 ( 
.A1(n_5098),
.A2(n_5126),
.B1(n_5132),
.B2(n_5053),
.Y(n_6965)
);

AO21x1_ASAP7_75t_L g6966 ( 
.A1(n_5890),
.A2(n_5900),
.B(n_5446),
.Y(n_6966)
);

AOI21xp5_ASAP7_75t_L g6967 ( 
.A1(n_6204),
.A2(n_6200),
.B(n_5293),
.Y(n_6967)
);

OAI21xp5_ASAP7_75t_L g6968 ( 
.A1(n_5733),
.A2(n_5675),
.B(n_5528),
.Y(n_6968)
);

BUFx6f_ASAP7_75t_L g6969 ( 
.A(n_4846),
.Y(n_6969)
);

INVx6_ASAP7_75t_SL g6970 ( 
.A(n_5251),
.Y(n_6970)
);

NOR2xp33_ASAP7_75t_L g6971 ( 
.A(n_4973),
.B(n_4976),
.Y(n_6971)
);

INVx1_ASAP7_75t_L g6972 ( 
.A(n_5153),
.Y(n_6972)
);

INVx2_ASAP7_75t_L g6973 ( 
.A(n_6018),
.Y(n_6973)
);

OAI21x1_ASAP7_75t_L g6974 ( 
.A1(n_5962),
.A2(n_5981),
.B(n_5977),
.Y(n_6974)
);

AOI21xp5_ASAP7_75t_L g6975 ( 
.A1(n_6204),
.A2(n_5293),
.B(n_5391),
.Y(n_6975)
);

OAI21x1_ASAP7_75t_L g6976 ( 
.A1(n_5962),
.A2(n_5981),
.B(n_5977),
.Y(n_6976)
);

AOI21xp5_ASAP7_75t_L g6977 ( 
.A1(n_5420),
.A2(n_5422),
.B(n_4997),
.Y(n_6977)
);

OAI22xp5_ASAP7_75t_L g6978 ( 
.A1(n_5132),
.A2(n_5275),
.B1(n_5134),
.B2(n_5174),
.Y(n_6978)
);

BUFx2_ASAP7_75t_L g6979 ( 
.A(n_5879),
.Y(n_6979)
);

NAND2xp33_ASAP7_75t_SL g6980 ( 
.A(n_5321),
.B(n_6214),
.Y(n_6980)
);

AOI21xp5_ASAP7_75t_SL g6981 ( 
.A1(n_6040),
.A2(n_6053),
.B(n_6023),
.Y(n_6981)
);

OAI21xp5_ASAP7_75t_L g6982 ( 
.A1(n_5528),
.A2(n_5645),
.B(n_5120),
.Y(n_6982)
);

INVx1_ASAP7_75t_L g6983 ( 
.A(n_5180),
.Y(n_6983)
);

AOI22xp5_ASAP7_75t_L g6984 ( 
.A1(n_5448),
.A2(n_5518),
.B1(n_5517),
.B2(n_5530),
.Y(n_6984)
);

BUFx3_ASAP7_75t_L g6985 ( 
.A(n_5573),
.Y(n_6985)
);

NAND2xp5_ASAP7_75t_L g6986 ( 
.A(n_4976),
.B(n_4997),
.Y(n_6986)
);

NAND2xp5_ASAP7_75t_L g6987 ( 
.A(n_5003),
.B(n_5004),
.Y(n_6987)
);

NAND2xp5_ASAP7_75t_L g6988 ( 
.A(n_5003),
.B(n_5004),
.Y(n_6988)
);

NOR2xp33_ASAP7_75t_SL g6989 ( 
.A(n_4761),
.B(n_5756),
.Y(n_6989)
);

A2O1A1Ixp33_ASAP7_75t_L g6990 ( 
.A1(n_5186),
.A2(n_5190),
.B(n_5187),
.C(n_5283),
.Y(n_6990)
);

AOI21xp5_ASAP7_75t_SL g6991 ( 
.A1(n_6023),
.A2(n_5966),
.B(n_6192),
.Y(n_6991)
);

OAI21x1_ASAP7_75t_L g6992 ( 
.A1(n_5984),
.A2(n_6004),
.B(n_5996),
.Y(n_6992)
);

NOR2xp33_ASAP7_75t_L g6993 ( 
.A(n_5009),
.B(n_5016),
.Y(n_6993)
);

AND2x2_ASAP7_75t_L g6994 ( 
.A(n_5483),
.B(n_5510),
.Y(n_6994)
);

AO21x2_ASAP7_75t_L g6995 ( 
.A1(n_5900),
.A2(n_5996),
.B(n_5984),
.Y(n_6995)
);

AOI21xp5_ASAP7_75t_L g6996 ( 
.A1(n_5422),
.A2(n_5016),
.B(n_5009),
.Y(n_6996)
);

AO31x2_ASAP7_75t_L g6997 ( 
.A1(n_6004),
.A2(n_6015),
.A3(n_6017),
.B(n_6012),
.Y(n_6997)
);

AOI21xp5_ASAP7_75t_L g6998 ( 
.A1(n_5018),
.A2(n_5032),
.B(n_5030),
.Y(n_6998)
);

AOI21xp5_ASAP7_75t_L g6999 ( 
.A1(n_5018),
.A2(n_5032),
.B(n_5030),
.Y(n_6999)
);

OAI21x1_ASAP7_75t_L g7000 ( 
.A1(n_6012),
.A2(n_6017),
.B(n_6015),
.Y(n_7000)
);

OAI21x1_ASAP7_75t_L g7001 ( 
.A1(n_6019),
.A2(n_6024),
.B(n_6021),
.Y(n_7001)
);

OAI21x1_ASAP7_75t_L g7002 ( 
.A1(n_6019),
.A2(n_6024),
.B(n_6021),
.Y(n_7002)
);

OAI21x1_ASAP7_75t_L g7003 ( 
.A1(n_6030),
.A2(n_6033),
.B(n_6031),
.Y(n_7003)
);

AOI21x1_ASAP7_75t_L g7004 ( 
.A1(n_6030),
.A2(n_6033),
.B(n_6031),
.Y(n_7004)
);

OAI21xp5_ASAP7_75t_L g7005 ( 
.A1(n_5229),
.A2(n_5684),
.B(n_5130),
.Y(n_7005)
);

AOI21x1_ASAP7_75t_L g7006 ( 
.A1(n_6045),
.A2(n_6050),
.B(n_6047),
.Y(n_7006)
);

OAI21x1_ASAP7_75t_L g7007 ( 
.A1(n_6045),
.A2(n_6050),
.B(n_6047),
.Y(n_7007)
);

OAI21x1_ASAP7_75t_L g7008 ( 
.A1(n_6054),
.A2(n_6067),
.B(n_6057),
.Y(n_7008)
);

NAND2xp5_ASAP7_75t_L g7009 ( 
.A(n_5038),
.B(n_5043),
.Y(n_7009)
);

AOI21xp5_ASAP7_75t_L g7010 ( 
.A1(n_5038),
.A2(n_5043),
.B(n_6008),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_5180),
.Y(n_7011)
);

AND2x4_ASAP7_75t_L g7012 ( 
.A(n_4756),
.B(n_4782),
.Y(n_7012)
);

NOR2xp33_ASAP7_75t_SL g7013 ( 
.A(n_4761),
.B(n_5215),
.Y(n_7013)
);

AOI21xp5_ASAP7_75t_L g7014 ( 
.A1(n_6008),
.A2(n_5488),
.B(n_6054),
.Y(n_7014)
);

NAND2xp5_ASAP7_75t_L g7015 ( 
.A(n_5203),
.B(n_5212),
.Y(n_7015)
);

BUFx3_ASAP7_75t_L g7016 ( 
.A(n_5722),
.Y(n_7016)
);

NAND2xp5_ASAP7_75t_L g7017 ( 
.A(n_5203),
.B(n_5212),
.Y(n_7017)
);

NAND2xp5_ASAP7_75t_L g7018 ( 
.A(n_5216),
.B(n_5217),
.Y(n_7018)
);

NAND2xp5_ASAP7_75t_L g7019 ( 
.A(n_5216),
.B(n_5217),
.Y(n_7019)
);

INVx5_ASAP7_75t_L g7020 ( 
.A(n_4846),
.Y(n_7020)
);

OAI21x1_ASAP7_75t_L g7021 ( 
.A1(n_6057),
.A2(n_6077),
.B(n_6067),
.Y(n_7021)
);

INVxp67_ASAP7_75t_L g7022 ( 
.A(n_5311),
.Y(n_7022)
);

NAND2x1p5_ASAP7_75t_L g7023 ( 
.A(n_4846),
.B(n_4907),
.Y(n_7023)
);

AOI21xp5_ASAP7_75t_L g7024 ( 
.A1(n_6077),
.A2(n_6097),
.B(n_6094),
.Y(n_7024)
);

NAND2xp5_ASAP7_75t_L g7025 ( 
.A(n_5228),
.B(n_5241),
.Y(n_7025)
);

AOI21xp5_ASAP7_75t_L g7026 ( 
.A1(n_6094),
.A2(n_6099),
.B(n_6097),
.Y(n_7026)
);

AND2x2_ASAP7_75t_L g7027 ( 
.A(n_5510),
.B(n_5520),
.Y(n_7027)
);

CKINVDCx5p33_ASAP7_75t_R g7028 ( 
.A(n_4739),
.Y(n_7028)
);

AND2x4_ASAP7_75t_L g7029 ( 
.A(n_4782),
.B(n_4783),
.Y(n_7029)
);

OAI21x1_ASAP7_75t_L g7030 ( 
.A1(n_6099),
.A2(n_6103),
.B(n_5099),
.Y(n_7030)
);

OAI21xp5_ASAP7_75t_L g7031 ( 
.A1(n_5684),
.A2(n_5194),
.B(n_5113),
.Y(n_7031)
);

NAND2xp5_ASAP7_75t_L g7032 ( 
.A(n_5228),
.B(n_5241),
.Y(n_7032)
);

INVx4_ASAP7_75t_L g7033 ( 
.A(n_5463),
.Y(n_7033)
);

OAI21x1_ASAP7_75t_L g7034 ( 
.A1(n_6103),
.A2(n_5099),
.B(n_5084),
.Y(n_7034)
);

O2A1O1Ixp5_ASAP7_75t_L g7035 ( 
.A1(n_5540),
.A2(n_5592),
.B(n_5618),
.C(n_5658),
.Y(n_7035)
);

BUFx2_ASAP7_75t_L g7036 ( 
.A(n_5879),
.Y(n_7036)
);

NAND2xp5_ASAP7_75t_L g7037 ( 
.A(n_5472),
.B(n_5473),
.Y(n_7037)
);

AOI21x1_ASAP7_75t_L g7038 ( 
.A1(n_5317),
.A2(n_5323),
.B(n_5906),
.Y(n_7038)
);

AND3x4_ASAP7_75t_L g7039 ( 
.A(n_5846),
.B(n_5909),
.C(n_5531),
.Y(n_7039)
);

A2O1A1Ixp33_ASAP7_75t_L g7040 ( 
.A1(n_5595),
.A2(n_5717),
.B(n_5663),
.C(n_5829),
.Y(n_7040)
);

OAI21x1_ASAP7_75t_SL g7041 ( 
.A1(n_6209),
.A2(n_6243),
.B(n_5487),
.Y(n_7041)
);

AND2x2_ASAP7_75t_L g7042 ( 
.A(n_5510),
.B(n_5520),
.Y(n_7042)
);

OAI21x1_ASAP7_75t_L g7043 ( 
.A1(n_5084),
.A2(n_5136),
.B(n_5099),
.Y(n_7043)
);

OAI21xp5_ASAP7_75t_L g7044 ( 
.A1(n_5316),
.A2(n_5347),
.B(n_5652),
.Y(n_7044)
);

BUFx12f_ASAP7_75t_L g7045 ( 
.A(n_5082),
.Y(n_7045)
);

BUFx2_ASAP7_75t_L g7046 ( 
.A(n_5879),
.Y(n_7046)
);

AOI21x1_ASAP7_75t_L g7047 ( 
.A1(n_5317),
.A2(n_5323),
.B(n_5906),
.Y(n_7047)
);

AOI21xp5_ASAP7_75t_L g7048 ( 
.A1(n_6239),
.A2(n_6244),
.B(n_5515),
.Y(n_7048)
);

INVx1_ASAP7_75t_L g7049 ( 
.A(n_5200),
.Y(n_7049)
);

NAND2xp5_ASAP7_75t_L g7050 ( 
.A(n_5472),
.B(n_5473),
.Y(n_7050)
);

HB1xp67_ASAP7_75t_L g7051 ( 
.A(n_6026),
.Y(n_7051)
);

AO31x2_ASAP7_75t_L g7052 ( 
.A1(n_6248),
.A2(n_6072),
.A3(n_6142),
.B(n_6126),
.Y(n_7052)
);

INVx2_ASAP7_75t_L g7053 ( 
.A(n_6078),
.Y(n_7053)
);

AOI21xp5_ASAP7_75t_L g7054 ( 
.A1(n_5576),
.A2(n_5964),
.B(n_5290),
.Y(n_7054)
);

NOR2x1_ASAP7_75t_SL g7055 ( 
.A(n_5291),
.B(n_5251),
.Y(n_7055)
);

AOI21xp5_ASAP7_75t_L g7056 ( 
.A1(n_5576),
.A2(n_5964),
.B(n_5306),
.Y(n_7056)
);

NAND2xp5_ASAP7_75t_SL g7057 ( 
.A(n_5628),
.B(n_5933),
.Y(n_7057)
);

AOI21xp5_ASAP7_75t_L g7058 ( 
.A1(n_5576),
.A2(n_5964),
.B(n_5333),
.Y(n_7058)
);

NAND3xp33_ASAP7_75t_SL g7059 ( 
.A(n_5053),
.B(n_5956),
.C(n_5918),
.Y(n_7059)
);

NAND2xp5_ASAP7_75t_L g7060 ( 
.A(n_5474),
.B(n_5497),
.Y(n_7060)
);

OAI21x1_ASAP7_75t_L g7061 ( 
.A1(n_5084),
.A2(n_5136),
.B(n_5099),
.Y(n_7061)
);

INVx1_ASAP7_75t_SL g7062 ( 
.A(n_5757),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_5205),
.Y(n_7063)
);

NAND2xp5_ASAP7_75t_L g7064 ( 
.A(n_5474),
.B(n_5497),
.Y(n_7064)
);

AND3x4_ASAP7_75t_L g7065 ( 
.A(n_5628),
.B(n_5064),
.C(n_5647),
.Y(n_7065)
);

NOR2x1_ASAP7_75t_SL g7066 ( 
.A(n_5291),
.B(n_5251),
.Y(n_7066)
);

AOI21xp5_ASAP7_75t_L g7067 ( 
.A1(n_5576),
.A2(n_5964),
.B(n_5344),
.Y(n_7067)
);

CKINVDCx20_ASAP7_75t_R g7068 ( 
.A(n_6235),
.Y(n_7068)
);

OAI21x1_ASAP7_75t_L g7069 ( 
.A1(n_5084),
.A2(n_5136),
.B(n_6151),
.Y(n_7069)
);

NAND2xp5_ASAP7_75t_L g7070 ( 
.A(n_5503),
.B(n_5504),
.Y(n_7070)
);

INVx1_ASAP7_75t_L g7071 ( 
.A(n_5214),
.Y(n_7071)
);

INVxp67_ASAP7_75t_L g7072 ( 
.A(n_5151),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_5214),
.Y(n_7073)
);

NAND2xp5_ASAP7_75t_L g7074 ( 
.A(n_5503),
.B(n_5504),
.Y(n_7074)
);

OAI21x1_ASAP7_75t_L g7075 ( 
.A1(n_5136),
.A2(n_6151),
.B(n_5658),
.Y(n_7075)
);

AOI21xp5_ASAP7_75t_SL g7076 ( 
.A1(n_5883),
.A2(n_6080),
.B(n_6066),
.Y(n_7076)
);

NAND2xp5_ASAP7_75t_L g7077 ( 
.A(n_5506),
.B(n_5507),
.Y(n_7077)
);

AOI22x1_ASAP7_75t_L g7078 ( 
.A1(n_5647),
.A2(n_5304),
.B1(n_5438),
.B2(n_4762),
.Y(n_7078)
);

OAI21x1_ASAP7_75t_L g7079 ( 
.A1(n_6155),
.A2(n_6029),
.B(n_5967),
.Y(n_7079)
);

NAND2xp5_ASAP7_75t_L g7080 ( 
.A(n_5506),
.B(n_5507),
.Y(n_7080)
);

OAI21x1_ASAP7_75t_L g7081 ( 
.A1(n_6155),
.A2(n_6029),
.B(n_5967),
.Y(n_7081)
);

AOI21xp5_ASAP7_75t_L g7082 ( 
.A1(n_5279),
.A2(n_5400),
.B(n_5345),
.Y(n_7082)
);

AOI21xp33_ASAP7_75t_L g7083 ( 
.A1(n_5663),
.A2(n_5841),
.B(n_5741),
.Y(n_7083)
);

NAND2x1p5_ASAP7_75t_L g7084 ( 
.A(n_4846),
.B(n_4907),
.Y(n_7084)
);

NAND2xp5_ASAP7_75t_L g7085 ( 
.A(n_5509),
.B(n_5522),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_5509),
.B(n_5522),
.Y(n_7086)
);

AOI21xp5_ASAP7_75t_L g7087 ( 
.A1(n_5412),
.A2(n_6242),
.B(n_6228),
.Y(n_7087)
);

O2A1O1Ixp5_ASAP7_75t_L g7088 ( 
.A1(n_5698),
.A2(n_5700),
.B(n_5727),
.C(n_5837),
.Y(n_7088)
);

NAND2xp5_ASAP7_75t_L g7089 ( 
.A(n_5534),
.B(n_5543),
.Y(n_7089)
);

INVx2_ASAP7_75t_SL g7090 ( 
.A(n_5990),
.Y(n_7090)
);

NOR2xp33_ASAP7_75t_L g7091 ( 
.A(n_5135),
.B(n_5150),
.Y(n_7091)
);

AO31x2_ASAP7_75t_L g7092 ( 
.A1(n_6072),
.A2(n_6126),
.A3(n_6159),
.B(n_6142),
.Y(n_7092)
);

CKINVDCx5p33_ASAP7_75t_R g7093 ( 
.A(n_5082),
.Y(n_7093)
);

OAI21xp5_ASAP7_75t_L g7094 ( 
.A1(n_5704),
.A2(n_5746),
.B(n_5741),
.Y(n_7094)
);

AOI21x1_ASAP7_75t_L g7095 ( 
.A1(n_5551),
.A2(n_5064),
.B(n_5236),
.Y(n_7095)
);

OAI21x1_ASAP7_75t_L g7096 ( 
.A1(n_5867),
.A2(n_5697),
.B(n_5696),
.Y(n_7096)
);

OAI22xp5_ASAP7_75t_L g7097 ( 
.A1(n_5134),
.A2(n_5237),
.B1(n_5438),
.B2(n_5142),
.Y(n_7097)
);

A2O1A1Ixp33_ASAP7_75t_L g7098 ( 
.A1(n_5595),
.A2(n_5717),
.B(n_6129),
.C(n_5578),
.Y(n_7098)
);

OAI21x1_ASAP7_75t_L g7099 ( 
.A1(n_5867),
.A2(n_5760),
.B(n_5759),
.Y(n_7099)
);

NAND2xp5_ASAP7_75t_SL g7100 ( 
.A(n_5956),
.B(n_5854),
.Y(n_7100)
);

NAND2xp5_ASAP7_75t_L g7101 ( 
.A(n_5534),
.B(n_5543),
.Y(n_7101)
);

INVx1_ASAP7_75t_L g7102 ( 
.A(n_5240),
.Y(n_7102)
);

AOI21x1_ASAP7_75t_SL g7103 ( 
.A1(n_5445),
.A2(n_5893),
.B(n_5891),
.Y(n_7103)
);

OAI21x1_ASAP7_75t_L g7104 ( 
.A1(n_5867),
.A2(n_5760),
.B(n_5759),
.Y(n_7104)
);

AND2x2_ASAP7_75t_L g7105 ( 
.A(n_5520),
.B(n_4783),
.Y(n_7105)
);

NAND2xp5_ASAP7_75t_SL g7106 ( 
.A(n_5854),
.B(n_5930),
.Y(n_7106)
);

BUFx6f_ASAP7_75t_L g7107 ( 
.A(n_4907),
.Y(n_7107)
);

OAI21xp5_ASAP7_75t_SL g7108 ( 
.A1(n_5607),
.A2(n_5406),
.B(n_5313),
.Y(n_7108)
);

OAI21xp5_ASAP7_75t_L g7109 ( 
.A1(n_5704),
.A2(n_5767),
.B(n_5746),
.Y(n_7109)
);

OAI21xp5_ASAP7_75t_L g7110 ( 
.A1(n_5767),
.A2(n_5784),
.B(n_5801),
.Y(n_7110)
);

OAI21xp5_ASAP7_75t_L g7111 ( 
.A1(n_5784),
.A2(n_5801),
.B(n_5935),
.Y(n_7111)
);

OAI21x1_ASAP7_75t_L g7112 ( 
.A1(n_5764),
.A2(n_5833),
.B(n_5807),
.Y(n_7112)
);

NAND2xp5_ASAP7_75t_L g7113 ( 
.A(n_5545),
.B(n_5556),
.Y(n_7113)
);

OAI21x1_ASAP7_75t_L g7114 ( 
.A1(n_5764),
.A2(n_5833),
.B(n_5807),
.Y(n_7114)
);

INVx1_ASAP7_75t_L g7115 ( 
.A(n_5240),
.Y(n_7115)
);

AO31x2_ASAP7_75t_L g7116 ( 
.A1(n_6159),
.A2(n_6162),
.A3(n_6044),
.B(n_5312),
.Y(n_7116)
);

OAI21xp5_ASAP7_75t_L g7117 ( 
.A1(n_5841),
.A2(n_5487),
.B(n_5475),
.Y(n_7117)
);

AOI21xp5_ASAP7_75t_L g7118 ( 
.A1(n_6167),
.A2(n_5437),
.B(n_5434),
.Y(n_7118)
);

NAND2xp5_ASAP7_75t_L g7119 ( 
.A(n_5545),
.B(n_5556),
.Y(n_7119)
);

AOI21xp5_ASAP7_75t_L g7120 ( 
.A1(n_5434),
.A2(n_5442),
.B(n_5437),
.Y(n_7120)
);

INVxp67_ASAP7_75t_L g7121 ( 
.A(n_5151),
.Y(n_7121)
);

AOI21xp5_ASAP7_75t_L g7122 ( 
.A1(n_5442),
.A2(n_5536),
.B(n_5208),
.Y(n_7122)
);

AOI21xp5_ASAP7_75t_L g7123 ( 
.A1(n_5930),
.A2(n_5957),
.B(n_5300),
.Y(n_7123)
);

BUFx2_ASAP7_75t_L g7124 ( 
.A(n_5879),
.Y(n_7124)
);

CKINVDCx16_ASAP7_75t_R g7125 ( 
.A(n_5722),
.Y(n_7125)
);

OAI21x1_ASAP7_75t_L g7126 ( 
.A1(n_5880),
.A2(n_6064),
.B(n_4808),
.Y(n_7126)
);

OR2x2_ASAP7_75t_L g7127 ( 
.A(n_5634),
.B(n_5679),
.Y(n_7127)
);

CKINVDCx20_ASAP7_75t_R g7128 ( 
.A(n_5514),
.Y(n_7128)
);

OAI21x1_ASAP7_75t_L g7129 ( 
.A1(n_5880),
.A2(n_6064),
.B(n_4808),
.Y(n_7129)
);

AOI21xp5_ASAP7_75t_L g7130 ( 
.A1(n_5982),
.A2(n_5340),
.B(n_5335),
.Y(n_7130)
);

AOI21xp5_ASAP7_75t_L g7131 ( 
.A1(n_5335),
.A2(n_5352),
.B(n_5340),
.Y(n_7131)
);

BUFx8_ASAP7_75t_SL g7132 ( 
.A(n_5865),
.Y(n_7132)
);

O2A1O1Ixp5_ASAP7_75t_L g7133 ( 
.A1(n_5527),
.A2(n_5571),
.B(n_5546),
.C(n_5761),
.Y(n_7133)
);

AO21x1_ASAP7_75t_L g7134 ( 
.A1(n_6230),
.A2(n_6249),
.B(n_6044),
.Y(n_7134)
);

OAI22xp5_ASAP7_75t_L g7135 ( 
.A1(n_5134),
.A2(n_5145),
.B1(n_5172),
.B2(n_5154),
.Y(n_7135)
);

CKINVDCx5p33_ASAP7_75t_R g7136 ( 
.A(n_5082),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_5358),
.Y(n_7137)
);

AOI21xp5_ASAP7_75t_L g7138 ( 
.A1(n_5352),
.A2(n_5371),
.B(n_5357),
.Y(n_7138)
);

NAND2xp5_ASAP7_75t_L g7139 ( 
.A(n_5578),
.B(n_5601),
.Y(n_7139)
);

NAND2xp5_ASAP7_75t_SL g7140 ( 
.A(n_5357),
.B(n_5371),
.Y(n_7140)
);

OAI21xp5_ASAP7_75t_L g7141 ( 
.A1(n_5475),
.A2(n_5591),
.B(n_5587),
.Y(n_7141)
);

AOI21x1_ASAP7_75t_L g7142 ( 
.A1(n_5551),
.A2(n_5363),
.B(n_5361),
.Y(n_7142)
);

AOI21xp5_ASAP7_75t_L g7143 ( 
.A1(n_5375),
.A2(n_5381),
.B(n_5376),
.Y(n_7143)
);

OAI21xp5_ASAP7_75t_L g7144 ( 
.A1(n_5587),
.A2(n_5591),
.B(n_5601),
.Y(n_7144)
);

OAI21x1_ASAP7_75t_L g7145 ( 
.A1(n_6064),
.A2(n_4808),
.B(n_4734),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_5361),
.Y(n_7146)
);

OAI21x1_ASAP7_75t_L g7147 ( 
.A1(n_6064),
.A2(n_4808),
.B(n_4734),
.Y(n_7147)
);

INVxp67_ASAP7_75t_L g7148 ( 
.A(n_5182),
.Y(n_7148)
);

NAND2xp5_ASAP7_75t_L g7149 ( 
.A(n_5331),
.B(n_5248),
.Y(n_7149)
);

BUFx2_ASAP7_75t_L g7150 ( 
.A(n_5879),
.Y(n_7150)
);

OAI21xp5_ASAP7_75t_L g7151 ( 
.A1(n_5557),
.A2(n_5518),
.B(n_5855),
.Y(n_7151)
);

CKINVDCx5p33_ASAP7_75t_R g7152 ( 
.A(n_5360),
.Y(n_7152)
);

BUFx3_ASAP7_75t_L g7153 ( 
.A(n_5722),
.Y(n_7153)
);

AOI22xp33_ASAP7_75t_L g7154 ( 
.A1(n_5090),
.A2(n_5094),
.B1(n_5226),
.B2(n_5517),
.Y(n_7154)
);

OAI21x1_ASAP7_75t_L g7155 ( 
.A1(n_4734),
.A2(n_4974),
.B(n_4939),
.Y(n_7155)
);

AOI21x1_ASAP7_75t_L g7156 ( 
.A1(n_5370),
.A2(n_5455),
.B(n_5435),
.Y(n_7156)
);

NAND2xp5_ASAP7_75t_L g7157 ( 
.A(n_5331),
.B(n_5248),
.Y(n_7157)
);

OAI21x1_ASAP7_75t_L g7158 ( 
.A1(n_4734),
.A2(n_4974),
.B(n_4939),
.Y(n_7158)
);

INVxp67_ASAP7_75t_SL g7159 ( 
.A(n_5435),
.Y(n_7159)
);

INVx1_ASAP7_75t_L g7160 ( 
.A(n_5455),
.Y(n_7160)
);

NAND2xp5_ASAP7_75t_L g7161 ( 
.A(n_5089),
.B(n_5103),
.Y(n_7161)
);

BUFx2_ASAP7_75t_L g7162 ( 
.A(n_5879),
.Y(n_7162)
);

AOI21xp5_ASAP7_75t_L g7163 ( 
.A1(n_5375),
.A2(n_5381),
.B(n_5376),
.Y(n_7163)
);

AOI21xp5_ASAP7_75t_L g7164 ( 
.A1(n_5385),
.A2(n_5395),
.B(n_5394),
.Y(n_7164)
);

NAND2xp5_ASAP7_75t_L g7165 ( 
.A(n_5089),
.B(n_5103),
.Y(n_7165)
);

AOI21xp5_ASAP7_75t_L g7166 ( 
.A1(n_5385),
.A2(n_5395),
.B(n_5394),
.Y(n_7166)
);

O2A1O1Ixp5_ASAP7_75t_L g7167 ( 
.A1(n_5761),
.A2(n_6184),
.B(n_6081),
.C(n_6090),
.Y(n_7167)
);

AO21x1_ASAP7_75t_L g7168 ( 
.A1(n_6249),
.A2(n_5720),
.B(n_5694),
.Y(n_7168)
);

AOI21xp5_ASAP7_75t_L g7169 ( 
.A1(n_5408),
.A2(n_5413),
.B(n_6048),
.Y(n_7169)
);

OAI21x1_ASAP7_75t_L g7170 ( 
.A1(n_4939),
.A2(n_4996),
.B(n_4974),
.Y(n_7170)
);

NOR2x1_ASAP7_75t_L g7171 ( 
.A(n_5958),
.B(n_5882),
.Y(n_7171)
);

OAI21x1_ASAP7_75t_L g7172 ( 
.A1(n_4939),
.A2(n_4996),
.B(n_4974),
.Y(n_7172)
);

OAI21x1_ASAP7_75t_L g7173 ( 
.A1(n_4996),
.A2(n_5060),
.B(n_5047),
.Y(n_7173)
);

NAND2xp5_ASAP7_75t_SL g7174 ( 
.A(n_5408),
.B(n_5413),
.Y(n_7174)
);

NAND2xp5_ASAP7_75t_L g7175 ( 
.A(n_5144),
.B(n_5170),
.Y(n_7175)
);

OAI21x1_ASAP7_75t_L g7176 ( 
.A1(n_4996),
.A2(n_5060),
.B(n_5047),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_5471),
.Y(n_7177)
);

AOI21xp33_ASAP7_75t_L g7178 ( 
.A1(n_5498),
.A2(n_5616),
.B(n_5557),
.Y(n_7178)
);

OAI21xp5_ASAP7_75t_L g7179 ( 
.A1(n_5855),
.A2(n_5616),
.B(n_5830),
.Y(n_7179)
);

OAI22xp5_ASAP7_75t_L g7180 ( 
.A1(n_5135),
.A2(n_6214),
.B1(n_5321),
.B2(n_5170),
.Y(n_7180)
);

AO21x1_ASAP7_75t_L g7181 ( 
.A1(n_5694),
.A2(n_5720),
.B(n_6162),
.Y(n_7181)
);

OAI21x1_ASAP7_75t_L g7182 ( 
.A1(n_5047),
.A2(n_5068),
.B(n_5060),
.Y(n_7182)
);

OR2x6_ASAP7_75t_L g7183 ( 
.A(n_5251),
.B(n_4733),
.Y(n_7183)
);

INVx1_ASAP7_75t_SL g7184 ( 
.A(n_5757),
.Y(n_7184)
);

OAI21x1_ASAP7_75t_SL g7185 ( 
.A1(n_6209),
.A2(n_6243),
.B(n_5889),
.Y(n_7185)
);

INVx1_ASAP7_75t_L g7186 ( 
.A(n_5471),
.Y(n_7186)
);

AOI21xp5_ASAP7_75t_L g7187 ( 
.A1(n_6048),
.A2(n_6037),
.B(n_4938),
.Y(n_7187)
);

NAND2xp5_ASAP7_75t_L g7188 ( 
.A(n_5144),
.B(n_5565),
.Y(n_7188)
);

NAND2xp5_ASAP7_75t_SL g7189 ( 
.A(n_5830),
.B(n_5550),
.Y(n_7189)
);

NOR2xp67_ASAP7_75t_SL g7190 ( 
.A(n_4761),
.B(n_5360),
.Y(n_7190)
);

NAND2xp5_ASAP7_75t_SL g7191 ( 
.A(n_5550),
.B(n_6229),
.Y(n_7191)
);

NAND2xp5_ASAP7_75t_SL g7192 ( 
.A(n_6180),
.B(n_6037),
.Y(n_7192)
);

AO21x1_ASAP7_75t_L g7193 ( 
.A1(n_5480),
.A2(n_5529),
.B(n_5501),
.Y(n_7193)
);

AND2x4_ASAP7_75t_L g7194 ( 
.A(n_4783),
.B(n_4792),
.Y(n_7194)
);

NAND2xp5_ASAP7_75t_L g7195 ( 
.A(n_5565),
.B(n_5328),
.Y(n_7195)
);

HB1xp67_ASAP7_75t_L g7196 ( 
.A(n_6026),
.Y(n_7196)
);

AOI21xp33_ASAP7_75t_L g7197 ( 
.A1(n_5498),
.A2(n_5537),
.B(n_5502),
.Y(n_7197)
);

INVx1_ASAP7_75t_SL g7198 ( 
.A(n_5182),
.Y(n_7198)
);

NAND2xp5_ASAP7_75t_L g7199 ( 
.A(n_5328),
.B(n_5330),
.Y(n_7199)
);

OAI22xp5_ASAP7_75t_L g7200 ( 
.A1(n_5321),
.A2(n_6214),
.B1(n_5549),
.B2(n_5541),
.Y(n_7200)
);

NAND2x1p5_ASAP7_75t_L g7201 ( 
.A(n_4907),
.B(n_5017),
.Y(n_7201)
);

AOI21x1_ASAP7_75t_L g7202 ( 
.A1(n_5501),
.A2(n_5539),
.B(n_5529),
.Y(n_7202)
);

AOI21xp5_ASAP7_75t_L g7203 ( 
.A1(n_6048),
.A2(n_4938),
.B(n_4889),
.Y(n_7203)
);

AO31x2_ASAP7_75t_L g7204 ( 
.A1(n_5539),
.A2(n_5563),
.A3(n_5580),
.B(n_5552),
.Y(n_7204)
);

OAI21x1_ASAP7_75t_L g7205 ( 
.A1(n_5047),
.A2(n_5068),
.B(n_5060),
.Y(n_7205)
);

NAND3xp33_ASAP7_75t_L g7206 ( 
.A(n_5918),
.B(n_5864),
.C(n_5537),
.Y(n_7206)
);

AOI22xp5_ASAP7_75t_L g7207 ( 
.A1(n_5502),
.A2(n_5498),
.B1(n_6180),
.B2(n_5643),
.Y(n_7207)
);

AND2x4_ASAP7_75t_L g7208 ( 
.A(n_4792),
.B(n_4800),
.Y(n_7208)
);

BUFx12f_ASAP7_75t_L g7209 ( 
.A(n_5360),
.Y(n_7209)
);

NAND2xp5_ASAP7_75t_L g7210 ( 
.A(n_5330),
.B(n_5253),
.Y(n_7210)
);

AND2x2_ASAP7_75t_L g7211 ( 
.A(n_4800),
.B(n_4862),
.Y(n_7211)
);

OAI21x1_ASAP7_75t_L g7212 ( 
.A1(n_5068),
.A2(n_5382),
.B(n_5222),
.Y(n_7212)
);

AOI21xp5_ASAP7_75t_L g7213 ( 
.A1(n_6048),
.A2(n_4938),
.B(n_4889),
.Y(n_7213)
);

NAND2xp5_ASAP7_75t_L g7214 ( 
.A(n_5253),
.B(n_5899),
.Y(n_7214)
);

AND2x2_ASAP7_75t_L g7215 ( 
.A(n_4862),
.B(n_4881),
.Y(n_7215)
);

OAI21xp5_ASAP7_75t_L g7216 ( 
.A1(n_5958),
.A2(n_5798),
.B(n_5795),
.Y(n_7216)
);

OAI21xp5_ASAP7_75t_L g7217 ( 
.A1(n_5995),
.A2(n_6083),
.B(n_6068),
.Y(n_7217)
);

NAND2xp5_ASAP7_75t_L g7218 ( 
.A(n_5899),
.B(n_5903),
.Y(n_7218)
);

OAI21x1_ASAP7_75t_L g7219 ( 
.A1(n_5068),
.A2(n_5382),
.B(n_5222),
.Y(n_7219)
);

AOI21x1_ASAP7_75t_L g7220 ( 
.A1(n_5563),
.A2(n_5586),
.B(n_5580),
.Y(n_7220)
);

INVx1_ASAP7_75t_SL g7221 ( 
.A(n_5219),
.Y(n_7221)
);

AO31x2_ASAP7_75t_L g7222 ( 
.A1(n_5594),
.A2(n_5598),
.A3(n_5608),
.B(n_5596),
.Y(n_7222)
);

OAI21x1_ASAP7_75t_L g7223 ( 
.A1(n_5222),
.A2(n_5432),
.B(n_5382),
.Y(n_7223)
);

NAND2xp5_ASAP7_75t_SL g7224 ( 
.A(n_5731),
.B(n_5498),
.Y(n_7224)
);

AOI21xp5_ASAP7_75t_L g7225 ( 
.A1(n_4938),
.A2(n_5191),
.B(n_5138),
.Y(n_7225)
);

AND2x4_ASAP7_75t_L g7226 ( 
.A(n_4962),
.B(n_4968),
.Y(n_7226)
);

INVx1_ASAP7_75t_L g7227 ( 
.A(n_5598),
.Y(n_7227)
);

NAND2xp5_ASAP7_75t_L g7228 ( 
.A(n_5423),
.B(n_5428),
.Y(n_7228)
);

BUFx3_ASAP7_75t_L g7229 ( 
.A(n_5876),
.Y(n_7229)
);

NAND2x1p5_ASAP7_75t_L g7230 ( 
.A(n_4907),
.B(n_5017),
.Y(n_7230)
);

AND2x4_ASAP7_75t_L g7231 ( 
.A(n_4962),
.B(n_4968),
.Y(n_7231)
);

INVx4_ASAP7_75t_L g7232 ( 
.A(n_5251),
.Y(n_7232)
);

BUFx6f_ASAP7_75t_L g7233 ( 
.A(n_4907),
.Y(n_7233)
);

AND2x4_ASAP7_75t_L g7234 ( 
.A(n_4968),
.B(n_5001),
.Y(n_7234)
);

OAI21xp5_ASAP7_75t_L g7235 ( 
.A1(n_5995),
.A2(n_6083),
.B(n_6068),
.Y(n_7235)
);

OAI22xp5_ASAP7_75t_L g7236 ( 
.A1(n_5541),
.A2(n_5549),
.B1(n_5486),
.B2(n_5485),
.Y(n_7236)
);

OAI21xp5_ASAP7_75t_L g7237 ( 
.A1(n_5633),
.A2(n_6042),
.B(n_5864),
.Y(n_7237)
);

OAI21x1_ASAP7_75t_L g7238 ( 
.A1(n_5613),
.A2(n_6169),
.B(n_5615),
.Y(n_7238)
);

INVx2_ASAP7_75t_L g7239 ( 
.A(n_5612),
.Y(n_7239)
);

OAI21x1_ASAP7_75t_L g7240 ( 
.A1(n_5613),
.A2(n_6169),
.B(n_5615),
.Y(n_7240)
);

AOI21xp5_ASAP7_75t_L g7241 ( 
.A1(n_5138),
.A2(n_5191),
.B(n_4889),
.Y(n_7241)
);

NOR2xp33_ASAP7_75t_SL g7242 ( 
.A(n_5756),
.B(n_4889),
.Y(n_7242)
);

NAND2xp5_ASAP7_75t_SL g7243 ( 
.A(n_5731),
.B(n_6128),
.Y(n_7243)
);

OAI21xp5_ASAP7_75t_L g7244 ( 
.A1(n_6042),
.A2(n_6187),
.B(n_5889),
.Y(n_7244)
);

AOI21xp5_ASAP7_75t_L g7245 ( 
.A1(n_5138),
.A2(n_5191),
.B(n_5668),
.Y(n_7245)
);

OR2x6_ASAP7_75t_L g7246 ( 
.A(n_4733),
.B(n_4763),
.Y(n_7246)
);

OAI21x1_ASAP7_75t_L g7247 ( 
.A1(n_5612),
.A2(n_5619),
.B(n_5617),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_SL g7248 ( 
.A(n_6128),
.B(n_6210),
.Y(n_7248)
);

A2O1A1Ixp33_ASAP7_75t_L g7249 ( 
.A1(n_5647),
.A2(n_5040),
.B(n_4899),
.C(n_6210),
.Y(n_7249)
);

AO21x1_ASAP7_75t_L g7250 ( 
.A1(n_5617),
.A2(n_5631),
.B(n_5619),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_5631),
.Y(n_7251)
);

OAI21x1_ASAP7_75t_L g7252 ( 
.A1(n_5659),
.A2(n_5674),
.B(n_5667),
.Y(n_7252)
);

INVx2_ASAP7_75t_SL g7253 ( 
.A(n_6056),
.Y(n_7253)
);

AOI21xp5_ASAP7_75t_L g7254 ( 
.A1(n_5191),
.A2(n_5138),
.B(n_5668),
.Y(n_7254)
);

INVx1_ASAP7_75t_L g7255 ( 
.A(n_5659),
.Y(n_7255)
);

OAI21xp5_ASAP7_75t_L g7256 ( 
.A1(n_6187),
.A2(n_5887),
.B(n_6161),
.Y(n_7256)
);

INVx1_ASAP7_75t_L g7257 ( 
.A(n_5667),
.Y(n_7257)
);

NAND2xp5_ASAP7_75t_L g7258 ( 
.A(n_5428),
.B(n_5150),
.Y(n_7258)
);

OAI21x1_ASAP7_75t_L g7259 ( 
.A1(n_5674),
.A2(n_5699),
.B(n_5688),
.Y(n_7259)
);

NAND2xp5_ASAP7_75t_SL g7260 ( 
.A(n_6134),
.B(n_5762),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_5699),
.Y(n_7261)
);

INVxp67_ASAP7_75t_L g7262 ( 
.A(n_5219),
.Y(n_7262)
);

CKINVDCx11_ASAP7_75t_R g7263 ( 
.A(n_6196),
.Y(n_7263)
);

OAI21x1_ASAP7_75t_L g7264 ( 
.A1(n_5701),
.A2(n_5726),
.B(n_5725),
.Y(n_7264)
);

AOI21xp5_ASAP7_75t_L g7265 ( 
.A1(n_6107),
.A2(n_6207),
.B(n_5261),
.Y(n_7265)
);

INVxp67_ASAP7_75t_SL g7266 ( 
.A(n_5701),
.Y(n_7266)
);

OAI21xp5_ASAP7_75t_L g7267 ( 
.A1(n_5887),
.A2(n_6177),
.B(n_5762),
.Y(n_7267)
);

NAND2xp5_ASAP7_75t_L g7268 ( 
.A(n_5157),
.B(n_5163),
.Y(n_7268)
);

O2A1O1Ixp33_ASAP7_75t_L g7269 ( 
.A1(n_4880),
.A2(n_4949),
.B(n_5010),
.C(n_4943),
.Y(n_7269)
);

INVx3_ASAP7_75t_L g7270 ( 
.A(n_6056),
.Y(n_7270)
);

NAND2x1p5_ASAP7_75t_L g7271 ( 
.A(n_4907),
.B(n_5017),
.Y(n_7271)
);

AOI21xp5_ASAP7_75t_L g7272 ( 
.A1(n_6107),
.A2(n_5261),
.B(n_5122),
.Y(n_7272)
);

AOI21xp5_ASAP7_75t_L g7273 ( 
.A1(n_6107),
.A2(n_5261),
.B(n_5122),
.Y(n_7273)
);

AOI21xp5_ASAP7_75t_L g7274 ( 
.A1(n_5122),
.A2(n_5453),
.B(n_5329),
.Y(n_7274)
);

NAND2xp5_ASAP7_75t_L g7275 ( 
.A(n_5164),
.B(n_5168),
.Y(n_7275)
);

AOI22xp5_ASAP7_75t_L g7276 ( 
.A1(n_5638),
.A2(n_6111),
.B1(n_5742),
.B2(n_6236),
.Y(n_7276)
);

OAI21x1_ASAP7_75t_L g7277 ( 
.A1(n_5725),
.A2(n_5729),
.B(n_5726),
.Y(n_7277)
);

NAND2xp5_ASAP7_75t_L g7278 ( 
.A(n_5189),
.B(n_5062),
.Y(n_7278)
);

AOI21xp5_ASAP7_75t_L g7279 ( 
.A1(n_5329),
.A2(n_5453),
.B(n_5676),
.Y(n_7279)
);

NOR2xp33_ASAP7_75t_L g7280 ( 
.A(n_5189),
.B(n_6134),
.Y(n_7280)
);

INVx1_ASAP7_75t_L g7281 ( 
.A(n_5729),
.Y(n_7281)
);

AOI21x1_ASAP7_75t_L g7282 ( 
.A1(n_5748),
.A2(n_5765),
.B(n_5749),
.Y(n_7282)
);

AOI221xp5_ASAP7_75t_SL g7283 ( 
.A1(n_5743),
.A2(n_5755),
.B1(n_5721),
.B2(n_5278),
.C(n_5589),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_5748),
.Y(n_7284)
);

NAND2x1p5_ASAP7_75t_L g7285 ( 
.A(n_5017),
.B(n_5049),
.Y(n_7285)
);

OAI21xp5_ASAP7_75t_L g7286 ( 
.A1(n_5562),
.A2(n_5610),
.B(n_5882),
.Y(n_7286)
);

OAI21x1_ASAP7_75t_L g7287 ( 
.A1(n_5749),
.A2(n_5803),
.B(n_5765),
.Y(n_7287)
);

NOR2xp33_ASAP7_75t_L g7288 ( 
.A(n_5758),
.B(n_5776),
.Y(n_7288)
);

NAND2xp5_ASAP7_75t_L g7289 ( 
.A(n_5062),
.B(n_5063),
.Y(n_7289)
);

INVx1_ASAP7_75t_L g7290 ( 
.A(n_5803),
.Y(n_7290)
);

AOI21x1_ASAP7_75t_L g7291 ( 
.A1(n_5835),
.A2(n_5847),
.B(n_5836),
.Y(n_7291)
);

OAI21x1_ASAP7_75t_L g7292 ( 
.A1(n_5835),
.A2(n_5847),
.B(n_5836),
.Y(n_7292)
);

OAI21x1_ASAP7_75t_L g7293 ( 
.A1(n_5859),
.A2(n_5907),
.B(n_5873),
.Y(n_7293)
);

INVx1_ASAP7_75t_L g7294 ( 
.A(n_5859),
.Y(n_7294)
);

NAND2xp5_ASAP7_75t_L g7295 ( 
.A(n_5062),
.B(n_5063),
.Y(n_7295)
);

NAND2xp5_ASAP7_75t_L g7296 ( 
.A(n_5063),
.B(n_5080),
.Y(n_7296)
);

AOI21xp5_ASAP7_75t_L g7297 ( 
.A1(n_5329),
.A2(n_5453),
.B(n_5901),
.Y(n_7297)
);

A2O1A1Ixp33_ASAP7_75t_L g7298 ( 
.A1(n_4762),
.A2(n_4804),
.B(n_4818),
.C(n_4767),
.Y(n_7298)
);

AOI21x1_ASAP7_75t_L g7299 ( 
.A1(n_5873),
.A2(n_5919),
.B(n_5907),
.Y(n_7299)
);

AO31x2_ASAP7_75t_L g7300 ( 
.A1(n_5919),
.A2(n_4767),
.A3(n_4818),
.B(n_4804),
.Y(n_7300)
);

AOI21xp5_ASAP7_75t_L g7301 ( 
.A1(n_6056),
.A2(n_6135),
.B(n_6112),
.Y(n_7301)
);

INVx2_ASAP7_75t_SL g7302 ( 
.A(n_6056),
.Y(n_7302)
);

OAI21xp5_ASAP7_75t_L g7303 ( 
.A1(n_5931),
.A2(n_6140),
.B(n_6114),
.Y(n_7303)
);

NOR2xp33_ASAP7_75t_L g7304 ( 
.A(n_5842),
.B(n_5897),
.Y(n_7304)
);

AOI21xp5_ASAP7_75t_L g7305 ( 
.A1(n_6112),
.A2(n_6135),
.B(n_5751),
.Y(n_7305)
);

A2O1A1Ixp33_ASAP7_75t_L g7306 ( 
.A1(n_4834),
.A2(n_5058),
.B(n_5041),
.C(n_6006),
.Y(n_7306)
);

OAI21xp5_ASAP7_75t_L g7307 ( 
.A1(n_5931),
.A2(n_6140),
.B(n_6114),
.Y(n_7307)
);

INVx5_ASAP7_75t_L g7308 ( 
.A(n_5017),
.Y(n_7308)
);

NOR2x1_ASAP7_75t_L g7309 ( 
.A(n_5973),
.B(n_5840),
.Y(n_7309)
);

NAND2xp5_ASAP7_75t_L g7310 ( 
.A(n_4791),
.B(n_4811),
.Y(n_7310)
);

BUFx2_ASAP7_75t_L g7311 ( 
.A(n_5558),
.Y(n_7311)
);

AOI21xp5_ASAP7_75t_L g7312 ( 
.A1(n_6112),
.A2(n_6135),
.B(n_5766),
.Y(n_7312)
);

AO31x2_ASAP7_75t_L g7313 ( 
.A1(n_4834),
.A2(n_5058),
.A3(n_5041),
.B(n_6122),
.Y(n_7313)
);

AOI21xp5_ASAP7_75t_L g7314 ( 
.A1(n_6112),
.A2(n_6135),
.B(n_5780),
.Y(n_7314)
);

AND2x4_ASAP7_75t_L g7315 ( 
.A(n_5006),
.B(n_5026),
.Y(n_7315)
);

OAI21x1_ASAP7_75t_L g7316 ( 
.A1(n_5649),
.A2(n_5777),
.B(n_5715),
.Y(n_7316)
);

AOI21xp5_ASAP7_75t_L g7317 ( 
.A1(n_6112),
.A2(n_6135),
.B(n_5713),
.Y(n_7317)
);

CKINVDCx6p67_ASAP7_75t_R g7318 ( 
.A(n_4832),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_6116),
.Y(n_7319)
);

OAI21xp33_ASAP7_75t_L g7320 ( 
.A1(n_5567),
.A2(n_6181),
.B(n_5533),
.Y(n_7320)
);

BUFx6f_ASAP7_75t_L g7321 ( 
.A(n_5017),
.Y(n_7321)
);

NAND2xp5_ASAP7_75t_L g7322 ( 
.A(n_4791),
.B(n_4811),
.Y(n_7322)
);

NAND2xp5_ASAP7_75t_SL g7323 ( 
.A(n_6171),
.B(n_6251),
.Y(n_7323)
);

BUFx6f_ASAP7_75t_L g7324 ( 
.A(n_5017),
.Y(n_7324)
);

OAI21x1_ASAP7_75t_L g7325 ( 
.A1(n_5649),
.A2(n_5777),
.B(n_5715),
.Y(n_7325)
);

NAND2xp5_ASAP7_75t_L g7326 ( 
.A(n_4815),
.B(n_4835),
.Y(n_7326)
);

AOI21x1_ASAP7_75t_L g7327 ( 
.A1(n_5831),
.A2(n_6123),
.B(n_5973),
.Y(n_7327)
);

A2O1A1Ixp33_ASAP7_75t_L g7328 ( 
.A1(n_6171),
.A2(n_6251),
.B(n_5817),
.C(n_5304),
.Y(n_7328)
);

AOI22xp5_ASAP7_75t_L g7329 ( 
.A1(n_5710),
.A2(n_5927),
.B1(n_5932),
.B2(n_6088),
.Y(n_7329)
);

OAI21xp5_ASAP7_75t_L g7330 ( 
.A1(n_6101),
.A2(n_5817),
.B(n_5936),
.Y(n_7330)
);

OAI21xp33_ASAP7_75t_L g7331 ( 
.A1(n_6181),
.A2(n_5468),
.B(n_5794),
.Y(n_7331)
);

CKINVDCx5p33_ASAP7_75t_R g7332 ( 
.A(n_5692),
.Y(n_7332)
);

OR2x2_ASAP7_75t_L g7333 ( 
.A(n_5634),
.B(n_5679),
.Y(n_7333)
);

A2O1A1Ixp33_ASAP7_75t_L g7334 ( 
.A1(n_5706),
.A2(n_5636),
.B(n_5648),
.C(n_5721),
.Y(n_7334)
);

OAI21x1_ASAP7_75t_L g7335 ( 
.A1(n_5848),
.A2(n_5894),
.B(n_5863),
.Y(n_7335)
);

OAI21xp5_ASAP7_75t_L g7336 ( 
.A1(n_6101),
.A2(n_5980),
.B(n_5936),
.Y(n_7336)
);

AOI21xp5_ASAP7_75t_L g7337 ( 
.A1(n_6112),
.A2(n_6135),
.B(n_5055),
.Y(n_7337)
);

INVx4_ASAP7_75t_L g7338 ( 
.A(n_5049),
.Y(n_7338)
);

INVx3_ASAP7_75t_L g7339 ( 
.A(n_6112),
.Y(n_7339)
);

HB1xp67_ASAP7_75t_L g7340 ( 
.A(n_6026),
.Y(n_7340)
);

OAI21xp5_ASAP7_75t_L g7341 ( 
.A1(n_5980),
.A2(n_5997),
.B(n_5033),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_4815),
.B(n_4835),
.Y(n_7342)
);

O2A1O1Ixp5_ASAP7_75t_L g7343 ( 
.A1(n_6052),
.A2(n_6121),
.B(n_6133),
.C(n_6110),
.Y(n_7343)
);

NAND2xp5_ASAP7_75t_SL g7344 ( 
.A(n_5997),
.B(n_6145),
.Y(n_7344)
);

NAND2xp5_ASAP7_75t_L g7345 ( 
.A(n_4845),
.B(n_5327),
.Y(n_7345)
);

INVx3_ASAP7_75t_L g7346 ( 
.A(n_6135),
.Y(n_7346)
);

INVx4_ASAP7_75t_L g7347 ( 
.A(n_5049),
.Y(n_7347)
);

INVx5_ASAP7_75t_L g7348 ( 
.A(n_5049),
.Y(n_7348)
);

OAI21xp33_ASAP7_75t_L g7349 ( 
.A1(n_5184),
.A2(n_5302),
.B(n_5244),
.Y(n_7349)
);

AND2x4_ASAP7_75t_L g7350 ( 
.A(n_5036),
.B(n_5044),
.Y(n_7350)
);

OR2x6_ASAP7_75t_L g7351 ( 
.A(n_4733),
.B(n_4763),
.Y(n_7351)
);

AND2x2_ASAP7_75t_L g7352 ( 
.A(n_5036),
.B(n_5044),
.Y(n_7352)
);

A2O1A1Ixp33_ASAP7_75t_L g7353 ( 
.A1(n_5743),
.A2(n_5755),
.B(n_5738),
.C(n_6145),
.Y(n_7353)
);

AOI21xp5_ASAP7_75t_L g7354 ( 
.A1(n_5049),
.A2(n_5088),
.B(n_5055),
.Y(n_7354)
);

AOI21xp5_ASAP7_75t_L g7355 ( 
.A1(n_5049),
.A2(n_5088),
.B(n_5055),
.Y(n_7355)
);

NAND2xp5_ASAP7_75t_SL g7356 ( 
.A(n_5998),
.B(n_6070),
.Y(n_7356)
);

NAND2xp5_ASAP7_75t_L g7357 ( 
.A(n_4845),
.B(n_5327),
.Y(n_7357)
);

OAI21x1_ASAP7_75t_L g7358 ( 
.A1(n_5848),
.A2(n_5894),
.B(n_5863),
.Y(n_7358)
);

BUFx6f_ASAP7_75t_L g7359 ( 
.A(n_5049),
.Y(n_7359)
);

INVx5_ASAP7_75t_L g7360 ( 
.A(n_5055),
.Y(n_7360)
);

OAI21xp5_ASAP7_75t_L g7361 ( 
.A1(n_4764),
.A2(n_5048),
.B(n_5033),
.Y(n_7361)
);

NAND2xp5_ASAP7_75t_L g7362 ( 
.A(n_5372),
.B(n_5384),
.Y(n_7362)
);

OAI21x1_ASAP7_75t_L g7363 ( 
.A1(n_5911),
.A2(n_5558),
.B(n_6122),
.Y(n_7363)
);

BUFx3_ASAP7_75t_L g7364 ( 
.A(n_5558),
.Y(n_7364)
);

OAI21x1_ASAP7_75t_L g7365 ( 
.A1(n_5911),
.A2(n_5558),
.B(n_6122),
.Y(n_7365)
);

NAND2xp5_ASAP7_75t_L g7366 ( 
.A(n_5372),
.B(n_5384),
.Y(n_7366)
);

OAI21x1_ASAP7_75t_L g7367 ( 
.A1(n_5911),
.A2(n_6157),
.B(n_6131),
.Y(n_7367)
);

OAI22xp33_ASAP7_75t_L g7368 ( 
.A1(n_5077),
.A2(n_5932),
.B1(n_5927),
.B2(n_6196),
.Y(n_7368)
);

INVx2_ASAP7_75t_SL g7369 ( 
.A(n_5752),
.Y(n_7369)
);

CKINVDCx5p33_ASAP7_75t_R g7370 ( 
.A(n_5719),
.Y(n_7370)
);

OAI21x1_ASAP7_75t_SL g7371 ( 
.A1(n_6049),
.A2(n_6055),
.B(n_6051),
.Y(n_7371)
);

AOI21xp5_ASAP7_75t_L g7372 ( 
.A1(n_5055),
.A2(n_5114),
.B(n_5088),
.Y(n_7372)
);

AOI21xp33_ASAP7_75t_L g7373 ( 
.A1(n_5928),
.A2(n_5913),
.B(n_5926),
.Y(n_7373)
);

OAI21x1_ASAP7_75t_L g7374 ( 
.A1(n_5911),
.A2(n_6157),
.B(n_6131),
.Y(n_7374)
);

AOI21xp5_ASAP7_75t_L g7375 ( 
.A1(n_5055),
.A2(n_5114),
.B(n_5088),
.Y(n_7375)
);

AOI21xp5_ASAP7_75t_L g7376 ( 
.A1(n_5088),
.A2(n_5123),
.B(n_5114),
.Y(n_7376)
);

AOI21x1_ASAP7_75t_L g7377 ( 
.A1(n_5831),
.A2(n_6123),
.B(n_5654),
.Y(n_7377)
);

AOI21xp5_ASAP7_75t_L g7378 ( 
.A1(n_5088),
.A2(n_5123),
.B(n_5114),
.Y(n_7378)
);

NAND2xp5_ASAP7_75t_L g7379 ( 
.A(n_5274),
.B(n_5289),
.Y(n_7379)
);

INVx3_ASAP7_75t_L g7380 ( 
.A(n_4771),
.Y(n_7380)
);

OAI21x1_ASAP7_75t_L g7381 ( 
.A1(n_6131),
.A2(n_6165),
.B(n_6157),
.Y(n_7381)
);

AOI21xp5_ASAP7_75t_L g7382 ( 
.A1(n_5114),
.A2(n_5124),
.B(n_5123),
.Y(n_7382)
);

BUFx12f_ASAP7_75t_L g7383 ( 
.A(n_5514),
.Y(n_7383)
);

NOR2xp67_ASAP7_75t_L g7384 ( 
.A(n_5044),
.B(n_5067),
.Y(n_7384)
);

NAND2xp5_ASAP7_75t_L g7385 ( 
.A(n_5289),
.B(n_5297),
.Y(n_7385)
);

NAND2xp5_ASAP7_75t_SL g7386 ( 
.A(n_5998),
.B(n_6070),
.Y(n_7386)
);

OAI21xp5_ASAP7_75t_L g7387 ( 
.A1(n_4764),
.A2(n_5076),
.B(n_5048),
.Y(n_7387)
);

A2O1A1Ixp33_ASAP7_75t_L g7388 ( 
.A1(n_6218),
.A2(n_6232),
.B(n_6231),
.C(n_6241),
.Y(n_7388)
);

NAND2xp5_ASAP7_75t_L g7389 ( 
.A(n_5297),
.B(n_5299),
.Y(n_7389)
);

NAND2xp5_ASAP7_75t_L g7390 ( 
.A(n_5299),
.B(n_5303),
.Y(n_7390)
);

OAI21xp5_ASAP7_75t_L g7391 ( 
.A1(n_5076),
.A2(n_6125),
.B(n_6124),
.Y(n_7391)
);

AND2x2_ASAP7_75t_L g7392 ( 
.A(n_5067),
.B(n_5100),
.Y(n_7392)
);

AOI21xp5_ASAP7_75t_L g7393 ( 
.A1(n_5114),
.A2(n_5124),
.B(n_5123),
.Y(n_7393)
);

OAI21xp5_ASAP7_75t_L g7394 ( 
.A1(n_6124),
.A2(n_6206),
.B(n_6125),
.Y(n_7394)
);

OAI21x1_ASAP7_75t_L g7395 ( 
.A1(n_6185),
.A2(n_6186),
.B(n_6143),
.Y(n_7395)
);

OAI21x1_ASAP7_75t_L g7396 ( 
.A1(n_6143),
.A2(n_5951),
.B(n_5100),
.Y(n_7396)
);

NAND2xp5_ASAP7_75t_L g7397 ( 
.A(n_5303),
.B(n_5309),
.Y(n_7397)
);

AOI21x1_ASAP7_75t_L g7398 ( 
.A1(n_5641),
.A2(n_6084),
.B(n_6079),
.Y(n_7398)
);

AO31x2_ASAP7_75t_L g7399 ( 
.A1(n_5067),
.A2(n_5100),
.A3(n_5162),
.B(n_5140),
.Y(n_7399)
);

OA21x2_ASAP7_75t_L g7400 ( 
.A1(n_6065),
.A2(n_6084),
.B(n_6079),
.Y(n_7400)
);

NAND2xp5_ASAP7_75t_L g7401 ( 
.A(n_5309),
.B(n_5310),
.Y(n_7401)
);

INVx3_ASAP7_75t_L g7402 ( 
.A(n_4771),
.Y(n_7402)
);

NOR2xp33_ASAP7_75t_L g7403 ( 
.A(n_5850),
.B(n_5871),
.Y(n_7403)
);

CKINVDCx5p33_ASAP7_75t_R g7404 ( 
.A(n_5806),
.Y(n_7404)
);

AOI21xp5_ASAP7_75t_L g7405 ( 
.A1(n_5123),
.A2(n_5152),
.B(n_5124),
.Y(n_7405)
);

AOI21xp5_ASAP7_75t_L g7406 ( 
.A1(n_5123),
.A2(n_5152),
.B(n_5124),
.Y(n_7406)
);

AOI221xp5_ASAP7_75t_SL g7407 ( 
.A1(n_5542),
.A2(n_5589),
.B1(n_6234),
.B2(n_5853),
.C(n_6020),
.Y(n_7407)
);

OAI21x1_ASAP7_75t_L g7408 ( 
.A1(n_6143),
.A2(n_5951),
.B(n_5185),
.Y(n_7408)
);

BUFx2_ASAP7_75t_L g7409 ( 
.A(n_5686),
.Y(n_7409)
);

A2O1A1Ixp33_ASAP7_75t_L g7410 ( 
.A1(n_6218),
.A2(n_6232),
.B(n_6231),
.C(n_5651),
.Y(n_7410)
);

OAI22x1_ASAP7_75t_L g7411 ( 
.A1(n_6234),
.A2(n_5941),
.B1(n_5440),
.B2(n_5460),
.Y(n_7411)
);

OAI21x1_ASAP7_75t_L g7412 ( 
.A1(n_5951),
.A2(n_5185),
.B(n_5162),
.Y(n_7412)
);

OAI21x1_ASAP7_75t_L g7413 ( 
.A1(n_5162),
.A2(n_5197),
.B(n_5185),
.Y(n_7413)
);

OAI21x1_ASAP7_75t_L g7414 ( 
.A1(n_5197),
.A2(n_5252),
.B(n_5246),
.Y(n_7414)
);

AOI21x1_ASAP7_75t_L g7415 ( 
.A1(n_6085),
.A2(n_6108),
.B(n_6089),
.Y(n_7415)
);

NAND2xp5_ASAP7_75t_L g7416 ( 
.A(n_5310),
.B(n_5314),
.Y(n_7416)
);

AOI21xp5_ASAP7_75t_L g7417 ( 
.A1(n_5124),
.A2(n_5193),
.B(n_5152),
.Y(n_7417)
);

OAI21xp5_ASAP7_75t_L g7418 ( 
.A1(n_6206),
.A2(n_5853),
.B(n_5826),
.Y(n_7418)
);

NOR2x1_ASAP7_75t_SL g7419 ( 
.A(n_5124),
.B(n_5152),
.Y(n_7419)
);

AOI21x1_ASAP7_75t_L g7420 ( 
.A1(n_6085),
.A2(n_6108),
.B(n_6089),
.Y(n_7420)
);

NAND2xp5_ASAP7_75t_L g7421 ( 
.A(n_5314),
.B(n_5322),
.Y(n_7421)
);

NAND2xp5_ASAP7_75t_SL g7422 ( 
.A(n_5998),
.B(n_6070),
.Y(n_7422)
);

BUFx2_ASAP7_75t_L g7423 ( 
.A(n_5686),
.Y(n_7423)
);

AOI21x1_ASAP7_75t_L g7424 ( 
.A1(n_6026),
.A2(n_6173),
.B(n_6141),
.Y(n_7424)
);

AOI21xp5_ASAP7_75t_L g7425 ( 
.A1(n_5124),
.A2(n_5193),
.B(n_5152),
.Y(n_7425)
);

O2A1O1Ixp5_ASAP7_75t_L g7426 ( 
.A1(n_6182),
.A2(n_6065),
.B(n_5892),
.C(n_5246),
.Y(n_7426)
);

OAI211xp5_ASAP7_75t_SL g7427 ( 
.A1(n_5972),
.A2(n_5963),
.B(n_5845),
.C(n_6178),
.Y(n_7427)
);

NAND2x1_ASAP7_75t_L g7428 ( 
.A(n_4924),
.B(n_5265),
.Y(n_7428)
);

AOI21xp5_ASAP7_75t_L g7429 ( 
.A1(n_5152),
.A2(n_5242),
.B(n_5193),
.Y(n_7429)
);

AND2x4_ASAP7_75t_L g7430 ( 
.A(n_5197),
.B(n_5246),
.Y(n_7430)
);

AND2x4_ASAP7_75t_L g7431 ( 
.A(n_5256),
.B(n_5266),
.Y(n_7431)
);

AND2x4_ASAP7_75t_L g7432 ( 
.A(n_5266),
.B(n_5346),
.Y(n_7432)
);

OAI21xp5_ASAP7_75t_L g7433 ( 
.A1(n_5826),
.A2(n_6020),
.B(n_5575),
.Y(n_7433)
);

AOI22xp33_ASAP7_75t_SL g7434 ( 
.A1(n_6010),
.A2(n_6100),
.B1(n_5184),
.B2(n_5302),
.Y(n_7434)
);

AOI21xp5_ASAP7_75t_L g7435 ( 
.A1(n_5152),
.A2(n_5242),
.B(n_5193),
.Y(n_7435)
);

AOI21xp5_ASAP7_75t_L g7436 ( 
.A1(n_5193),
.A2(n_5255),
.B(n_5242),
.Y(n_7436)
);

INVx6_ASAP7_75t_L g7437 ( 
.A(n_5193),
.Y(n_7437)
);

NAND2xp5_ASAP7_75t_L g7438 ( 
.A(n_5244),
.B(n_5302),
.Y(n_7438)
);

AOI21xp5_ASAP7_75t_L g7439 ( 
.A1(n_5193),
.A2(n_5255),
.B(n_5242),
.Y(n_7439)
);

A2O1A1Ixp33_ASAP7_75t_L g7440 ( 
.A1(n_5635),
.A2(n_5735),
.B(n_5651),
.C(n_5857),
.Y(n_7440)
);

AOI21xp5_ASAP7_75t_L g7441 ( 
.A1(n_5242),
.A2(n_5255),
.B(n_6026),
.Y(n_7441)
);

INVx2_ASAP7_75t_L g7442 ( 
.A(n_5346),
.Y(n_7442)
);

NAND2xp5_ASAP7_75t_L g7443 ( 
.A(n_5244),
.B(n_5308),
.Y(n_7443)
);

OR2x2_ASAP7_75t_L g7444 ( 
.A(n_5707),
.B(n_5739),
.Y(n_7444)
);

OAI22xp5_ASAP7_75t_L g7445 ( 
.A1(n_6010),
.A2(n_6100),
.B1(n_6226),
.B2(n_5670),
.Y(n_7445)
);

BUFx3_ASAP7_75t_L g7446 ( 
.A(n_4771),
.Y(n_7446)
);

AOI21xp5_ASAP7_75t_L g7447 ( 
.A1(n_5242),
.A2(n_5255),
.B(n_4763),
.Y(n_7447)
);

INVx2_ASAP7_75t_L g7448 ( 
.A(n_5390),
.Y(n_7448)
);

AND2x6_ASAP7_75t_L g7449 ( 
.A(n_5255),
.B(n_5965),
.Y(n_7449)
);

NAND3xp33_ASAP7_75t_SL g7450 ( 
.A(n_6221),
.B(n_5728),
.C(n_6198),
.Y(n_7450)
);

AOI21x1_ASAP7_75t_L g7451 ( 
.A1(n_5904),
.A2(n_6038),
.B(n_5575),
.Y(n_7451)
);

AND2x4_ASAP7_75t_L g7452 ( 
.A(n_5417),
.B(n_5419),
.Y(n_7452)
);

BUFx6f_ASAP7_75t_L g7453 ( 
.A(n_5255),
.Y(n_7453)
);

OAI22xp5_ASAP7_75t_L g7454 ( 
.A1(n_6100),
.A2(n_5077),
.B1(n_6224),
.B2(n_5723),
.Y(n_7454)
);

NAND2xp5_ASAP7_75t_L g7455 ( 
.A(n_5308),
.B(n_5339),
.Y(n_7455)
);

OAI22xp5_ASAP7_75t_L g7456 ( 
.A1(n_5077),
.A2(n_6224),
.B1(n_5886),
.B2(n_5235),
.Y(n_7456)
);

OAI22xp5_ASAP7_75t_L g7457 ( 
.A1(n_5235),
.A2(n_5886),
.B1(n_6051),
.B2(n_6049),
.Y(n_7457)
);

NAND2xp5_ASAP7_75t_L g7458 ( 
.A(n_5308),
.B(n_5339),
.Y(n_7458)
);

AND2x4_ASAP7_75t_L g7459 ( 
.A(n_5489),
.B(n_5494),
.Y(n_7459)
);

INVx4_ASAP7_75t_L g7460 ( 
.A(n_5336),
.Y(n_7460)
);

NAND2xp5_ASAP7_75t_L g7461 ( 
.A(n_5339),
.B(n_4724),
.Y(n_7461)
);

A2O1A1Ixp33_ASAP7_75t_L g7462 ( 
.A1(n_5635),
.A2(n_5735),
.B(n_5969),
.C(n_4930),
.Y(n_7462)
);

NAND2xp5_ASAP7_75t_L g7463 ( 
.A(n_4724),
.B(n_4729),
.Y(n_7463)
);

OAI21xp5_ASAP7_75t_L g7464 ( 
.A1(n_5572),
.A2(n_5582),
.B(n_5579),
.Y(n_7464)
);

OA22x2_ASAP7_75t_L g7465 ( 
.A1(n_5998),
.A2(n_6070),
.B1(n_6076),
.B2(n_6075),
.Y(n_7465)
);

NAND2xp5_ASAP7_75t_L g7466 ( 
.A(n_4724),
.B(n_4729),
.Y(n_7466)
);

AND2x4_ASAP7_75t_L g7467 ( 
.A(n_5494),
.B(n_5495),
.Y(n_7467)
);

AO31x2_ASAP7_75t_L g7468 ( 
.A1(n_5495),
.A2(n_5499),
.A3(n_5505),
.B(n_5496),
.Y(n_7468)
);

BUFx6f_ASAP7_75t_L g7469 ( 
.A(n_5752),
.Y(n_7469)
);

AOI21xp5_ASAP7_75t_L g7470 ( 
.A1(n_4733),
.A2(n_5037),
.B(n_4763),
.Y(n_7470)
);

INVx2_ASAP7_75t_L g7471 ( 
.A(n_5499),
.Y(n_7471)
);

OR2x2_ASAP7_75t_L g7472 ( 
.A(n_5707),
.B(n_5739),
.Y(n_7472)
);

OAI21xp5_ASAP7_75t_L g7473 ( 
.A1(n_5572),
.A2(n_5582),
.B(n_5579),
.Y(n_7473)
);

NAND2xp5_ASAP7_75t_L g7474 ( 
.A(n_4729),
.B(n_4735),
.Y(n_7474)
);

AND2x2_ASAP7_75t_L g7475 ( 
.A(n_5505),
.B(n_5511),
.Y(n_7475)
);

OAI21x1_ASAP7_75t_SL g7476 ( 
.A1(n_6055),
.A2(n_6060),
.B(n_6058),
.Y(n_7476)
);

NAND2xp5_ASAP7_75t_L g7477 ( 
.A(n_4735),
.B(n_4801),
.Y(n_7477)
);

AOI22xp33_ASAP7_75t_L g7478 ( 
.A1(n_6196),
.A2(n_5514),
.B1(n_5987),
.B2(n_5881),
.Y(n_7478)
);

OA22x2_ASAP7_75t_L g7479 ( 
.A1(n_6075),
.A2(n_6076),
.B1(n_5686),
.B2(n_5965),
.Y(n_7479)
);

BUFx2_ASAP7_75t_L g7480 ( 
.A(n_5686),
.Y(n_7480)
);

AO21x2_ASAP7_75t_L g7481 ( 
.A1(n_5941),
.A2(n_5585),
.B(n_5584),
.Y(n_7481)
);

INVx2_ASAP7_75t_L g7482 ( 
.A(n_5511),
.Y(n_7482)
);

INVxp67_ASAP7_75t_L g7483 ( 
.A(n_5844),
.Y(n_7483)
);

CKINVDCx5p33_ASAP7_75t_R g7484 ( 
.A(n_5898),
.Y(n_7484)
);

OAI21x1_ASAP7_75t_SL g7485 ( 
.A1(n_6058),
.A2(n_6071),
.B(n_6060),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_L g7486 ( 
.A(n_4735),
.B(n_4801),
.Y(n_7486)
);

OAI21xp5_ASAP7_75t_L g7487 ( 
.A1(n_5584),
.A2(n_5593),
.B(n_5585),
.Y(n_7487)
);

A2O1A1Ixp33_ASAP7_75t_L g7488 ( 
.A1(n_5969),
.A2(n_4930),
.B(n_4985),
.C(n_4960),
.Y(n_7488)
);

BUFx6f_ASAP7_75t_L g7489 ( 
.A(n_5752),
.Y(n_7489)
);

NAND2x1p5_ASAP7_75t_L g7490 ( 
.A(n_5839),
.B(n_5037),
.Y(n_7490)
);

AND2x4_ASAP7_75t_L g7491 ( 
.A(n_5553),
.B(n_5566),
.Y(n_7491)
);

NAND2xp5_ASAP7_75t_L g7492 ( 
.A(n_4801),
.B(n_4905),
.Y(n_7492)
);

OAI22xp5_ASAP7_75t_L g7493 ( 
.A1(n_5235),
.A2(n_5886),
.B1(n_6073),
.B2(n_6071),
.Y(n_7493)
);

OAI21xp5_ASAP7_75t_L g7494 ( 
.A1(n_5593),
.A2(n_5604),
.B(n_5599),
.Y(n_7494)
);

AOI21xp5_ASAP7_75t_L g7495 ( 
.A1(n_5037),
.A2(n_5815),
.B(n_5337),
.Y(n_7495)
);

OAI21xp5_ASAP7_75t_L g7496 ( 
.A1(n_5599),
.A2(n_5605),
.B(n_5604),
.Y(n_7496)
);

INVx3_ASAP7_75t_L g7497 ( 
.A(n_4928),
.Y(n_7497)
);

AOI21xp5_ASAP7_75t_L g7498 ( 
.A1(n_5037),
.A2(n_5815),
.B(n_5337),
.Y(n_7498)
);

AOI22xp33_ASAP7_75t_L g7499 ( 
.A1(n_5881),
.A2(n_6109),
.B1(n_6223),
.B2(n_5987),
.Y(n_7499)
);

AOI21xp5_ASAP7_75t_L g7500 ( 
.A1(n_5337),
.A2(n_5815),
.B(n_5969),
.Y(n_7500)
);

OAI22x1_ASAP7_75t_L g7501 ( 
.A1(n_5409),
.A2(n_5460),
.B1(n_5600),
.B2(n_5440),
.Y(n_7501)
);

OAI21x1_ASAP7_75t_L g7502 ( 
.A1(n_5553),
.A2(n_5588),
.B(n_5566),
.Y(n_7502)
);

OAI21xp5_ASAP7_75t_L g7503 ( 
.A1(n_5605),
.A2(n_5620),
.B(n_5609),
.Y(n_7503)
);

OAI21xp5_ASAP7_75t_L g7504 ( 
.A1(n_5609),
.A2(n_5621),
.B(n_5620),
.Y(n_7504)
);

AOI21xp5_ASAP7_75t_L g7505 ( 
.A1(n_5337),
.A2(n_5815),
.B(n_6212),
.Y(n_7505)
);

OAI21x1_ASAP7_75t_L g7506 ( 
.A1(n_5553),
.A2(n_5588),
.B(n_5566),
.Y(n_7506)
);

AOI21xp5_ASAP7_75t_L g7507 ( 
.A1(n_6212),
.A2(n_5672),
.B(n_5664),
.Y(n_7507)
);

AOI21xp5_ASAP7_75t_L g7508 ( 
.A1(n_6212),
.A2(n_5691),
.B(n_4737),
.Y(n_7508)
);

OAI21x1_ASAP7_75t_L g7509 ( 
.A1(n_5588),
.A2(n_5622),
.B(n_5602),
.Y(n_7509)
);

AOI21xp5_ASAP7_75t_SL g7510 ( 
.A1(n_5840),
.A2(n_6062),
.B(n_6046),
.Y(n_7510)
);

AND2x2_ASAP7_75t_L g7511 ( 
.A(n_5602),
.B(n_5622),
.Y(n_7511)
);

AND2x2_ASAP7_75t_L g7512 ( 
.A(n_5661),
.B(n_5673),
.Y(n_7512)
);

OAI22x1_ASAP7_75t_L g7513 ( 
.A1(n_5409),
.A2(n_5600),
.B1(n_5895),
.B2(n_5639),
.Y(n_7513)
);

AND2x2_ASAP7_75t_L g7514 ( 
.A(n_5661),
.B(n_5673),
.Y(n_7514)
);

INVx5_ASAP7_75t_L g7515 ( 
.A(n_4924),
.Y(n_7515)
);

INVx1_ASAP7_75t_SL g7516 ( 
.A(n_5834),
.Y(n_7516)
);

AOI21x1_ASAP7_75t_L g7517 ( 
.A1(n_5621),
.A2(n_5629),
.B(n_5623),
.Y(n_7517)
);

NAND2xp5_ASAP7_75t_L g7518 ( 
.A(n_4905),
.B(n_4917),
.Y(n_7518)
);

BUFx2_ASAP7_75t_L g7519 ( 
.A(n_5686),
.Y(n_7519)
);

NAND2xp5_ASAP7_75t_L g7520 ( 
.A(n_4905),
.B(n_4917),
.Y(n_7520)
);

AOI21xp5_ASAP7_75t_L g7521 ( 
.A1(n_4730),
.A2(n_4737),
.B(n_4732),
.Y(n_7521)
);

AO31x2_ASAP7_75t_L g7522 ( 
.A1(n_5680),
.A2(n_5693),
.A3(n_5763),
.B(n_5732),
.Y(n_7522)
);

OAI21x1_ASAP7_75t_L g7523 ( 
.A1(n_5680),
.A2(n_5732),
.B(n_5693),
.Y(n_7523)
);

A2O1A1Ixp33_ASAP7_75t_L g7524 ( 
.A1(n_4930),
.A2(n_4960),
.B(n_5057),
.C(n_4985),
.Y(n_7524)
);

CKINVDCx5p33_ASAP7_75t_R g7525 ( 
.A(n_6011),
.Y(n_7525)
);

NAND2xp5_ASAP7_75t_L g7526 ( 
.A(n_5948),
.B(n_5968),
.Y(n_7526)
);

OAI21xp5_ASAP7_75t_L g7527 ( 
.A1(n_5623),
.A2(n_5637),
.B(n_5629),
.Y(n_7527)
);

NAND2xp5_ASAP7_75t_L g7528 ( 
.A(n_5948),
.B(n_5968),
.Y(n_7528)
);

OAI21x1_ASAP7_75t_L g7529 ( 
.A1(n_5763),
.A2(n_5788),
.B(n_5773),
.Y(n_7529)
);

AOI21xp5_ASAP7_75t_L g7530 ( 
.A1(n_4732),
.A2(n_5839),
.B(n_5686),
.Y(n_7530)
);

INVx4_ASAP7_75t_L g7531 ( 
.A(n_5336),
.Y(n_7531)
);

AND2x2_ASAP7_75t_L g7532 ( 
.A(n_5773),
.B(n_5788),
.Y(n_7532)
);

AOI21xp33_ASAP7_75t_L g7533 ( 
.A1(n_5929),
.A2(n_5942),
.B(n_5656),
.Y(n_7533)
);

OAI21xp33_ASAP7_75t_L g7534 ( 
.A1(n_5929),
.A2(n_5942),
.B(n_6073),
.Y(n_7534)
);

OAI21xp5_ASAP7_75t_L g7535 ( 
.A1(n_5637),
.A2(n_5657),
.B(n_5656),
.Y(n_7535)
);

OR2x6_ASAP7_75t_L g7536 ( 
.A(n_4924),
.B(n_5265),
.Y(n_7536)
);

NAND2xp5_ASAP7_75t_L g7537 ( 
.A(n_5978),
.B(n_5986),
.Y(n_7537)
);

AOI21xp33_ASAP7_75t_L g7538 ( 
.A1(n_5657),
.A2(n_5666),
.B(n_5665),
.Y(n_7538)
);

INVx3_ASAP7_75t_L g7539 ( 
.A(n_4928),
.Y(n_7539)
);

OAI21x1_ASAP7_75t_L g7540 ( 
.A1(n_5788),
.A2(n_5812),
.B(n_5811),
.Y(n_7540)
);

AOI21xp5_ASAP7_75t_L g7541 ( 
.A1(n_4732),
.A2(n_5839),
.B(n_6175),
.Y(n_7541)
);

AOI21x1_ASAP7_75t_L g7542 ( 
.A1(n_5665),
.A2(n_5678),
.B(n_5666),
.Y(n_7542)
);

NAND2xp5_ASAP7_75t_L g7543 ( 
.A(n_5978),
.B(n_5986),
.Y(n_7543)
);

OAI21x1_ASAP7_75t_L g7544 ( 
.A1(n_5811),
.A2(n_5827),
.B(n_5812),
.Y(n_7544)
);

OR2x6_ASAP7_75t_L g7545 ( 
.A(n_4924),
.B(n_5265),
.Y(n_7545)
);

NAND2xp5_ASAP7_75t_L g7546 ( 
.A(n_5993),
.B(n_6001),
.Y(n_7546)
);

AOI21x1_ASAP7_75t_L g7547 ( 
.A1(n_5678),
.A2(n_5683),
.B(n_5681),
.Y(n_7547)
);

OAI21xp33_ASAP7_75t_L g7548 ( 
.A1(n_6091),
.A2(n_6098),
.B(n_6096),
.Y(n_7548)
);

BUFx3_ASAP7_75t_L g7549 ( 
.A(n_4928),
.Y(n_7549)
);

A2O1A1Ixp33_ASAP7_75t_L g7550 ( 
.A1(n_4960),
.A2(n_4985),
.B(n_5343),
.C(n_5057),
.Y(n_7550)
);

AOI21x1_ASAP7_75t_L g7551 ( 
.A1(n_5681),
.A2(n_5690),
.B(n_5683),
.Y(n_7551)
);

NAND2xp5_ASAP7_75t_L g7552 ( 
.A(n_5993),
.B(n_6001),
.Y(n_7552)
);

NAND2xp5_ASAP7_75t_SL g7553 ( 
.A(n_6075),
.B(n_6076),
.Y(n_7553)
);

NAND2xp5_ASAP7_75t_L g7554 ( 
.A(n_6003),
.B(n_6022),
.Y(n_7554)
);

INVx1_ASAP7_75t_L g7555 ( 
.A(n_6176),
.Y(n_7555)
);

BUFx4_ASAP7_75t_SL g7556 ( 
.A(n_6082),
.Y(n_7556)
);

NAND2xp5_ASAP7_75t_L g7557 ( 
.A(n_6003),
.B(n_6022),
.Y(n_7557)
);

NAND2xp5_ASAP7_75t_L g7558 ( 
.A(n_5690),
.B(n_5695),
.Y(n_7558)
);

OAI22x1_ASAP7_75t_L g7559 ( 
.A1(n_5639),
.A2(n_5895),
.B1(n_5914),
.B2(n_6183),
.Y(n_7559)
);

OAI21x1_ASAP7_75t_L g7560 ( 
.A1(n_5914),
.A2(n_6093),
.B(n_6028),
.Y(n_7560)
);

OAI21x1_ASAP7_75t_L g7561 ( 
.A1(n_6028),
.A2(n_6093),
.B(n_5702),
.Y(n_7561)
);

AO21x1_ASAP7_75t_L g7562 ( 
.A1(n_5695),
.A2(n_5712),
.B(n_5702),
.Y(n_7562)
);

AOI21xp5_ASAP7_75t_L g7563 ( 
.A1(n_5839),
.A2(n_6227),
.B(n_6175),
.Y(n_7563)
);

OAI21x1_ASAP7_75t_L g7564 ( 
.A1(n_6093),
.A2(n_5730),
.B(n_5714),
.Y(n_7564)
);

OAI21x1_ASAP7_75t_L g7565 ( 
.A1(n_5730),
.A2(n_5768),
.B(n_5744),
.Y(n_7565)
);

AND2x2_ASAP7_75t_L g7566 ( 
.A(n_5953),
.B(n_5992),
.Y(n_7566)
);

INVx1_ASAP7_75t_SL g7567 ( 
.A(n_5834),
.Y(n_7567)
);

AOI21xp5_ASAP7_75t_L g7568 ( 
.A1(n_5839),
.A2(n_6227),
.B(n_6175),
.Y(n_7568)
);

AND2x4_ASAP7_75t_L g7569 ( 
.A(n_5953),
.B(n_5992),
.Y(n_7569)
);

INVx1_ASAP7_75t_L g7570 ( 
.A(n_6176),
.Y(n_7570)
);

OAI21x1_ASAP7_75t_SL g7571 ( 
.A1(n_6091),
.A2(n_6098),
.B(n_6096),
.Y(n_7571)
);

AOI21x1_ASAP7_75t_L g7572 ( 
.A1(n_5778),
.A2(n_5793),
.B(n_5789),
.Y(n_7572)
);

NAND2xp5_ASAP7_75t_SL g7573 ( 
.A(n_6075),
.B(n_6076),
.Y(n_7573)
);

AOI21xp5_ASAP7_75t_L g7574 ( 
.A1(n_5839),
.A2(n_6227),
.B(n_6175),
.Y(n_7574)
);

OAI21xp5_ASAP7_75t_L g7575 ( 
.A1(n_5778),
.A2(n_5793),
.B(n_5789),
.Y(n_7575)
);

AOI21xp5_ASAP7_75t_L g7576 ( 
.A1(n_5839),
.A2(n_6227),
.B(n_6175),
.Y(n_7576)
);

OAI22xp5_ASAP7_75t_L g7577 ( 
.A1(n_6102),
.A2(n_6253),
.B1(n_6252),
.B2(n_6250),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_6183),
.Y(n_7578)
);

OAI21xp5_ASAP7_75t_L g7579 ( 
.A1(n_5820),
.A2(n_5832),
.B(n_5828),
.Y(n_7579)
);

OAI21x1_ASAP7_75t_L g7580 ( 
.A1(n_5843),
.A2(n_5860),
.B(n_5858),
.Y(n_7580)
);

BUFx10_ASAP7_75t_L g7581 ( 
.A(n_5265),
.Y(n_7581)
);

AOI21x1_ASAP7_75t_SL g7582 ( 
.A1(n_5581),
.A2(n_5875),
.B(n_5790),
.Y(n_7582)
);

NAND2xp33_ASAP7_75t_L g7583 ( 
.A(n_5373),
.B(n_5148),
.Y(n_7583)
);

NAND2xp5_ASAP7_75t_L g7584 ( 
.A(n_5861),
.B(n_5862),
.Y(n_7584)
);

NAND2xp5_ASAP7_75t_SL g7585 ( 
.A(n_5934),
.B(n_5752),
.Y(n_7585)
);

AOI21xp5_ASAP7_75t_L g7586 ( 
.A1(n_6175),
.A2(n_6227),
.B(n_5028),
.Y(n_7586)
);

AND2x2_ASAP7_75t_L g7587 ( 
.A(n_5953),
.B(n_5992),
.Y(n_7587)
);

OR2x6_ASAP7_75t_L g7588 ( 
.A(n_5057),
.B(n_5343),
.Y(n_7588)
);

OAI21x1_ASAP7_75t_L g7589 ( 
.A1(n_5861),
.A2(n_5866),
.B(n_5862),
.Y(n_7589)
);

BUFx6f_ASAP7_75t_L g7590 ( 
.A(n_5752),
.Y(n_7590)
);

NAND3xp33_ASAP7_75t_L g7591 ( 
.A(n_6102),
.B(n_6106),
.C(n_6104),
.Y(n_7591)
);

AOI21xp5_ASAP7_75t_L g7592 ( 
.A1(n_6175),
.A2(n_6227),
.B(n_5028),
.Y(n_7592)
);

INVx1_ASAP7_75t_L g7593 ( 
.A(n_6205),
.Y(n_7593)
);

OAI21x1_ASAP7_75t_L g7594 ( 
.A1(n_5866),
.A2(n_5878),
.B(n_5868),
.Y(n_7594)
);

AOI21xp5_ASAP7_75t_L g7595 ( 
.A1(n_5028),
.A2(n_5286),
.B(n_5896),
.Y(n_7595)
);

AOI21xp5_ASAP7_75t_L g7596 ( 
.A1(n_5028),
.A2(n_5940),
.B(n_5917),
.Y(n_7596)
);

INVx1_ASAP7_75t_L g7597 ( 
.A(n_6213),
.Y(n_7597)
);

OAI21xp5_ASAP7_75t_L g7598 ( 
.A1(n_5884),
.A2(n_6202),
.B(n_5999),
.Y(n_7598)
);

INVx1_ASAP7_75t_SL g7599 ( 
.A(n_5834),
.Y(n_7599)
);

OAI21x1_ASAP7_75t_L g7600 ( 
.A1(n_6202),
.A2(n_5945),
.B(n_5943),
.Y(n_7600)
);

NAND2xp5_ASAP7_75t_L g7601 ( 
.A(n_6149),
.B(n_6160),
.Y(n_7601)
);

AO31x2_ASAP7_75t_L g7602 ( 
.A1(n_6213),
.A2(n_6238),
.A3(n_6220),
.B(n_5994),
.Y(n_7602)
);

AOI21xp5_ASAP7_75t_SL g7603 ( 
.A1(n_5840),
.A2(n_6062),
.B(n_6046),
.Y(n_7603)
);

OAI21xp5_ASAP7_75t_L g7604 ( 
.A1(n_6202),
.A2(n_5999),
.B(n_5785),
.Y(n_7604)
);

NAND2xp5_ASAP7_75t_SL g7605 ( 
.A(n_5934),
.B(n_5752),
.Y(n_7605)
);

OAI21x1_ASAP7_75t_L g7606 ( 
.A1(n_5943),
.A2(n_5960),
.B(n_5945),
.Y(n_7606)
);

NAND3xp33_ASAP7_75t_L g7607 ( 
.A(n_6104),
.B(n_6253),
.C(n_6252),
.Y(n_7607)
);

OAI22x1_ASAP7_75t_L g7608 ( 
.A1(n_6220),
.A2(n_6238),
.B1(n_5999),
.B2(n_5946),
.Y(n_7608)
);

AOI21xp5_ASAP7_75t_L g7609 ( 
.A1(n_5028),
.A2(n_5950),
.B(n_6016),
.Y(n_7609)
);

BUFx2_ASAP7_75t_L g7610 ( 
.A(n_5752),
.Y(n_7610)
);

AOI21xp5_ASAP7_75t_SL g7611 ( 
.A1(n_5840),
.A2(n_6062),
.B(n_6025),
.Y(n_7611)
);

AOI21xp5_ASAP7_75t_L g7612 ( 
.A1(n_5961),
.A2(n_5970),
.B(n_6000),
.Y(n_7612)
);

CKINVDCx20_ASAP7_75t_R g7613 ( 
.A(n_5881),
.Y(n_7613)
);

INVx2_ASAP7_75t_SL g7614 ( 
.A(n_5792),
.Y(n_7614)
);

OAI21x1_ASAP7_75t_L g7615 ( 
.A1(n_5960),
.A2(n_5974),
.B(n_6014),
.Y(n_7615)
);

AOI21xp5_ASAP7_75t_L g7616 ( 
.A1(n_6013),
.A2(n_5974),
.B(n_5976),
.Y(n_7616)
);

NAND2xp5_ASAP7_75t_SL g7617 ( 
.A(n_5934),
.B(n_5792),
.Y(n_7617)
);

OAI21x1_ASAP7_75t_L g7618 ( 
.A1(n_5976),
.A2(n_5983),
.B(n_5994),
.Y(n_7618)
);

NAND2xp5_ASAP7_75t_L g7619 ( 
.A(n_6222),
.B(n_5983),
.Y(n_7619)
);

NAND2xp5_ASAP7_75t_L g7620 ( 
.A(n_6002),
.B(n_6014),
.Y(n_7620)
);

OAI21x1_ASAP7_75t_L g7621 ( 
.A1(n_6002),
.A2(n_6059),
.B(n_6113),
.Y(n_7621)
);

INVx3_ASAP7_75t_SL g7622 ( 
.A(n_5336),
.Y(n_7622)
);

INVx1_ASAP7_75t_L g7623 ( 
.A(n_5792),
.Y(n_7623)
);

HB1xp67_ASAP7_75t_L g7624 ( 
.A(n_6115),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_5792),
.Y(n_7625)
);

OR2x6_ASAP7_75t_L g7626 ( 
.A(n_5343),
.B(n_5805),
.Y(n_7626)
);

NAND2xp5_ASAP7_75t_L g7627 ( 
.A(n_6113),
.B(n_6118),
.Y(n_7627)
);

OAI21x1_ASAP7_75t_L g7628 ( 
.A1(n_6118),
.A2(n_6250),
.B(n_6132),
.Y(n_7628)
);

NAND2xp5_ASAP7_75t_L g7629 ( 
.A(n_6132),
.B(n_6136),
.Y(n_7629)
);

AND2x4_ASAP7_75t_L g7630 ( 
.A(n_4928),
.B(n_5104),
.Y(n_7630)
);

BUFx2_ASAP7_75t_L g7631 ( 
.A(n_5792),
.Y(n_7631)
);

INVx1_ASAP7_75t_L g7632 ( 
.A(n_5792),
.Y(n_7632)
);

OAI21x1_ASAP7_75t_L g7633 ( 
.A1(n_6136),
.A2(n_6174),
.B(n_6246),
.Y(n_7633)
);

NAND2xp5_ASAP7_75t_L g7634 ( 
.A(n_6147),
.B(n_6163),
.Y(n_7634)
);

NAND2xp5_ASAP7_75t_L g7635 ( 
.A(n_6147),
.B(n_6163),
.Y(n_7635)
);

NAND3xp33_ASAP7_75t_L g7636 ( 
.A(n_6164),
.B(n_6170),
.C(n_6246),
.Y(n_7636)
);

OAI21x1_ASAP7_75t_L g7637 ( 
.A1(n_6164),
.A2(n_6216),
.B(n_6245),
.Y(n_7637)
);

NOR2x1_ASAP7_75t_SL g7638 ( 
.A(n_5805),
.B(n_5825),
.Y(n_7638)
);

AOI21xp5_ASAP7_75t_L g7639 ( 
.A1(n_6168),
.A2(n_6211),
.B(n_6245),
.Y(n_7639)
);

OAI21xp5_ASAP7_75t_L g7640 ( 
.A1(n_5781),
.A2(n_6174),
.B(n_6240),
.Y(n_7640)
);

NAND2xp5_ASAP7_75t_L g7641 ( 
.A(n_6168),
.B(n_6170),
.Y(n_7641)
);

OA22x2_ASAP7_75t_L g7642 ( 
.A1(n_5965),
.A2(n_5790),
.B1(n_5875),
.B2(n_5581),
.Y(n_7642)
);

OAI21x1_ASAP7_75t_L g7643 ( 
.A1(n_6172),
.A2(n_6203),
.B(n_6240),
.Y(n_7643)
);

INVx1_ASAP7_75t_SL g7644 ( 
.A(n_6086),
.Y(n_7644)
);

NAND2xp5_ASAP7_75t_L g7645 ( 
.A(n_6172),
.B(n_6190),
.Y(n_7645)
);

NOR2xp33_ASAP7_75t_L g7646 ( 
.A(n_5934),
.B(n_5792),
.Y(n_7646)
);

INVx2_ASAP7_75t_L g7647 ( 
.A(n_5796),
.Y(n_7647)
);

AOI21xp5_ASAP7_75t_L g7648 ( 
.A1(n_6190),
.A2(n_6211),
.B(n_6217),
.Y(n_7648)
);

AND2x4_ASAP7_75t_L g7649 ( 
.A(n_5104),
.B(n_5225),
.Y(n_7649)
);

OAI21xp5_ASAP7_75t_L g7650 ( 
.A1(n_6193),
.A2(n_6217),
.B(n_6216),
.Y(n_7650)
);

OAI21x1_ASAP7_75t_L g7651 ( 
.A1(n_6193),
.A2(n_6208),
.B(n_6203),
.Y(n_7651)
);

OAI21x1_ASAP7_75t_L g7652 ( 
.A1(n_6197),
.A2(n_6208),
.B(n_6130),
.Y(n_7652)
);

INVx1_ASAP7_75t_L g7653 ( 
.A(n_5796),
.Y(n_7653)
);

OAI21xp5_ASAP7_75t_L g7654 ( 
.A1(n_6086),
.A2(n_5734),
.B(n_5737),
.Y(n_7654)
);

AOI21xp5_ASAP7_75t_L g7655 ( 
.A1(n_5805),
.A2(n_5825),
.B(n_6062),
.Y(n_7655)
);

OAI21x1_ASAP7_75t_L g7656 ( 
.A1(n_5946),
.A2(n_6247),
.B(n_5740),
.Y(n_7656)
);

OAI21x1_ASAP7_75t_L g7657 ( 
.A1(n_5946),
.A2(n_5373),
.B(n_5774),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_5796),
.Y(n_7658)
);

NAND2xp5_ASAP7_75t_L g7659 ( 
.A(n_5934),
.B(n_5796),
.Y(n_7659)
);

AOI21xp5_ASAP7_75t_L g7660 ( 
.A1(n_5825),
.A2(n_5796),
.B(n_5934),
.Y(n_7660)
);

A2O1A1Ixp33_ASAP7_75t_L g7661 ( 
.A1(n_5745),
.A2(n_6087),
.B(n_6069),
.C(n_5938),
.Y(n_7661)
);

NOR2xp33_ASAP7_75t_L g7662 ( 
.A(n_5934),
.B(n_5796),
.Y(n_7662)
);

NAND2xp5_ASAP7_75t_L g7663 ( 
.A(n_5796),
.B(n_5597),
.Y(n_7663)
);

OAI21xp5_ASAP7_75t_L g7664 ( 
.A1(n_5965),
.A2(n_6138),
.B(n_6137),
.Y(n_7664)
);

INVx2_ASAP7_75t_L g7665 ( 
.A(n_5104),
.Y(n_7665)
);

NAND2xp5_ASAP7_75t_L g7666 ( 
.A(n_5307),
.B(n_5640),
.Y(n_7666)
);

NOR2xp67_ASAP7_75t_L g7667 ( 
.A(n_5104),
.B(n_5513),
.Y(n_7667)
);

OAI21xp5_ASAP7_75t_L g7668 ( 
.A1(n_6137),
.A2(n_6138),
.B(n_5513),
.Y(n_7668)
);

NAND2xp5_ASAP7_75t_L g7669 ( 
.A(n_5307),
.B(n_5640),
.Y(n_7669)
);

INVx3_ASAP7_75t_L g7670 ( 
.A(n_5225),
.Y(n_7670)
);

OAI22x1_ASAP7_75t_L g7671 ( 
.A1(n_5225),
.A2(n_5513),
.B1(n_6138),
.B2(n_6137),
.Y(n_7671)
);

OAI21x1_ASAP7_75t_L g7672 ( 
.A1(n_5373),
.A2(n_5838),
.B(n_5954),
.Y(n_7672)
);

A2O1A1Ixp33_ASAP7_75t_L g7673 ( 
.A1(n_5753),
.A2(n_5823),
.B(n_5869),
.C(n_6036),
.Y(n_7673)
);

AOI21xp33_ASAP7_75t_L g7674 ( 
.A1(n_6025),
.A2(n_6046),
.B(n_6137),
.Y(n_7674)
);

AOI21x1_ASAP7_75t_SL g7675 ( 
.A1(n_5225),
.A2(n_5513),
.B(n_4934),
.Y(n_7675)
);

OAI21x1_ASAP7_75t_L g7676 ( 
.A1(n_5373),
.A2(n_5822),
.B(n_5877),
.Y(n_7676)
);

OAI21xp5_ASAP7_75t_L g7677 ( 
.A1(n_6138),
.A2(n_6025),
.B(n_5770),
.Y(n_7677)
);

OAI21xp5_ASAP7_75t_L g7678 ( 
.A1(n_5772),
.A2(n_5804),
.B(n_5851),
.Y(n_7678)
);

OAI21x1_ASAP7_75t_L g7679 ( 
.A1(n_5373),
.A2(n_5800),
.B(n_6035),
.Y(n_7679)
);

NAND2xp5_ASAP7_75t_L g7680 ( 
.A(n_5307),
.B(n_5640),
.Y(n_7680)
);

CKINVDCx6p67_ASAP7_75t_R g7681 ( 
.A(n_4832),
.Y(n_7681)
);

AOI21xp5_ASAP7_75t_L g7682 ( 
.A1(n_5307),
.A2(n_5559),
.B(n_5640),
.Y(n_7682)
);

OAI21xp5_ASAP7_75t_L g7683 ( 
.A1(n_5856),
.A2(n_5988),
.B(n_5885),
.Y(n_7683)
);

AOI21xp5_ASAP7_75t_L g7684 ( 
.A1(n_6352),
.A2(n_5606),
.B(n_5640),
.Y(n_7684)
);

OAI21xp5_ASAP7_75t_L g7685 ( 
.A1(n_6364),
.A2(n_5989),
.B(n_5874),
.Y(n_7685)
);

INVx5_ASAP7_75t_L g7686 ( 
.A(n_6602),
.Y(n_7686)
);

NOR2xp33_ASAP7_75t_L g7687 ( 
.A(n_6527),
.B(n_5597),
.Y(n_7687)
);

NAND2xp5_ASAP7_75t_L g7688 ( 
.A(n_6996),
.B(n_5597),
.Y(n_7688)
);

AO21x2_ASAP7_75t_L g7689 ( 
.A1(n_6351),
.A2(n_5373),
.B(n_5606),
.Y(n_7689)
);

AOI21xp5_ASAP7_75t_L g7690 ( 
.A1(n_6352),
.A2(n_5597),
.B(n_5640),
.Y(n_7690)
);

NAND2xp5_ASAP7_75t_L g7691 ( 
.A(n_6996),
.B(n_5597),
.Y(n_7691)
);

OAI21x1_ASAP7_75t_L g7692 ( 
.A1(n_6747),
.A2(n_5373),
.B(n_5336),
.Y(n_7692)
);

CKINVDCx5p33_ASAP7_75t_R g7693 ( 
.A(n_7556),
.Y(n_7693)
);

AOI21xp5_ASAP7_75t_L g7694 ( 
.A1(n_6391),
.A2(n_5597),
.B(n_5640),
.Y(n_7694)
);

INVx3_ASAP7_75t_L g7695 ( 
.A(n_6854),
.Y(n_7695)
);

INVxp67_ASAP7_75t_L g7696 ( 
.A(n_6723),
.Y(n_7696)
);

AOI22xp33_ASAP7_75t_L g7697 ( 
.A1(n_6696),
.A2(n_5987),
.B1(n_5881),
.B2(n_6109),
.Y(n_7697)
);

AOI21xp5_ASAP7_75t_L g7698 ( 
.A1(n_6391),
.A2(n_5570),
.B(n_5606),
.Y(n_7698)
);

O2A1O1Ixp5_ASAP7_75t_SL g7699 ( 
.A1(n_6781),
.A2(n_4934),
.B(n_5849),
.C(n_5564),
.Y(n_7699)
);

NAND2xp5_ASAP7_75t_L g7700 ( 
.A(n_6977),
.B(n_5570),
.Y(n_7700)
);

A2O1A1Ixp33_ASAP7_75t_L g7701 ( 
.A1(n_6364),
.A2(n_5910),
.B(n_5307),
.C(n_5570),
.Y(n_7701)
);

INVx2_ASAP7_75t_L g7702 ( 
.A(n_7395),
.Y(n_7702)
);

NAND2xp5_ASAP7_75t_L g7703 ( 
.A(n_6977),
.B(n_5570),
.Y(n_7703)
);

NAND2xp5_ASAP7_75t_L g7704 ( 
.A(n_6436),
.B(n_5570),
.Y(n_7704)
);

OAI21x1_ASAP7_75t_SL g7705 ( 
.A1(n_7216),
.A2(n_5564),
.B(n_5421),
.Y(n_7705)
);

BUFx6f_ASAP7_75t_L g7706 ( 
.A(n_6578),
.Y(n_7706)
);

AOI21x1_ASAP7_75t_L g7707 ( 
.A1(n_6265),
.A2(n_5849),
.B(n_5421),
.Y(n_7707)
);

AOI21x1_ASAP7_75t_L g7708 ( 
.A1(n_6265),
.A2(n_6502),
.B(n_6685),
.Y(n_7708)
);

NAND2xp5_ASAP7_75t_L g7709 ( 
.A(n_6436),
.B(n_5606),
.Y(n_7709)
);

OAI21xp5_ASAP7_75t_L g7710 ( 
.A1(n_6527),
.A2(n_5148),
.B(n_5925),
.Y(n_7710)
);

OR2x2_ASAP7_75t_L g7711 ( 
.A(n_6934),
.B(n_6979),
.Y(n_7711)
);

AOI21xp33_ASAP7_75t_L g7712 ( 
.A1(n_6304),
.A2(n_6459),
.B(n_6696),
.Y(n_7712)
);

AOI21xp5_ASAP7_75t_L g7713 ( 
.A1(n_6401),
.A2(n_5606),
.B(n_5526),
.Y(n_7713)
);

INVx5_ASAP7_75t_L g7714 ( 
.A(n_6602),
.Y(n_7714)
);

BUFx3_ASAP7_75t_L g7715 ( 
.A(n_7449),
.Y(n_7715)
);

AOI22xp5_ASAP7_75t_L g7716 ( 
.A1(n_6459),
.A2(n_6642),
.B1(n_6748),
.B2(n_6693),
.Y(n_7716)
);

AOI21xp5_ASAP7_75t_SL g7717 ( 
.A1(n_6745),
.A2(n_6233),
.B(n_5559),
.Y(n_7717)
);

BUFx4f_ASAP7_75t_L g7718 ( 
.A(n_6531),
.Y(n_7718)
);

NAND2xp5_ASAP7_75t_SL g7719 ( 
.A(n_6704),
.B(n_5559),
.Y(n_7719)
);

AOI22xp5_ASAP7_75t_L g7720 ( 
.A1(n_6459),
.A2(n_5336),
.B1(n_5373),
.B2(n_5148),
.Y(n_7720)
);

OAI21x1_ASAP7_75t_L g7721 ( 
.A1(n_6747),
.A2(n_5148),
.B(n_5454),
.Y(n_7721)
);

NAND2xp5_ASAP7_75t_L g7722 ( 
.A(n_6998),
.B(n_5559),
.Y(n_7722)
);

NAND2xp5_ASAP7_75t_L g7723 ( 
.A(n_6998),
.B(n_5526),
.Y(n_7723)
);

AOI21xp5_ASAP7_75t_L g7724 ( 
.A1(n_6401),
.A2(n_5451),
.B(n_5526),
.Y(n_7724)
);

NAND2xp5_ASAP7_75t_L g7725 ( 
.A(n_6999),
.B(n_7188),
.Y(n_7725)
);

OAI22xp5_ASAP7_75t_L g7726 ( 
.A1(n_6748),
.A2(n_6888),
.B1(n_6709),
.B2(n_6693),
.Y(n_7726)
);

HB1xp67_ASAP7_75t_L g7727 ( 
.A(n_7399),
.Y(n_7727)
);

NOR2x1_ASAP7_75t_SL g7728 ( 
.A(n_6327),
.B(n_5451),
.Y(n_7728)
);

HB1xp67_ASAP7_75t_L g7729 ( 
.A(n_7399),
.Y(n_7729)
);

AOI21xp5_ASAP7_75t_L g7730 ( 
.A1(n_6751),
.A2(n_5451),
.B(n_5526),
.Y(n_7730)
);

NAND2xp5_ASAP7_75t_L g7731 ( 
.A(n_6999),
.B(n_5526),
.Y(n_7731)
);

HB1xp67_ASAP7_75t_L g7732 ( 
.A(n_7399),
.Y(n_7732)
);

NAND2xp5_ASAP7_75t_SL g7733 ( 
.A(n_6704),
.B(n_5526),
.Y(n_7733)
);

NAND2xp5_ASAP7_75t_L g7734 ( 
.A(n_7188),
.B(n_7118),
.Y(n_7734)
);

BUFx8_ASAP7_75t_L g7735 ( 
.A(n_6292),
.Y(n_7735)
);

NAND2xp5_ASAP7_75t_L g7736 ( 
.A(n_7118),
.B(n_5526),
.Y(n_7736)
);

AOI21xp5_ASAP7_75t_L g7737 ( 
.A1(n_6751),
.A2(n_5451),
.B(n_5524),
.Y(n_7737)
);

NAND2xp5_ASAP7_75t_L g7738 ( 
.A(n_7131),
.B(n_5524),
.Y(n_7738)
);

AO21x1_ASAP7_75t_L g7739 ( 
.A1(n_6822),
.A2(n_5910),
.B(n_5925),
.Y(n_7739)
);

AOI21xp5_ASAP7_75t_L g7740 ( 
.A1(n_6708),
.A2(n_5451),
.B(n_5524),
.Y(n_7740)
);

A2O1A1Ixp33_ASAP7_75t_L g7741 ( 
.A1(n_6467),
.A2(n_5451),
.B(n_5524),
.C(n_6237),
.Y(n_7741)
);

AOI21xp5_ASAP7_75t_SL g7742 ( 
.A1(n_6745),
.A2(n_6849),
.B(n_6479),
.Y(n_7742)
);

NAND2xp5_ASAP7_75t_L g7743 ( 
.A(n_7131),
.B(n_7138),
.Y(n_7743)
);

OR2x6_ASAP7_75t_L g7744 ( 
.A(n_6602),
.B(n_6623),
.Y(n_7744)
);

NAND2xp5_ASAP7_75t_L g7745 ( 
.A(n_7138),
.B(n_5524),
.Y(n_7745)
);

OAI21x1_ASAP7_75t_L g7746 ( 
.A1(n_6747),
.A2(n_5148),
.B(n_5454),
.Y(n_7746)
);

NOR2xp33_ASAP7_75t_L g7747 ( 
.A(n_6642),
.B(n_6748),
.Y(n_7747)
);

NAND2xp5_ASAP7_75t_SL g7748 ( 
.A(n_6694),
.B(n_5524),
.Y(n_7748)
);

INVx2_ASAP7_75t_SL g7749 ( 
.A(n_7642),
.Y(n_7749)
);

OAI21x1_ASAP7_75t_SL g7750 ( 
.A1(n_7216),
.A2(n_5148),
.B(n_5454),
.Y(n_7750)
);

NOR3xp33_ASAP7_75t_SL g7751 ( 
.A(n_6856),
.B(n_5987),
.C(n_6109),
.Y(n_7751)
);

AND2x4_ASAP7_75t_L g7752 ( 
.A(n_6258),
.B(n_5148),
.Y(n_7752)
);

NOR2x1_ASAP7_75t_SL g7753 ( 
.A(n_6327),
.B(n_5148),
.Y(n_7753)
);

INVx3_ASAP7_75t_L g7754 ( 
.A(n_6854),
.Y(n_7754)
);

NAND2xp5_ASAP7_75t_L g7755 ( 
.A(n_7143),
.B(n_5454),
.Y(n_7755)
);

OA22x2_ASAP7_75t_L g7756 ( 
.A1(n_6479),
.A2(n_5454),
.B1(n_5925),
.B2(n_6109),
.Y(n_7756)
);

OA21x2_ASAP7_75t_L g7757 ( 
.A1(n_6747),
.A2(n_5454),
.B(n_5925),
.Y(n_7757)
);

AOI221xp5_ASAP7_75t_L g7758 ( 
.A1(n_6642),
.A2(n_6741),
.B1(n_6738),
.B2(n_6711),
.C(n_6709),
.Y(n_7758)
);

OAI21x1_ASAP7_75t_L g7759 ( 
.A1(n_6555),
.A2(n_5454),
.B(n_5925),
.Y(n_7759)
);

OAI21x1_ASAP7_75t_L g7760 ( 
.A1(n_6555),
.A2(n_5454),
.B(n_5925),
.Y(n_7760)
);

INVx2_ASAP7_75t_SL g7761 ( 
.A(n_7642),
.Y(n_7761)
);

BUFx6f_ASAP7_75t_L g7762 ( 
.A(n_6578),
.Y(n_7762)
);

AOI21xp5_ASAP7_75t_L g7763 ( 
.A1(n_6708),
.A2(n_5925),
.B(n_6043),
.Y(n_7763)
);

OAI22xp5_ASAP7_75t_L g7764 ( 
.A1(n_6888),
.A2(n_5925),
.B1(n_6223),
.B2(n_6678),
.Y(n_7764)
);

NOR2xp33_ASAP7_75t_L g7765 ( 
.A(n_6856),
.B(n_6223),
.Y(n_7765)
);

OAI21x1_ASAP7_75t_L g7766 ( 
.A1(n_6555),
.A2(n_5925),
.B(n_6223),
.Y(n_7766)
);

NAND2xp5_ASAP7_75t_L g7767 ( 
.A(n_7143),
.B(n_7163),
.Y(n_7767)
);

O2A1O1Ixp33_ASAP7_75t_SL g7768 ( 
.A1(n_6830),
.A2(n_6736),
.B(n_6514),
.C(n_6796),
.Y(n_7768)
);

NAND2xp5_ASAP7_75t_L g7769 ( 
.A(n_7163),
.B(n_7164),
.Y(n_7769)
);

AOI22xp5_ASAP7_75t_L g7770 ( 
.A1(n_6711),
.A2(n_6777),
.B1(n_6785),
.B2(n_6666),
.Y(n_7770)
);

AND2x4_ASAP7_75t_L g7771 ( 
.A(n_6258),
.B(n_6463),
.Y(n_7771)
);

NAND2xp33_ASAP7_75t_R g7772 ( 
.A(n_6928),
.B(n_6301),
.Y(n_7772)
);

A2O1A1Ixp33_ASAP7_75t_L g7773 ( 
.A1(n_6467),
.A2(n_6276),
.B(n_6630),
.C(n_6304),
.Y(n_7773)
);

AND2x2_ASAP7_75t_L g7774 ( 
.A(n_7311),
.B(n_7560),
.Y(n_7774)
);

INVx2_ASAP7_75t_L g7775 ( 
.A(n_7395),
.Y(n_7775)
);

AO21x1_ASAP7_75t_L g7776 ( 
.A1(n_6822),
.A2(n_7100),
.B(n_6873),
.Y(n_7776)
);

A2O1A1Ixp33_ASAP7_75t_L g7777 ( 
.A1(n_6276),
.A2(n_6630),
.B(n_6673),
.C(n_6738),
.Y(n_7777)
);

AOI21xp5_ASAP7_75t_L g7778 ( 
.A1(n_6733),
.A2(n_6739),
.B(n_6737),
.Y(n_7778)
);

INVxp67_ASAP7_75t_SL g7779 ( 
.A(n_6416),
.Y(n_7779)
);

OAI21x1_ASAP7_75t_L g7780 ( 
.A1(n_6555),
.A2(n_6657),
.B(n_6265),
.Y(n_7780)
);

A2O1A1Ixp33_ASAP7_75t_L g7781 ( 
.A1(n_6673),
.A2(n_6741),
.B(n_6777),
.C(n_6678),
.Y(n_7781)
);

BUFx10_ASAP7_75t_L g7782 ( 
.A(n_6301),
.Y(n_7782)
);

NAND2xp5_ASAP7_75t_L g7783 ( 
.A(n_7164),
.B(n_7166),
.Y(n_7783)
);

AND2x2_ASAP7_75t_L g7784 ( 
.A(n_7560),
.B(n_7396),
.Y(n_7784)
);

AND2x4_ASAP7_75t_L g7785 ( 
.A(n_6258),
.B(n_6463),
.Y(n_7785)
);

O2A1O1Ixp33_ASAP7_75t_L g7786 ( 
.A1(n_6796),
.A2(n_6830),
.B(n_6736),
.C(n_6849),
.Y(n_7786)
);

INVx2_ASAP7_75t_L g7787 ( 
.A(n_7395),
.Y(n_7787)
);

OAI21x1_ASAP7_75t_L g7788 ( 
.A1(n_6350),
.A2(n_6437),
.B(n_6359),
.Y(n_7788)
);

OAI21xp5_ASAP7_75t_L g7789 ( 
.A1(n_6479),
.A2(n_6968),
.B(n_6718),
.Y(n_7789)
);

OAI21x1_ASAP7_75t_L g7790 ( 
.A1(n_6350),
.A2(n_6437),
.B(n_6359),
.Y(n_7790)
);

NOR2xp33_ASAP7_75t_SL g7791 ( 
.A(n_7320),
.B(n_6687),
.Y(n_7791)
);

INVx4_ASAP7_75t_L g7792 ( 
.A(n_6480),
.Y(n_7792)
);

AND2x2_ASAP7_75t_L g7793 ( 
.A(n_7560),
.B(n_7396),
.Y(n_7793)
);

OAI21x1_ASAP7_75t_L g7794 ( 
.A1(n_6437),
.A2(n_6625),
.B(n_6578),
.Y(n_7794)
);

O2A1O1Ixp5_ASAP7_75t_L g7795 ( 
.A1(n_7100),
.A2(n_6781),
.B(n_6873),
.C(n_6913),
.Y(n_7795)
);

AOI21xp5_ASAP7_75t_L g7796 ( 
.A1(n_6788),
.A2(n_6792),
.B(n_6896),
.Y(n_7796)
);

NAND3xp33_ASAP7_75t_L g7797 ( 
.A(n_6718),
.B(n_6755),
.C(n_6794),
.Y(n_7797)
);

OR2x6_ASAP7_75t_L g7798 ( 
.A(n_6602),
.B(n_6623),
.Y(n_7798)
);

AO21x1_ASAP7_75t_L g7799 ( 
.A1(n_6913),
.A2(n_7323),
.B(n_7106),
.Y(n_7799)
);

A2O1A1Ixp33_ASAP7_75t_L g7800 ( 
.A1(n_6755),
.A2(n_6694),
.B(n_6908),
.C(n_6896),
.Y(n_7800)
);

OA22x2_ASAP7_75t_L g7801 ( 
.A1(n_7065),
.A2(n_6439),
.B1(n_6620),
.B2(n_6771),
.Y(n_7801)
);

AOI21xp5_ASAP7_75t_L g7802 ( 
.A1(n_6788),
.A2(n_6792),
.B(n_6908),
.Y(n_7802)
);

AOI22xp5_ASAP7_75t_L g7803 ( 
.A1(n_6711),
.A2(n_6785),
.B1(n_6666),
.B2(n_6537),
.Y(n_7803)
);

CKINVDCx5p33_ASAP7_75t_R g7804 ( 
.A(n_7556),
.Y(n_7804)
);

OAI22xp5_ASAP7_75t_L g7805 ( 
.A1(n_6888),
.A2(n_6658),
.B1(n_6984),
.B2(n_6891),
.Y(n_7805)
);

AOI211xp5_ASAP7_75t_L g7806 ( 
.A1(n_6679),
.A2(n_6771),
.B(n_6795),
.C(n_6794),
.Y(n_7806)
);

NAND2xp5_ASAP7_75t_SL g7807 ( 
.A(n_6643),
.B(n_6689),
.Y(n_7807)
);

NOR2x1_ASAP7_75t_R g7808 ( 
.A(n_6581),
.B(n_6641),
.Y(n_7808)
);

OAI21xp33_ASAP7_75t_L g7809 ( 
.A1(n_6968),
.A2(n_6925),
.B(n_6984),
.Y(n_7809)
);

INVx5_ASAP7_75t_L g7810 ( 
.A(n_6602),
.Y(n_7810)
);

OAI22x1_ASAP7_75t_L g7811 ( 
.A1(n_7106),
.A2(n_7065),
.B1(n_6439),
.B2(n_7078),
.Y(n_7811)
);

NAND2xp5_ASAP7_75t_L g7812 ( 
.A(n_7166),
.B(n_7169),
.Y(n_7812)
);

NAND2xp5_ASAP7_75t_L g7813 ( 
.A(n_7169),
.B(n_6450),
.Y(n_7813)
);

INVx2_ASAP7_75t_L g7814 ( 
.A(n_7395),
.Y(n_7814)
);

BUFx3_ASAP7_75t_L g7815 ( 
.A(n_7449),
.Y(n_7815)
);

AOI211x1_ASAP7_75t_L g7816 ( 
.A1(n_6793),
.A2(n_6857),
.B(n_6795),
.C(n_7181),
.Y(n_7816)
);

NOR2x1_ASAP7_75t_SL g7817 ( 
.A(n_6327),
.B(n_6309),
.Y(n_7817)
);

NAND2xp5_ASAP7_75t_L g7818 ( 
.A(n_6450),
.B(n_7161),
.Y(n_7818)
);

AOI21xp5_ASAP7_75t_L g7819 ( 
.A1(n_6695),
.A2(n_6877),
.B(n_6874),
.Y(n_7819)
);

OR2x2_ASAP7_75t_L g7820 ( 
.A(n_6979),
.B(n_7036),
.Y(n_7820)
);

BUFx3_ASAP7_75t_L g7821 ( 
.A(n_7449),
.Y(n_7821)
);

OAI21x1_ASAP7_75t_L g7822 ( 
.A1(n_6625),
.A2(n_6631),
.B(n_6628),
.Y(n_7822)
);

NAND2xp5_ASAP7_75t_L g7823 ( 
.A(n_7161),
.B(n_7165),
.Y(n_7823)
);

OAI21xp5_ASAP7_75t_L g7824 ( 
.A1(n_6958),
.A2(n_6925),
.B(n_6669),
.Y(n_7824)
);

HB1xp67_ASAP7_75t_L g7825 ( 
.A(n_7399),
.Y(n_7825)
);

NAND2xp5_ASAP7_75t_L g7826 ( 
.A(n_7165),
.B(n_7175),
.Y(n_7826)
);

OA22x2_ASAP7_75t_L g7827 ( 
.A1(n_7065),
.A2(n_6439),
.B1(n_6984),
.B2(n_6929),
.Y(n_7827)
);

AOI21xp5_ASAP7_75t_L g7828 ( 
.A1(n_6351),
.A2(n_7048),
.B(n_7094),
.Y(n_7828)
);

NAND2xp5_ASAP7_75t_L g7829 ( 
.A(n_7175),
.B(n_6971),
.Y(n_7829)
);

O2A1O1Ixp5_ASAP7_75t_L g7830 ( 
.A1(n_7168),
.A2(n_6779),
.B(n_7181),
.C(n_6740),
.Y(n_7830)
);

BUFx10_ASAP7_75t_L g7831 ( 
.A(n_6706),
.Y(n_7831)
);

AOI21xp5_ASAP7_75t_L g7832 ( 
.A1(n_7048),
.A2(n_7109),
.B(n_7094),
.Y(n_7832)
);

AOI22xp5_ASAP7_75t_L g7833 ( 
.A1(n_6785),
.A2(n_6537),
.B1(n_6833),
.B2(n_6798),
.Y(n_7833)
);

OR2x2_ASAP7_75t_L g7834 ( 
.A(n_7036),
.B(n_7046),
.Y(n_7834)
);

OAI21x1_ASAP7_75t_L g7835 ( 
.A1(n_6625),
.A2(n_6631),
.B(n_6628),
.Y(n_7835)
);

NAND2xp5_ASAP7_75t_L g7836 ( 
.A(n_6971),
.B(n_6993),
.Y(n_7836)
);

NAND2xp5_ASAP7_75t_L g7837 ( 
.A(n_6993),
.B(n_7218),
.Y(n_7837)
);

AOI21xp5_ASAP7_75t_L g7838 ( 
.A1(n_7109),
.A2(n_7026),
.B(n_7024),
.Y(n_7838)
);

NOR2xp33_ASAP7_75t_SL g7839 ( 
.A(n_7320),
.B(n_6687),
.Y(n_7839)
);

NOR2x1_ASAP7_75t_L g7840 ( 
.A(n_6634),
.B(n_6723),
.Y(n_7840)
);

AOI22xp33_ASAP7_75t_L g7841 ( 
.A1(n_6793),
.A2(n_6883),
.B1(n_6844),
.B2(n_6798),
.Y(n_7841)
);

INVx2_ASAP7_75t_SL g7842 ( 
.A(n_7642),
.Y(n_7842)
);

OAI21xp5_ASAP7_75t_L g7843 ( 
.A1(n_6958),
.A2(n_6669),
.B(n_6779),
.Y(n_7843)
);

AOI21x1_ASAP7_75t_L g7844 ( 
.A1(n_6502),
.A2(n_6685),
.B(n_6647),
.Y(n_7844)
);

AOI21xp5_ASAP7_75t_L g7845 ( 
.A1(n_7024),
.A2(n_7026),
.B(n_6472),
.Y(n_7845)
);

OAI21xp5_ASAP7_75t_L g7846 ( 
.A1(n_6669),
.A2(n_6658),
.B(n_6682),
.Y(n_7846)
);

NOR2xp67_ASAP7_75t_L g7847 ( 
.A(n_7671),
.B(n_7515),
.Y(n_7847)
);

AND2x2_ASAP7_75t_L g7848 ( 
.A(n_7560),
.B(n_7396),
.Y(n_7848)
);

AO31x2_ASAP7_75t_L g7849 ( 
.A1(n_6966),
.A2(n_7134),
.A3(n_7181),
.B(n_7168),
.Y(n_7849)
);

OAI21x1_ASAP7_75t_L g7850 ( 
.A1(n_6628),
.A2(n_6635),
.B(n_6631),
.Y(n_7850)
);

AOI21xp5_ASAP7_75t_L g7851 ( 
.A1(n_6472),
.A2(n_7110),
.B(n_6624),
.Y(n_7851)
);

NAND2xp5_ASAP7_75t_L g7852 ( 
.A(n_7218),
.B(n_7120),
.Y(n_7852)
);

OAI21xp5_ASAP7_75t_L g7853 ( 
.A1(n_6669),
.A2(n_6682),
.B(n_6634),
.Y(n_7853)
);

NAND2xp5_ASAP7_75t_L g7854 ( 
.A(n_7120),
.B(n_6948),
.Y(n_7854)
);

OAI21x1_ASAP7_75t_L g7855 ( 
.A1(n_6631),
.A2(n_6638),
.B(n_6635),
.Y(n_7855)
);

AOI21xp5_ASAP7_75t_L g7856 ( 
.A1(n_7110),
.A2(n_6624),
.B(n_6621),
.Y(n_7856)
);

HB1xp67_ASAP7_75t_L g7857 ( 
.A(n_7399),
.Y(n_7857)
);

OAI21xp33_ASAP7_75t_SL g7858 ( 
.A1(n_7323),
.A2(n_6740),
.B(n_6855),
.Y(n_7858)
);

OAI21x1_ASAP7_75t_L g7859 ( 
.A1(n_6635),
.A2(n_6645),
.B(n_6638),
.Y(n_7859)
);

BUFx6f_ASAP7_75t_L g7860 ( 
.A(n_6635),
.Y(n_7860)
);

INVx5_ASAP7_75t_L g7861 ( 
.A(n_6602),
.Y(n_7861)
);

INVx3_ASAP7_75t_L g7862 ( 
.A(n_6854),
.Y(n_7862)
);

OAI21xp5_ASAP7_75t_L g7863 ( 
.A1(n_6634),
.A2(n_6729),
.B(n_6910),
.Y(n_7863)
);

INVx2_ASAP7_75t_SL g7864 ( 
.A(n_7642),
.Y(n_7864)
);

OAI21xp33_ASAP7_75t_L g7865 ( 
.A1(n_6643),
.A2(n_6689),
.B(n_6910),
.Y(n_7865)
);

AOI22xp5_ASAP7_75t_L g7866 ( 
.A1(n_6833),
.A2(n_6726),
.B1(n_7097),
.B2(n_6857),
.Y(n_7866)
);

NOR2x1_ASAP7_75t_SL g7867 ( 
.A(n_6309),
.B(n_6310),
.Y(n_7867)
);

OAI21x1_ASAP7_75t_L g7868 ( 
.A1(n_6638),
.A2(n_6650),
.B(n_6645),
.Y(n_7868)
);

INVxp67_ASAP7_75t_L g7869 ( 
.A(n_6723),
.Y(n_7869)
);

INVx3_ASAP7_75t_L g7870 ( 
.A(n_6854),
.Y(n_7870)
);

A2O1A1Ixp33_ASAP7_75t_L g7871 ( 
.A1(n_7088),
.A2(n_6753),
.B(n_6855),
.C(n_6663),
.Y(n_7871)
);

OR2x2_ASAP7_75t_L g7872 ( 
.A(n_7036),
.B(n_7046),
.Y(n_7872)
);

AOI21x1_ASAP7_75t_L g7873 ( 
.A1(n_6502),
.A2(n_6685),
.B(n_6647),
.Y(n_7873)
);

NOR2xp33_ASAP7_75t_L g7874 ( 
.A(n_6883),
.B(n_7044),
.Y(n_7874)
);

AO21x2_ASAP7_75t_L g7875 ( 
.A1(n_6665),
.A2(n_6672),
.B(n_6668),
.Y(n_7875)
);

INVx3_ASAP7_75t_L g7876 ( 
.A(n_6866),
.Y(n_7876)
);

OAI21x1_ASAP7_75t_L g7877 ( 
.A1(n_6638),
.A2(n_6650),
.B(n_6645),
.Y(n_7877)
);

OAI21x1_ASAP7_75t_L g7878 ( 
.A1(n_6645),
.A2(n_6651),
.B(n_6650),
.Y(n_7878)
);

NAND2xp5_ASAP7_75t_L g7879 ( 
.A(n_6948),
.B(n_6956),
.Y(n_7879)
);

INVx2_ASAP7_75t_SL g7880 ( 
.A(n_7642),
.Y(n_7880)
);

BUFx2_ASAP7_75t_L g7881 ( 
.A(n_7479),
.Y(n_7881)
);

NOR2xp33_ASAP7_75t_L g7882 ( 
.A(n_7044),
.B(n_6851),
.Y(n_7882)
);

AND2x2_ASAP7_75t_SL g7883 ( 
.A(n_7125),
.B(n_6528),
.Y(n_7883)
);

INVx3_ASAP7_75t_L g7884 ( 
.A(n_6866),
.Y(n_7884)
);

A2O1A1Ixp33_ASAP7_75t_L g7885 ( 
.A1(n_7088),
.A2(n_6753),
.B(n_6663),
.C(n_6990),
.Y(n_7885)
);

BUFx3_ASAP7_75t_L g7886 ( 
.A(n_7449),
.Y(n_7886)
);

AOI21xp5_ASAP7_75t_L g7887 ( 
.A1(n_6674),
.A2(n_6681),
.B(n_6475),
.Y(n_7887)
);

OAI21x1_ASAP7_75t_L g7888 ( 
.A1(n_6651),
.A2(n_6659),
.B(n_6656),
.Y(n_7888)
);

NOR2x1_ASAP7_75t_L g7889 ( 
.A(n_7206),
.B(n_6871),
.Y(n_7889)
);

OAI21x1_ASAP7_75t_L g7890 ( 
.A1(n_6651),
.A2(n_6659),
.B(n_6656),
.Y(n_7890)
);

AOI211x1_ASAP7_75t_L g7891 ( 
.A1(n_7181),
.A2(n_7168),
.B(n_6846),
.C(n_6836),
.Y(n_7891)
);

AND2x2_ASAP7_75t_L g7892 ( 
.A(n_7396),
.B(n_7408),
.Y(n_7892)
);

NAND2xp5_ASAP7_75t_L g7893 ( 
.A(n_6956),
.B(n_7091),
.Y(n_7893)
);

AND2x2_ASAP7_75t_L g7894 ( 
.A(n_7408),
.B(n_7364),
.Y(n_7894)
);

INVx3_ASAP7_75t_L g7895 ( 
.A(n_6866),
.Y(n_7895)
);

OAI21x1_ASAP7_75t_L g7896 ( 
.A1(n_6651),
.A2(n_6659),
.B(n_6656),
.Y(n_7896)
);

NAND2xp5_ASAP7_75t_L g7897 ( 
.A(n_7091),
.B(n_7534),
.Y(n_7897)
);

NAND2xp5_ASAP7_75t_L g7898 ( 
.A(n_7534),
.B(n_7149),
.Y(n_7898)
);

NAND2xp5_ASAP7_75t_L g7899 ( 
.A(n_7534),
.B(n_7149),
.Y(n_7899)
);

OAI21x1_ASAP7_75t_L g7900 ( 
.A1(n_6656),
.A2(n_6662),
.B(n_6659),
.Y(n_7900)
);

INVx5_ASAP7_75t_L g7901 ( 
.A(n_6602),
.Y(n_7901)
);

OAI22x1_ASAP7_75t_L g7902 ( 
.A1(n_7065),
.A2(n_6439),
.B1(n_7078),
.B2(n_7039),
.Y(n_7902)
);

INVx3_ASAP7_75t_L g7903 ( 
.A(n_6866),
.Y(n_7903)
);

INVx4_ASAP7_75t_L g7904 ( 
.A(n_6480),
.Y(n_7904)
);

OAI21x1_ASAP7_75t_L g7905 ( 
.A1(n_6662),
.A2(n_6698),
.B(n_6717),
.Y(n_7905)
);

OAI21x1_ASAP7_75t_L g7906 ( 
.A1(n_6662),
.A2(n_6698),
.B(n_6717),
.Y(n_7906)
);

AOI21x1_ASAP7_75t_SL g7907 ( 
.A1(n_7139),
.A2(n_6534),
.B(n_6500),
.Y(n_7907)
);

OAI22xp5_ASAP7_75t_L g7908 ( 
.A1(n_6891),
.A2(n_6851),
.B1(n_6729),
.B2(n_6726),
.Y(n_7908)
);

AOI22xp5_ASAP7_75t_L g7909 ( 
.A1(n_6726),
.A2(n_7097),
.B1(n_6804),
.B2(n_6962),
.Y(n_7909)
);

AOI21xp5_ASAP7_75t_L g7910 ( 
.A1(n_6911),
.A2(n_6912),
.B(n_7111),
.Y(n_7910)
);

O2A1O1Ixp33_ASAP7_75t_SL g7911 ( 
.A1(n_6514),
.A2(n_7249),
.B(n_6362),
.C(n_6360),
.Y(n_7911)
);

BUFx2_ASAP7_75t_L g7912 ( 
.A(n_7479),
.Y(n_7912)
);

AOI21x1_ASAP7_75t_L g7913 ( 
.A1(n_6647),
.A2(n_6575),
.B(n_6329),
.Y(n_7913)
);

AOI21xp5_ASAP7_75t_L g7914 ( 
.A1(n_7111),
.A2(n_6257),
.B(n_6670),
.Y(n_7914)
);

AND2x4_ASAP7_75t_L g7915 ( 
.A(n_6258),
.B(n_6463),
.Y(n_7915)
);

NAND2xp5_ASAP7_75t_L g7916 ( 
.A(n_7157),
.B(n_6917),
.Y(n_7916)
);

NAND2xp5_ASAP7_75t_L g7917 ( 
.A(n_7157),
.B(n_6917),
.Y(n_7917)
);

INVxp67_ASAP7_75t_SL g7918 ( 
.A(n_6416),
.Y(n_7918)
);

AOI21xp5_ASAP7_75t_L g7919 ( 
.A1(n_6257),
.A2(n_6670),
.B(n_6654),
.Y(n_7919)
);

AOI21xp5_ASAP7_75t_L g7920 ( 
.A1(n_6670),
.A2(n_6654),
.B(n_6632),
.Y(n_7920)
);

NOR2xp67_ASAP7_75t_L g7921 ( 
.A(n_7671),
.B(n_7515),
.Y(n_7921)
);

NAND2xp5_ASAP7_75t_L g7922 ( 
.A(n_6917),
.B(n_6534),
.Y(n_7922)
);

NOR2xp33_ASAP7_75t_L g7923 ( 
.A(n_7057),
.B(n_7236),
.Y(n_7923)
);

NAND2xp5_ASAP7_75t_SL g7924 ( 
.A(n_6962),
.B(n_6894),
.Y(n_7924)
);

AOI21xp5_ASAP7_75t_L g7925 ( 
.A1(n_6670),
.A2(n_6632),
.B(n_6800),
.Y(n_7925)
);

OAI21x1_ASAP7_75t_L g7926 ( 
.A1(n_6791),
.A2(n_6797),
.B(n_6705),
.Y(n_7926)
);

AO21x1_ASAP7_75t_L g7927 ( 
.A1(n_7189),
.A2(n_7057),
.B(n_7248),
.Y(n_7927)
);

OAI21xp5_ASAP7_75t_L g7928 ( 
.A1(n_6655),
.A2(n_7098),
.B(n_7005),
.Y(n_7928)
);

BUFx4_ASAP7_75t_SL g7929 ( 
.A(n_7068),
.Y(n_7929)
);

INVx2_ASAP7_75t_SL g7930 ( 
.A(n_7479),
.Y(n_7930)
);

NOR2xp33_ASAP7_75t_L g7931 ( 
.A(n_7236),
.B(n_6949),
.Y(n_7931)
);

OAI21x1_ASAP7_75t_L g7932 ( 
.A1(n_6791),
.A2(n_6797),
.B(n_6705),
.Y(n_7932)
);

OAI21xp5_ASAP7_75t_L g7933 ( 
.A1(n_6655),
.A2(n_7098),
.B(n_7005),
.Y(n_7933)
);

NAND2xp5_ASAP7_75t_SL g7934 ( 
.A(n_6894),
.B(n_6871),
.Y(n_7934)
);

NAND2xp5_ASAP7_75t_L g7935 ( 
.A(n_7639),
.B(n_7648),
.Y(n_7935)
);

OAI21x1_ASAP7_75t_L g7936 ( 
.A1(n_6797),
.A2(n_6705),
.B(n_6774),
.Y(n_7936)
);

A2O1A1Ixp33_ASAP7_75t_L g7937 ( 
.A1(n_6886),
.A2(n_6675),
.B(n_7249),
.C(n_7040),
.Y(n_7937)
);

OAI21x1_ASAP7_75t_L g7938 ( 
.A1(n_6797),
.A2(n_6705),
.B(n_6774),
.Y(n_7938)
);

OAI21x1_ASAP7_75t_L g7939 ( 
.A1(n_6774),
.A2(n_6754),
.B(n_6749),
.Y(n_7939)
);

OAI21x1_ASAP7_75t_L g7940 ( 
.A1(n_6749),
.A2(n_6758),
.B(n_6754),
.Y(n_7940)
);

OAI21x1_ASAP7_75t_SL g7941 ( 
.A1(n_7225),
.A2(n_7241),
.B(n_7134),
.Y(n_7941)
);

NAND2xp5_ASAP7_75t_L g7942 ( 
.A(n_7639),
.B(n_7648),
.Y(n_7942)
);

NOR2xp33_ASAP7_75t_SL g7943 ( 
.A(n_7320),
.B(n_7190),
.Y(n_7943)
);

NAND3xp33_ASAP7_75t_L g7944 ( 
.A(n_6844),
.B(n_6886),
.C(n_6804),
.Y(n_7944)
);

OAI21x1_ASAP7_75t_L g7945 ( 
.A1(n_6749),
.A2(n_6758),
.B(n_6754),
.Y(n_7945)
);

OAI21x1_ASAP7_75t_L g7946 ( 
.A1(n_6749),
.A2(n_6758),
.B(n_6754),
.Y(n_7946)
);

AO21x1_ASAP7_75t_L g7947 ( 
.A1(n_7189),
.A2(n_7248),
.B(n_6881),
.Y(n_7947)
);

AND2x2_ASAP7_75t_L g7948 ( 
.A(n_7408),
.B(n_7364),
.Y(n_7948)
);

AND2x2_ASAP7_75t_L g7949 ( 
.A(n_7408),
.B(n_7364),
.Y(n_7949)
);

OAI21xp5_ASAP7_75t_L g7950 ( 
.A1(n_6655),
.A2(n_6787),
.B(n_6982),
.Y(n_7950)
);

A2O1A1Ixp33_ASAP7_75t_L g7951 ( 
.A1(n_6675),
.A2(n_7040),
.B(n_6881),
.C(n_7237),
.Y(n_7951)
);

AND2x4_ASAP7_75t_L g7952 ( 
.A(n_6463),
.B(n_6544),
.Y(n_7952)
);

NAND2xp33_ASAP7_75t_R g7953 ( 
.A(n_6928),
.B(n_6842),
.Y(n_7953)
);

AO31x2_ASAP7_75t_L g7954 ( 
.A1(n_6385),
.A2(n_6270),
.A3(n_7250),
.B(n_7193),
.Y(n_7954)
);

NOR4xp25_ASAP7_75t_L g7955 ( 
.A(n_7059),
.B(n_6965),
.C(n_6846),
.D(n_6802),
.Y(n_7955)
);

AOI22xp5_ASAP7_75t_L g7956 ( 
.A1(n_6726),
.A2(n_6804),
.B1(n_6978),
.B2(n_6802),
.Y(n_7956)
);

AO31x2_ASAP7_75t_L g7957 ( 
.A1(n_6385),
.A2(n_6270),
.A3(n_7250),
.B(n_7193),
.Y(n_7957)
);

AOI21xp5_ASAP7_75t_L g7958 ( 
.A1(n_6995),
.A2(n_6267),
.B(n_6770),
.Y(n_7958)
);

OAI22xp5_ASAP7_75t_L g7959 ( 
.A1(n_6726),
.A2(n_6872),
.B1(n_7154),
.B2(n_6605),
.Y(n_7959)
);

NOR2xp67_ASAP7_75t_L g7960 ( 
.A(n_7671),
.B(n_7515),
.Y(n_7960)
);

OAI21xp5_ASAP7_75t_L g7961 ( 
.A1(n_6655),
.A2(n_6787),
.B(n_6982),
.Y(n_7961)
);

CKINVDCx5p33_ASAP7_75t_R g7962 ( 
.A(n_6499),
.Y(n_7962)
);

NAND2xp5_ASAP7_75t_SL g7963 ( 
.A(n_6965),
.B(n_6836),
.Y(n_7963)
);

AOI21xp5_ASAP7_75t_L g7964 ( 
.A1(n_6995),
.A2(n_7117),
.B(n_7123),
.Y(n_7964)
);

NOR2xp33_ASAP7_75t_L g7965 ( 
.A(n_6949),
.B(n_6686),
.Y(n_7965)
);

CKINVDCx11_ASAP7_75t_R g7966 ( 
.A(n_6499),
.Y(n_7966)
);

AOI21xp5_ASAP7_75t_L g7967 ( 
.A1(n_6995),
.A2(n_6268),
.B(n_7014),
.Y(n_7967)
);

A2O1A1Ixp33_ASAP7_75t_L g7968 ( 
.A1(n_7237),
.A2(n_7031),
.B(n_7144),
.C(n_7151),
.Y(n_7968)
);

NOR4xp25_ASAP7_75t_L g7969 ( 
.A(n_7059),
.B(n_6686),
.C(n_7135),
.D(n_6978),
.Y(n_7969)
);

NAND2xp5_ASAP7_75t_L g7970 ( 
.A(n_7037),
.B(n_7050),
.Y(n_7970)
);

BUFx6f_ASAP7_75t_L g7971 ( 
.A(n_6355),
.Y(n_7971)
);

AOI21xp5_ASAP7_75t_L g7972 ( 
.A1(n_7014),
.A2(n_7179),
.B(n_6807),
.Y(n_7972)
);

AOI21xp5_ASAP7_75t_L g7973 ( 
.A1(n_7179),
.A2(n_6807),
.B(n_6801),
.Y(n_7973)
);

CKINVDCx20_ASAP7_75t_R g7974 ( 
.A(n_7068),
.Y(n_7974)
);

AOI21xp5_ASAP7_75t_L g7975 ( 
.A1(n_6801),
.A2(n_6817),
.B(n_6809),
.Y(n_7975)
);

NAND2xp5_ASAP7_75t_L g7976 ( 
.A(n_7037),
.B(n_7050),
.Y(n_7976)
);

NAND2x1_ASAP7_75t_L g7977 ( 
.A(n_7076),
.B(n_6732),
.Y(n_7977)
);

OAI21xp5_ASAP7_75t_L g7978 ( 
.A1(n_7031),
.A2(n_7151),
.B(n_7144),
.Y(n_7978)
);

OAI21x1_ASAP7_75t_L g7979 ( 
.A1(n_6764),
.A2(n_6782),
.B(n_6773),
.Y(n_7979)
);

NAND2xp5_ASAP7_75t_L g7980 ( 
.A(n_7060),
.B(n_7064),
.Y(n_7980)
);

NAND2xp5_ASAP7_75t_L g7981 ( 
.A(n_7060),
.B(n_7064),
.Y(n_7981)
);

AOI221xp5_ASAP7_75t_L g7982 ( 
.A1(n_6872),
.A2(n_6939),
.B1(n_7178),
.B2(n_7135),
.C(n_7197),
.Y(n_7982)
);

OAI22xp5_ASAP7_75t_L g7983 ( 
.A1(n_6872),
.A2(n_7154),
.B1(n_6605),
.B2(n_6766),
.Y(n_7983)
);

AOI31xp67_ASAP7_75t_L g7984 ( 
.A1(n_6320),
.A2(n_6322),
.A3(n_6348),
.B(n_6337),
.Y(n_7984)
);

OAI21xp5_ASAP7_75t_L g7985 ( 
.A1(n_7141),
.A2(n_6889),
.B(n_6805),
.Y(n_7985)
);

AO31x2_ASAP7_75t_L g7986 ( 
.A1(n_6270),
.A2(n_7193),
.A3(n_7250),
.B(n_7562),
.Y(n_7986)
);

A2O1A1Ixp33_ASAP7_75t_L g7987 ( 
.A1(n_7328),
.A2(n_6766),
.B(n_6820),
.C(n_7141),
.Y(n_7987)
);

OAI21xp5_ASAP7_75t_L g7988 ( 
.A1(n_6889),
.A2(n_6805),
.B(n_6862),
.Y(n_7988)
);

NOR2xp33_ASAP7_75t_L g7989 ( 
.A(n_7286),
.B(n_6589),
.Y(n_7989)
);

NOR2xp33_ASAP7_75t_L g7990 ( 
.A(n_7286),
.B(n_6589),
.Y(n_7990)
);

A2O1A1Ixp33_ASAP7_75t_L g7991 ( 
.A1(n_7328),
.A2(n_6820),
.B(n_6845),
.C(n_7206),
.Y(n_7991)
);

NAND2xp5_ASAP7_75t_L g7992 ( 
.A(n_7070),
.B(n_7074),
.Y(n_7992)
);

NOR2xp33_ASAP7_75t_L g7993 ( 
.A(n_6614),
.B(n_6619),
.Y(n_7993)
);

NOR2xp33_ASAP7_75t_L g7994 ( 
.A(n_6614),
.B(n_6619),
.Y(n_7994)
);

NAND2xp5_ASAP7_75t_L g7995 ( 
.A(n_7070),
.B(n_7074),
.Y(n_7995)
);

INVx6_ASAP7_75t_L g7996 ( 
.A(n_6952),
.Y(n_7996)
);

HB1xp67_ASAP7_75t_L g7997 ( 
.A(n_7399),
.Y(n_7997)
);

NOR3xp33_ASAP7_75t_L g7998 ( 
.A(n_6286),
.B(n_6939),
.C(n_7450),
.Y(n_7998)
);

NAND2xp5_ASAP7_75t_L g7999 ( 
.A(n_7077),
.B(n_7080),
.Y(n_7999)
);

NAND2xp5_ASAP7_75t_L g8000 ( 
.A(n_7077),
.B(n_7080),
.Y(n_8000)
);

NOR2xp33_ASAP7_75t_L g8001 ( 
.A(n_6636),
.B(n_6649),
.Y(n_8001)
);

NAND3xp33_ASAP7_75t_L g8002 ( 
.A(n_6845),
.B(n_7206),
.C(n_7178),
.Y(n_8002)
);

OAI21x1_ASAP7_75t_L g8003 ( 
.A1(n_6790),
.A2(n_6697),
.B(n_7079),
.Y(n_8003)
);

AOI21xp5_ASAP7_75t_L g8004 ( 
.A1(n_6809),
.A2(n_6818),
.B(n_6817),
.Y(n_8004)
);

AOI21xp5_ASAP7_75t_L g8005 ( 
.A1(n_6818),
.A2(n_6821),
.B(n_6543),
.Y(n_8005)
);

OAI21xp5_ASAP7_75t_L g8006 ( 
.A1(n_6862),
.A2(n_6981),
.B(n_6991),
.Y(n_8006)
);

INVx2_ASAP7_75t_SL g8007 ( 
.A(n_7479),
.Y(n_8007)
);

BUFx2_ASAP7_75t_L g8008 ( 
.A(n_7479),
.Y(n_8008)
);

INVx3_ASAP7_75t_L g8009 ( 
.A(n_6870),
.Y(n_8009)
);

OAI21x1_ASAP7_75t_L g8010 ( 
.A1(n_6697),
.A2(n_7081),
.B(n_7079),
.Y(n_8010)
);

NAND2xp5_ASAP7_75t_SL g8011 ( 
.A(n_7122),
.B(n_7256),
.Y(n_8011)
);

AOI22xp5_ASAP7_75t_L g8012 ( 
.A1(n_7191),
.A2(n_7276),
.B1(n_6862),
.B2(n_7207),
.Y(n_8012)
);

NAND3x1_ASAP7_75t_L g8013 ( 
.A(n_6392),
.B(n_7171),
.C(n_7267),
.Y(n_8013)
);

AOI21xp5_ASAP7_75t_L g8014 ( 
.A1(n_6821),
.A2(n_6543),
.B(n_6945),
.Y(n_8014)
);

INVxp67_ASAP7_75t_L g8015 ( 
.A(n_7371),
.Y(n_8015)
);

AOI21xp33_ASAP7_75t_L g8016 ( 
.A1(n_6861),
.A2(n_7139),
.B(n_7191),
.Y(n_8016)
);

NAND3xp33_ASAP7_75t_SL g8017 ( 
.A(n_6616),
.B(n_7256),
.C(n_7267),
.Y(n_8017)
);

NOR2x1_ASAP7_75t_SL g8018 ( 
.A(n_6309),
.B(n_6310),
.Y(n_8018)
);

AND2x2_ASAP7_75t_L g8019 ( 
.A(n_7124),
.B(n_7150),
.Y(n_8019)
);

INVx4_ASAP7_75t_L g8020 ( 
.A(n_6453),
.Y(n_8020)
);

OR2x6_ASAP7_75t_L g8021 ( 
.A(n_6623),
.B(n_7183),
.Y(n_8021)
);

BUFx12f_ASAP7_75t_L g8022 ( 
.A(n_6595),
.Y(n_8022)
);

A2O1A1Ixp33_ASAP7_75t_L g8023 ( 
.A1(n_6289),
.A2(n_6559),
.B(n_6588),
.C(n_7122),
.Y(n_8023)
);

O2A1O1Ixp33_ASAP7_75t_SL g8024 ( 
.A1(n_6360),
.A2(n_6362),
.B(n_6470),
.C(n_6454),
.Y(n_8024)
);

BUFx12f_ASAP7_75t_L g8025 ( 
.A(n_6595),
.Y(n_8025)
);

NAND2xp5_ASAP7_75t_L g8026 ( 
.A(n_7085),
.B(n_7086),
.Y(n_8026)
);

NOR2xp67_ASAP7_75t_L g8027 ( 
.A(n_7671),
.B(n_7515),
.Y(n_8027)
);

OAI21xp5_ASAP7_75t_L g8028 ( 
.A1(n_6862),
.A2(n_6286),
.B(n_6598),
.Y(n_8028)
);

AOI21xp5_ASAP7_75t_SL g8029 ( 
.A1(n_6390),
.A2(n_6470),
.B(n_6454),
.Y(n_8029)
);

OAI21x1_ASAP7_75t_L g8030 ( 
.A1(n_6697),
.A2(n_7081),
.B(n_7079),
.Y(n_8030)
);

A2O1A1Ixp33_ASAP7_75t_L g8031 ( 
.A1(n_6289),
.A2(n_6559),
.B(n_6588),
.C(n_6812),
.Y(n_8031)
);

OAI21x1_ASAP7_75t_SL g8032 ( 
.A1(n_7225),
.A2(n_7241),
.B(n_7055),
.Y(n_8032)
);

OAI21x1_ASAP7_75t_L g8033 ( 
.A1(n_7079),
.A2(n_7081),
.B(n_6710),
.Y(n_8033)
);

NAND2x1p5_ASAP7_75t_L g8034 ( 
.A(n_7020),
.B(n_7308),
.Y(n_8034)
);

AND2x2_ASAP7_75t_SL g8035 ( 
.A(n_7125),
.B(n_6528),
.Y(n_8035)
);

NAND2xp5_ASAP7_75t_L g8036 ( 
.A(n_7085),
.B(n_7086),
.Y(n_8036)
);

INVx6_ASAP7_75t_L g8037 ( 
.A(n_6952),
.Y(n_8037)
);

AND2x4_ASAP7_75t_L g8038 ( 
.A(n_6463),
.B(n_6544),
.Y(n_8038)
);

NAND2xp5_ASAP7_75t_L g8039 ( 
.A(n_7089),
.B(n_7101),
.Y(n_8039)
);

A2O1A1Ixp33_ASAP7_75t_L g8040 ( 
.A1(n_6812),
.A2(n_6545),
.B(n_6285),
.C(n_7207),
.Y(n_8040)
);

NOR2x1_ASAP7_75t_SL g8041 ( 
.A(n_6309),
.B(n_6310),
.Y(n_8041)
);

OAI21xp5_ASAP7_75t_L g8042 ( 
.A1(n_6598),
.A2(n_6285),
.B(n_7243),
.Y(n_8042)
);

NAND2xp5_ASAP7_75t_L g8043 ( 
.A(n_7089),
.B(n_7101),
.Y(n_8043)
);

INVx2_ASAP7_75t_SL g8044 ( 
.A(n_7465),
.Y(n_8044)
);

AOI21x1_ASAP7_75t_L g8045 ( 
.A1(n_6575),
.A2(n_6329),
.B(n_6326),
.Y(n_8045)
);

CKINVDCx14_ASAP7_75t_R g8046 ( 
.A(n_7263),
.Y(n_8046)
);

NAND2xp5_ASAP7_75t_SL g8047 ( 
.A(n_7125),
.B(n_7207),
.Y(n_8047)
);

AOI22xp33_ASAP7_75t_L g8048 ( 
.A1(n_6861),
.A2(n_7078),
.B1(n_7450),
.B2(n_7197),
.Y(n_8048)
);

NAND2xp5_ASAP7_75t_L g8049 ( 
.A(n_7113),
.B(n_7119),
.Y(n_8049)
);

NAND2x1p5_ASAP7_75t_L g8050 ( 
.A(n_7020),
.B(n_7308),
.Y(n_8050)
);

NAND2xp5_ASAP7_75t_L g8051 ( 
.A(n_7113),
.B(n_7119),
.Y(n_8051)
);

NAND2xp33_ASAP7_75t_L g8052 ( 
.A(n_6523),
.B(n_6926),
.Y(n_8052)
);

AOI21x1_ASAP7_75t_L g8053 ( 
.A1(n_6575),
.A2(n_6329),
.B(n_6326),
.Y(n_8053)
);

AOI21x1_ASAP7_75t_L g8054 ( 
.A1(n_6326),
.A2(n_6379),
.B(n_6367),
.Y(n_8054)
);

INVxp67_ASAP7_75t_L g8055 ( 
.A(n_7371),
.Y(n_8055)
);

OAI21x1_ASAP7_75t_L g8056 ( 
.A1(n_6710),
.A2(n_6498),
.B(n_6712),
.Y(n_8056)
);

AOI21xp5_ASAP7_75t_L g8057 ( 
.A1(n_6521),
.A2(n_6553),
.B(n_7083),
.Y(n_8057)
);

OAI22x1_ASAP7_75t_L g8058 ( 
.A1(n_6929),
.A2(n_7039),
.B1(n_6266),
.B2(n_6464),
.Y(n_8058)
);

BUFx12f_ASAP7_75t_L g8059 ( 
.A(n_7263),
.Y(n_8059)
);

OAI21x1_ASAP7_75t_L g8060 ( 
.A1(n_6498),
.A2(n_6712),
.B(n_6810),
.Y(n_8060)
);

A2O1A1Ixp33_ASAP7_75t_L g8061 ( 
.A1(n_6812),
.A2(n_6545),
.B(n_6417),
.C(n_6501),
.Y(n_8061)
);

NAND2xp5_ASAP7_75t_L g8062 ( 
.A(n_7258),
.B(n_7195),
.Y(n_8062)
);

AND2x4_ASAP7_75t_L g8063 ( 
.A(n_6463),
.B(n_6544),
.Y(n_8063)
);

AO21x1_ASAP7_75t_L g8064 ( 
.A1(n_7243),
.A2(n_7192),
.B(n_7180),
.Y(n_8064)
);

AOI21xp5_ASAP7_75t_L g8065 ( 
.A1(n_6521),
.A2(n_6553),
.B(n_7083),
.Y(n_8065)
);

OAI21x1_ASAP7_75t_L g8066 ( 
.A1(n_6712),
.A2(n_6810),
.B(n_6875),
.Y(n_8066)
);

NOR2x1_ASAP7_75t_L g8067 ( 
.A(n_6392),
.B(n_6330),
.Y(n_8067)
);

NAND2xp5_ASAP7_75t_L g8068 ( 
.A(n_7258),
.B(n_7195),
.Y(n_8068)
);

NAND2xp5_ASAP7_75t_SL g8069 ( 
.A(n_6926),
.B(n_6936),
.Y(n_8069)
);

BUFx6f_ASAP7_75t_L g8070 ( 
.A(n_6355),
.Y(n_8070)
);

AO22x2_ASAP7_75t_L g8071 ( 
.A1(n_6587),
.A2(n_7260),
.B1(n_7039),
.B2(n_6929),
.Y(n_8071)
);

NAND2xp5_ASAP7_75t_L g8072 ( 
.A(n_7199),
.B(n_6263),
.Y(n_8072)
);

NAND2xp5_ASAP7_75t_L g8073 ( 
.A(n_7199),
.B(n_6263),
.Y(n_8073)
);

AND2x4_ASAP7_75t_L g8074 ( 
.A(n_6544),
.B(n_7667),
.Y(n_8074)
);

AOI21x1_ASAP7_75t_L g8075 ( 
.A1(n_6367),
.A2(n_6393),
.B(n_6379),
.Y(n_8075)
);

NAND3xp33_ASAP7_75t_SL g8076 ( 
.A(n_6616),
.B(n_7276),
.C(n_7039),
.Y(n_8076)
);

OAI21x1_ASAP7_75t_L g8077 ( 
.A1(n_6810),
.A2(n_6875),
.B(n_6858),
.Y(n_8077)
);

CKINVDCx20_ASAP7_75t_R g8078 ( 
.A(n_6269),
.Y(n_8078)
);

AOI21xp5_ASAP7_75t_L g8079 ( 
.A1(n_6967),
.A2(n_6264),
.B(n_6519),
.Y(n_8079)
);

NAND2x1p5_ASAP7_75t_L g8080 ( 
.A(n_7020),
.B(n_7308),
.Y(n_8080)
);

OAI21xp5_ASAP7_75t_L g8081 ( 
.A1(n_7192),
.A2(n_6275),
.B(n_6277),
.Y(n_8081)
);

NOR2xp67_ASAP7_75t_L g8082 ( 
.A(n_7515),
.B(n_7660),
.Y(n_8082)
);

O2A1O1Ixp5_ASAP7_75t_L g8083 ( 
.A1(n_6417),
.A2(n_7224),
.B(n_7260),
.C(n_6813),
.Y(n_8083)
);

OAI21xp5_ASAP7_75t_SL g8084 ( 
.A1(n_7108),
.A2(n_6458),
.B(n_6842),
.Y(n_8084)
);

O2A1O1Ixp5_ASAP7_75t_L g8085 ( 
.A1(n_6417),
.A2(n_7224),
.B(n_6813),
.C(n_6431),
.Y(n_8085)
);

AOI21xp5_ASAP7_75t_L g8086 ( 
.A1(n_6264),
.A2(n_6519),
.B(n_6780),
.Y(n_8086)
);

NAND2xp5_ASAP7_75t_L g8087 ( 
.A(n_7214),
.B(n_7373),
.Y(n_8087)
);

INVx4_ASAP7_75t_L g8088 ( 
.A(n_6453),
.Y(n_8088)
);

OAI21x1_ASAP7_75t_L g8089 ( 
.A1(n_6810),
.A2(n_6875),
.B(n_6858),
.Y(n_8089)
);

INVx3_ASAP7_75t_SL g8090 ( 
.A(n_6935),
.Y(n_8090)
);

NAND2xp5_ASAP7_75t_SL g8091 ( 
.A(n_6926),
.B(n_6936),
.Y(n_8091)
);

A2O1A1Ixp33_ASAP7_75t_L g8092 ( 
.A1(n_6390),
.A2(n_6501),
.B(n_6277),
.C(n_6275),
.Y(n_8092)
);

AND2x2_ASAP7_75t_L g8093 ( 
.A(n_7124),
.B(n_7150),
.Y(n_8093)
);

NAND2xp5_ASAP7_75t_L g8094 ( 
.A(n_7214),
.B(n_7373),
.Y(n_8094)
);

AND2x4_ASAP7_75t_L g8095 ( 
.A(n_6544),
.B(n_7667),
.Y(n_8095)
);

INVx3_ASAP7_75t_L g8096 ( 
.A(n_6870),
.Y(n_8096)
);

OAI21x1_ASAP7_75t_L g8097 ( 
.A1(n_6858),
.A2(n_6853),
.B(n_6933),
.Y(n_8097)
);

BUFx2_ASAP7_75t_L g8098 ( 
.A(n_7465),
.Y(n_8098)
);

OAI21x1_ASAP7_75t_L g8099 ( 
.A1(n_6853),
.A2(n_6933),
.B(n_7004),
.Y(n_8099)
);

NAND2xp5_ASAP7_75t_L g8100 ( 
.A(n_7015),
.B(n_7017),
.Y(n_8100)
);

OAI21x1_ASAP7_75t_L g8101 ( 
.A1(n_6853),
.A2(n_6933),
.B(n_7004),
.Y(n_8101)
);

AOI21xp5_ASAP7_75t_L g8102 ( 
.A1(n_6780),
.A2(n_6569),
.B(n_6562),
.Y(n_8102)
);

INVx5_ASAP7_75t_L g8103 ( 
.A(n_7183),
.Y(n_8103)
);

NAND2xp5_ASAP7_75t_L g8104 ( 
.A(n_7015),
.B(n_7017),
.Y(n_8104)
);

AND2x6_ASAP7_75t_SL g8105 ( 
.A(n_6617),
.B(n_6935),
.Y(n_8105)
);

AOI21xp5_ASAP7_75t_L g8106 ( 
.A1(n_6562),
.A2(n_6572),
.B(n_6569),
.Y(n_8106)
);

OAI21xp5_ASAP7_75t_L g8107 ( 
.A1(n_6879),
.A2(n_7200),
.B(n_7108),
.Y(n_8107)
);

OAI21x1_ASAP7_75t_L g8108 ( 
.A1(n_6853),
.A2(n_6933),
.B(n_7004),
.Y(n_8108)
);

NAND2xp5_ASAP7_75t_L g8109 ( 
.A(n_7548),
.B(n_7577),
.Y(n_8109)
);

AOI21xp5_ASAP7_75t_L g8110 ( 
.A1(n_6572),
.A2(n_6576),
.B(n_6466),
.Y(n_8110)
);

OAI22xp5_ASAP7_75t_L g8111 ( 
.A1(n_7276),
.A2(n_6458),
.B1(n_6528),
.B2(n_6929),
.Y(n_8111)
);

NAND2xp5_ASAP7_75t_L g8112 ( 
.A(n_7548),
.B(n_7010),
.Y(n_8112)
);

AND2x2_ASAP7_75t_L g8113 ( 
.A(n_7162),
.B(n_6300),
.Y(n_8113)
);

NAND3x1_ASAP7_75t_L g8114 ( 
.A(n_6392),
.B(n_7171),
.C(n_6505),
.Y(n_8114)
);

OAI21x1_ASAP7_75t_L g8115 ( 
.A1(n_7006),
.A2(n_6954),
.B(n_6950),
.Y(n_8115)
);

AOI21xp5_ASAP7_75t_L g8116 ( 
.A1(n_6576),
.A2(n_6466),
.B(n_6316),
.Y(n_8116)
);

OAI21x1_ASAP7_75t_L g8117 ( 
.A1(n_7006),
.A2(n_6954),
.B(n_6950),
.Y(n_8117)
);

AOI21xp5_ASAP7_75t_L g8118 ( 
.A1(n_6314),
.A2(n_6323),
.B(n_6316),
.Y(n_8118)
);

AOI21xp5_ASAP7_75t_L g8119 ( 
.A1(n_6314),
.A2(n_6331),
.B(n_6323),
.Y(n_8119)
);

OR2x2_ASAP7_75t_L g8120 ( 
.A(n_7162),
.B(n_6438),
.Y(n_8120)
);

NAND2xp5_ASAP7_75t_SL g8121 ( 
.A(n_6926),
.B(n_6936),
.Y(n_8121)
);

NAND2xp5_ASAP7_75t_L g8122 ( 
.A(n_7548),
.B(n_7010),
.Y(n_8122)
);

OAI21x1_ASAP7_75t_L g8123 ( 
.A1(n_7006),
.A2(n_6954),
.B(n_6950),
.Y(n_8123)
);

BUFx10_ASAP7_75t_L g8124 ( 
.A(n_6706),
.Y(n_8124)
);

NAND2xp33_ASAP7_75t_R g8125 ( 
.A(n_6266),
.B(n_6410),
.Y(n_8125)
);

AOI22xp5_ASAP7_75t_L g8126 ( 
.A1(n_6861),
.A2(n_6336),
.B1(n_7331),
.B2(n_6370),
.Y(n_8126)
);

NAND2xp5_ASAP7_75t_L g8127 ( 
.A(n_7210),
.B(n_7228),
.Y(n_8127)
);

OAI21x1_ASAP7_75t_L g8128 ( 
.A1(n_6950),
.A2(n_6954),
.B(n_6893),
.Y(n_8128)
);

AOI221xp5_ASAP7_75t_SL g8129 ( 
.A1(n_7200),
.A2(n_6861),
.B1(n_6613),
.B2(n_6936),
.C(n_7454),
.Y(n_8129)
);

AOI21xp5_ASAP7_75t_L g8130 ( 
.A1(n_6331),
.A2(n_6975),
.B(n_6361),
.Y(n_8130)
);

NAND2xp33_ASAP7_75t_R g8131 ( 
.A(n_6266),
.B(n_6410),
.Y(n_8131)
);

BUFx3_ASAP7_75t_L g8132 ( 
.A(n_7449),
.Y(n_8132)
);

A2O1A1Ixp33_ASAP7_75t_L g8133 ( 
.A1(n_6583),
.A2(n_7353),
.B(n_6271),
.C(n_6547),
.Y(n_8133)
);

AOI21xp5_ASAP7_75t_L g8134 ( 
.A1(n_6975),
.A2(n_6361),
.B(n_6358),
.Y(n_8134)
);

OAI21xp5_ASAP7_75t_L g8135 ( 
.A1(n_7217),
.A2(n_7235),
.B(n_6308),
.Y(n_8135)
);

NAND2xp5_ASAP7_75t_L g8136 ( 
.A(n_7210),
.B(n_7228),
.Y(n_8136)
);

AOI21xp5_ASAP7_75t_SL g8137 ( 
.A1(n_6315),
.A2(n_7334),
.B(n_6600),
.Y(n_8137)
);

AND2x2_ASAP7_75t_L g8138 ( 
.A(n_7162),
.B(n_6300),
.Y(n_8138)
);

OAI21x1_ASAP7_75t_L g8139 ( 
.A1(n_6885),
.A2(n_6898),
.B(n_6893),
.Y(n_8139)
);

OAI22xp5_ASAP7_75t_L g8140 ( 
.A1(n_6528),
.A2(n_7353),
.B1(n_6636),
.B2(n_6671),
.Y(n_8140)
);

OAI21x1_ASAP7_75t_L g8141 ( 
.A1(n_6885),
.A2(n_6898),
.B(n_6893),
.Y(n_8141)
);

OAI21x1_ASAP7_75t_L g8142 ( 
.A1(n_6885),
.A2(n_6903),
.B(n_6898),
.Y(n_8142)
);

NOR4xp25_ASAP7_75t_L g8143 ( 
.A(n_6421),
.B(n_6441),
.C(n_6613),
.D(n_7331),
.Y(n_8143)
);

OAI21x1_ASAP7_75t_L g8144 ( 
.A1(n_6903),
.A2(n_6931),
.B(n_6824),
.Y(n_8144)
);

NAND2x1p5_ASAP7_75t_L g8145 ( 
.A(n_7020),
.B(n_7308),
.Y(n_8145)
);

INVx3_ASAP7_75t_L g8146 ( 
.A(n_6903),
.Y(n_8146)
);

AOI21xp5_ASAP7_75t_L g8147 ( 
.A1(n_6358),
.A2(n_6280),
.B(n_6279),
.Y(n_8147)
);

AOI21xp5_ASAP7_75t_L g8148 ( 
.A1(n_6279),
.A2(n_6294),
.B(n_6280),
.Y(n_8148)
);

OAI21x1_ASAP7_75t_SL g8149 ( 
.A1(n_6730),
.A2(n_7066),
.B(n_7055),
.Y(n_8149)
);

OAI21x1_ASAP7_75t_L g8150 ( 
.A1(n_6931),
.A2(n_6824),
.B(n_6815),
.Y(n_8150)
);

NOR2xp67_ASAP7_75t_SL g8151 ( 
.A(n_6581),
.B(n_6641),
.Y(n_8151)
);

OAI21xp5_ASAP7_75t_L g8152 ( 
.A1(n_7217),
.A2(n_7235),
.B(n_6308),
.Y(n_8152)
);

AOI211x1_ASAP7_75t_L g8153 ( 
.A1(n_6403),
.A2(n_7082),
.B(n_6380),
.C(n_7130),
.Y(n_8153)
);

CKINVDCx20_ASAP7_75t_R g8154 ( 
.A(n_6269),
.Y(n_8154)
);

AOI21xp5_ASAP7_75t_L g8155 ( 
.A1(n_6294),
.A2(n_6592),
.B(n_6328),
.Y(n_8155)
);

A2O1A1Ixp33_ASAP7_75t_L g8156 ( 
.A1(n_6271),
.A2(n_6546),
.B(n_6548),
.C(n_6547),
.Y(n_8156)
);

OAI22xp5_ASAP7_75t_L g8157 ( 
.A1(n_6528),
.A2(n_6671),
.B1(n_6676),
.B2(n_6649),
.Y(n_8157)
);

BUFx2_ASAP7_75t_L g8158 ( 
.A(n_7465),
.Y(n_8158)
);

BUFx3_ASAP7_75t_L g8159 ( 
.A(n_7449),
.Y(n_8159)
);

A2O1A1Ixp33_ASAP7_75t_L g8160 ( 
.A1(n_6271),
.A2(n_6546),
.B(n_6548),
.C(n_6368),
.Y(n_8160)
);

OAI21x1_ASAP7_75t_L g8161 ( 
.A1(n_6931),
.A2(n_6815),
.B(n_6814),
.Y(n_8161)
);

BUFx12f_ASAP7_75t_L g8162 ( 
.A(n_6859),
.Y(n_8162)
);

O2A1O1Ixp5_ASAP7_75t_L g8163 ( 
.A1(n_6431),
.A2(n_6533),
.B(n_6434),
.C(n_6380),
.Y(n_8163)
);

AOI21xp5_ASAP7_75t_L g8164 ( 
.A1(n_6592),
.A2(n_6328),
.B(n_6319),
.Y(n_8164)
);

BUFx6f_ASAP7_75t_L g8165 ( 
.A(n_6355),
.Y(n_8165)
);

AOI21xp5_ASAP7_75t_L g8166 ( 
.A1(n_6319),
.A2(n_6333),
.B(n_6332),
.Y(n_8166)
);

OAI21xp5_ASAP7_75t_SL g8167 ( 
.A1(n_7331),
.A2(n_6441),
.B(n_6421),
.Y(n_8167)
);

INVx2_ASAP7_75t_SL g8168 ( 
.A(n_7465),
.Y(n_8168)
);

A2O1A1Ixp33_ASAP7_75t_L g8169 ( 
.A1(n_6368),
.A2(n_6370),
.B(n_7334),
.C(n_7283),
.Y(n_8169)
);

NAND2xp5_ASAP7_75t_L g8170 ( 
.A(n_7130),
.B(n_7616),
.Y(n_8170)
);

AO32x2_ASAP7_75t_L g8171 ( 
.A1(n_7090),
.A2(n_7302),
.A3(n_7253),
.B1(n_6587),
.B2(n_7369),
.Y(n_8171)
);

AO21x2_ASAP7_75t_L g8172 ( 
.A1(n_6256),
.A2(n_6282),
.B(n_7187),
.Y(n_8172)
);

NAND2xp5_ASAP7_75t_L g8173 ( 
.A(n_7616),
.B(n_7018),
.Y(n_8173)
);

AOI22xp5_ASAP7_75t_L g8174 ( 
.A1(n_6336),
.A2(n_6342),
.B1(n_6347),
.B2(n_6418),
.Y(n_8174)
);

AOI21xp5_ASAP7_75t_L g8175 ( 
.A1(n_6332),
.A2(n_6333),
.B(n_6425),
.Y(n_8175)
);

NAND2xp5_ASAP7_75t_L g8176 ( 
.A(n_7018),
.B(n_7019),
.Y(n_8176)
);

OR2x2_ASAP7_75t_L g8177 ( 
.A(n_6438),
.B(n_7444),
.Y(n_8177)
);

INVx3_ASAP7_75t_L g8178 ( 
.A(n_7412),
.Y(n_8178)
);

NAND2xp5_ASAP7_75t_L g8179 ( 
.A(n_7019),
.B(n_7025),
.Y(n_8179)
);

AO22x2_ASAP7_75t_L g8180 ( 
.A1(n_7445),
.A2(n_6315),
.B1(n_7041),
.B2(n_7344),
.Y(n_8180)
);

BUFx2_ASAP7_75t_L g8181 ( 
.A(n_7465),
.Y(n_8181)
);

OAI22xp5_ASAP7_75t_L g8182 ( 
.A1(n_6676),
.A2(n_6699),
.B1(n_6720),
.B2(n_6719),
.Y(n_8182)
);

NOR3xp33_ASAP7_75t_SL g8183 ( 
.A(n_6859),
.B(n_7093),
.C(n_7028),
.Y(n_8183)
);

NOR2xp33_ASAP7_75t_L g8184 ( 
.A(n_6699),
.B(n_6719),
.Y(n_8184)
);

AOI21xp5_ASAP7_75t_L g8185 ( 
.A1(n_6425),
.A2(n_6491),
.B(n_6490),
.Y(n_8185)
);

AOI21xp5_ASAP7_75t_L g8186 ( 
.A1(n_6425),
.A2(n_6491),
.B(n_6490),
.Y(n_8186)
);

AOI21xp5_ASAP7_75t_L g8187 ( 
.A1(n_6497),
.A2(n_6503),
.B(n_6378),
.Y(n_8187)
);

AOI21xp5_ASAP7_75t_L g8188 ( 
.A1(n_6497),
.A2(n_6503),
.B(n_6378),
.Y(n_8188)
);

NAND2xp5_ASAP7_75t_L g8189 ( 
.A(n_7025),
.B(n_7032),
.Y(n_8189)
);

NOR2xp33_ASAP7_75t_L g8190 ( 
.A(n_6720),
.B(n_6728),
.Y(n_8190)
);

NOR2xp67_ASAP7_75t_SL g8191 ( 
.A(n_6581),
.B(n_6641),
.Y(n_8191)
);

NAND2xp5_ASAP7_75t_SL g8192 ( 
.A(n_7283),
.B(n_7082),
.Y(n_8192)
);

NOR3xp33_ASAP7_75t_L g8193 ( 
.A(n_6403),
.B(n_6608),
.C(n_7035),
.Y(n_8193)
);

OA22x2_ASAP7_75t_L g8194 ( 
.A1(n_6511),
.A2(n_6488),
.B1(n_6884),
.B2(n_7454),
.Y(n_8194)
);

OAI21x1_ASAP7_75t_L g8195 ( 
.A1(n_6814),
.A2(n_6959),
.B(n_6957),
.Y(n_8195)
);

AOI21xp5_ASAP7_75t_L g8196 ( 
.A1(n_6375),
.A2(n_6386),
.B(n_6381),
.Y(n_8196)
);

NOR2xp33_ASAP7_75t_SL g8197 ( 
.A(n_7190),
.B(n_6581),
.Y(n_8197)
);

OR2x2_ASAP7_75t_L g8198 ( 
.A(n_6438),
.B(n_7444),
.Y(n_8198)
);

NOR2xp33_ASAP7_75t_L g8199 ( 
.A(n_6728),
.B(n_6734),
.Y(n_8199)
);

NOR2xp67_ASAP7_75t_L g8200 ( 
.A(n_7515),
.B(n_7660),
.Y(n_8200)
);

A2O1A1Ixp33_ASAP7_75t_L g8201 ( 
.A1(n_7283),
.A2(n_7244),
.B(n_6561),
.C(n_7330),
.Y(n_8201)
);

INVx2_ASAP7_75t_SL g8202 ( 
.A(n_7515),
.Y(n_8202)
);

BUFx10_ASAP7_75t_L g8203 ( 
.A(n_6292),
.Y(n_8203)
);

OAI21x1_ASAP7_75t_L g8204 ( 
.A1(n_6957),
.A2(n_6961),
.B(n_6959),
.Y(n_8204)
);

OAI21x1_ASAP7_75t_L g8205 ( 
.A1(n_6959),
.A2(n_6974),
.B(n_6961),
.Y(n_8205)
);

BUFx10_ASAP7_75t_L g8206 ( 
.A(n_6292),
.Y(n_8206)
);

AND2x4_ASAP7_75t_L g8207 ( 
.A(n_6544),
.B(n_7667),
.Y(n_8207)
);

BUFx6f_ASAP7_75t_L g8208 ( 
.A(n_6355),
.Y(n_8208)
);

BUFx3_ASAP7_75t_L g8209 ( 
.A(n_7449),
.Y(n_8209)
);

NAND2xp33_ASAP7_75t_L g8210 ( 
.A(n_6523),
.B(n_6283),
.Y(n_8210)
);

OAI21x1_ASAP7_75t_L g8211 ( 
.A1(n_6959),
.A2(n_6974),
.B(n_6961),
.Y(n_8211)
);

INVx2_ASAP7_75t_SL g8212 ( 
.A(n_7515),
.Y(n_8212)
);

NOR2xp33_ASAP7_75t_R g8213 ( 
.A(n_6283),
.B(n_7128),
.Y(n_8213)
);

NAND2xp5_ASAP7_75t_L g8214 ( 
.A(n_6743),
.B(n_6757),
.Y(n_8214)
);

NAND2xp5_ASAP7_75t_L g8215 ( 
.A(n_6743),
.B(n_6757),
.Y(n_8215)
);

O2A1O1Ixp33_ASAP7_75t_SL g8216 ( 
.A1(n_7456),
.A2(n_7613),
.B(n_7128),
.C(n_6603),
.Y(n_8216)
);

NAND2xp5_ASAP7_75t_SL g8217 ( 
.A(n_7303),
.B(n_7307),
.Y(n_8217)
);

NAND2xp5_ASAP7_75t_L g8218 ( 
.A(n_6761),
.B(n_6763),
.Y(n_8218)
);

AOI22xp5_ASAP7_75t_L g8219 ( 
.A1(n_6342),
.A2(n_6347),
.B1(n_6418),
.B2(n_6349),
.Y(n_8219)
);

NAND2xp5_ASAP7_75t_L g8220 ( 
.A(n_6761),
.B(n_6763),
.Y(n_8220)
);

AOI21xp5_ASAP7_75t_L g8221 ( 
.A1(n_6375),
.A2(n_6386),
.B(n_6381),
.Y(n_8221)
);

CKINVDCx5p33_ASAP7_75t_R g8222 ( 
.A(n_6577),
.Y(n_8222)
);

AO21x2_ASAP7_75t_L g8223 ( 
.A1(n_6256),
.A2(n_6282),
.B(n_7187),
.Y(n_8223)
);

AOI22xp5_ASAP7_75t_L g8224 ( 
.A1(n_6349),
.A2(n_7280),
.B1(n_6524),
.B2(n_6487),
.Y(n_8224)
);

NAND2xp33_ASAP7_75t_L g8225 ( 
.A(n_6532),
.B(n_6612),
.Y(n_8225)
);

OAI21x1_ASAP7_75t_L g8226 ( 
.A1(n_6961),
.A2(n_6976),
.B(n_6974),
.Y(n_8226)
);

AOI21x1_ASAP7_75t_L g8227 ( 
.A1(n_6367),
.A2(n_6393),
.B(n_6379),
.Y(n_8227)
);

NAND2xp5_ASAP7_75t_SL g8228 ( 
.A(n_7303),
.B(n_7307),
.Y(n_8228)
);

OAI22x1_ASAP7_75t_L g8229 ( 
.A1(n_6410),
.A2(n_6680),
.B1(n_6806),
.B2(n_6464),
.Y(n_8229)
);

NAND2xp5_ASAP7_75t_L g8230 ( 
.A(n_6768),
.B(n_6803),
.Y(n_8230)
);

NAND2xp5_ASAP7_75t_L g8231 ( 
.A(n_6768),
.B(n_6803),
.Y(n_8231)
);

OAI21x1_ASAP7_75t_L g8232 ( 
.A1(n_6974),
.A2(n_6992),
.B(n_6976),
.Y(n_8232)
);

NAND2xp5_ASAP7_75t_L g8233 ( 
.A(n_6823),
.B(n_6827),
.Y(n_8233)
);

NAND3xp33_ASAP7_75t_L g8234 ( 
.A(n_7244),
.B(n_6819),
.C(n_6374),
.Y(n_8234)
);

OAI21xp5_ASAP7_75t_L g8235 ( 
.A1(n_7035),
.A2(n_7167),
.B(n_6593),
.Y(n_8235)
);

OAI21x1_ASAP7_75t_L g8236 ( 
.A1(n_6976),
.A2(n_7000),
.B(n_6992),
.Y(n_8236)
);

OAI21x1_ASAP7_75t_L g8237 ( 
.A1(n_6976),
.A2(n_7000),
.B(n_6992),
.Y(n_8237)
);

OAI21x1_ASAP7_75t_L g8238 ( 
.A1(n_6992),
.A2(n_7001),
.B(n_7000),
.Y(n_8238)
);

NAND3xp33_ASAP7_75t_SL g8239 ( 
.A(n_7499),
.B(n_7478),
.C(n_6533),
.Y(n_8239)
);

OAI22x1_ASAP7_75t_L g8240 ( 
.A1(n_6464),
.A2(n_6806),
.B1(n_6892),
.B2(n_6680),
.Y(n_8240)
);

NAND2xp5_ASAP7_75t_L g8241 ( 
.A(n_6823),
.B(n_6827),
.Y(n_8241)
);

AO21x2_ASAP7_75t_L g8242 ( 
.A1(n_6290),
.A2(n_6307),
.B(n_6297),
.Y(n_8242)
);

NAND2x1p5_ASAP7_75t_L g8243 ( 
.A(n_7020),
.B(n_7308),
.Y(n_8243)
);

NAND2xp5_ASAP7_75t_L g8244 ( 
.A(n_6834),
.B(n_6841),
.Y(n_8244)
);

AOI21x1_ASAP7_75t_L g8245 ( 
.A1(n_6393),
.A2(n_6422),
.B(n_6404),
.Y(n_8245)
);

AOI21xp5_ASAP7_75t_L g8246 ( 
.A1(n_6550),
.A2(n_6944),
.B(n_6918),
.Y(n_8246)
);

AOI21xp5_ASAP7_75t_L g8247 ( 
.A1(n_6550),
.A2(n_6944),
.B(n_6918),
.Y(n_8247)
);

BUFx6f_ASAP7_75t_L g8248 ( 
.A(n_7043),
.Y(n_8248)
);

OAI21x1_ASAP7_75t_L g8249 ( 
.A1(n_7000),
.A2(n_7002),
.B(n_7001),
.Y(n_8249)
);

AND2x4_ASAP7_75t_L g8250 ( 
.A(n_6730),
.B(n_7055),
.Y(n_8250)
);

CKINVDCx20_ASAP7_75t_R g8251 ( 
.A(n_7613),
.Y(n_8251)
);

AOI21x1_ASAP7_75t_L g8252 ( 
.A1(n_6404),
.A2(n_6444),
.B(n_6422),
.Y(n_8252)
);

AND2x2_ASAP7_75t_L g8253 ( 
.A(n_6300),
.B(n_6509),
.Y(n_8253)
);

CKINVDCx20_ASAP7_75t_R g8254 ( 
.A(n_6648),
.Y(n_8254)
);

AOI221x1_ASAP7_75t_L g8255 ( 
.A1(n_6760),
.A2(n_6600),
.B1(n_6518),
.B2(n_6819),
.C(n_6593),
.Y(n_8255)
);

OAI21xp5_ASAP7_75t_L g8256 ( 
.A1(n_7167),
.A2(n_6449),
.B(n_6374),
.Y(n_8256)
);

NAND2x1p5_ASAP7_75t_L g8257 ( 
.A(n_7020),
.B(n_7308),
.Y(n_8257)
);

OAI22xp5_ASAP7_75t_L g8258 ( 
.A1(n_6834),
.A2(n_6841),
.B1(n_6869),
.B2(n_6863),
.Y(n_8258)
);

OAI21xp5_ASAP7_75t_L g8259 ( 
.A1(n_6449),
.A2(n_7330),
.B(n_6443),
.Y(n_8259)
);

O2A1O1Ixp33_ASAP7_75t_SL g8260 ( 
.A1(n_7456),
.A2(n_6603),
.B(n_6539),
.C(n_7488),
.Y(n_8260)
);

NAND2xp5_ASAP7_75t_L g8261 ( 
.A(n_6863),
.B(n_6869),
.Y(n_8261)
);

AOI21xp5_ASAP7_75t_L g8262 ( 
.A1(n_6915),
.A2(n_6932),
.B(n_6922),
.Y(n_8262)
);

NAND3xp33_ASAP7_75t_SL g8263 ( 
.A(n_7499),
.B(n_7478),
.C(n_6533),
.Y(n_8263)
);

OAI21xp5_ASAP7_75t_L g8264 ( 
.A1(n_6427),
.A2(n_6443),
.B(n_6608),
.Y(n_8264)
);

AOI21xp5_ASAP7_75t_L g8265 ( 
.A1(n_6915),
.A2(n_6932),
.B(n_6922),
.Y(n_8265)
);

NOR4xp25_ASAP7_75t_L g8266 ( 
.A(n_7269),
.B(n_6515),
.C(n_7368),
.D(n_7344),
.Y(n_8266)
);

NAND3x1_ASAP7_75t_L g8267 ( 
.A(n_7171),
.B(n_6505),
.C(n_6494),
.Y(n_8267)
);

OAI21x1_ASAP7_75t_L g8268 ( 
.A1(n_7001),
.A2(n_7003),
.B(n_7002),
.Y(n_8268)
);

AO21x2_ASAP7_75t_L g8269 ( 
.A1(n_6290),
.A2(n_6307),
.B(n_6297),
.Y(n_8269)
);

NAND2xp5_ASAP7_75t_L g8270 ( 
.A(n_6876),
.B(n_6878),
.Y(n_8270)
);

OAI21xp5_ASAP7_75t_L g8271 ( 
.A1(n_6427),
.A2(n_7426),
.B(n_6539),
.Y(n_8271)
);

OAI21x1_ASAP7_75t_L g8272 ( 
.A1(n_7001),
.A2(n_7003),
.B(n_7002),
.Y(n_8272)
);

BUFx6f_ASAP7_75t_L g8273 ( 
.A(n_7043),
.Y(n_8273)
);

INVx3_ASAP7_75t_L g8274 ( 
.A(n_7412),
.Y(n_8274)
);

OAI21x1_ASAP7_75t_L g8275 ( 
.A1(n_7002),
.A2(n_7007),
.B(n_7003),
.Y(n_8275)
);

AOI21xp5_ASAP7_75t_L g8276 ( 
.A1(n_6940),
.A2(n_7013),
.B(n_7007),
.Y(n_8276)
);

INVxp67_ASAP7_75t_L g8277 ( 
.A(n_7371),
.Y(n_8277)
);

AOI21xp5_ASAP7_75t_L g8278 ( 
.A1(n_6940),
.A2(n_7013),
.B(n_7007),
.Y(n_8278)
);

AND2x4_ASAP7_75t_L g8279 ( 
.A(n_6730),
.B(n_7066),
.Y(n_8279)
);

AOI21x1_ASAP7_75t_L g8280 ( 
.A1(n_6404),
.A2(n_6444),
.B(n_6422),
.Y(n_8280)
);

AOI21xp5_ASAP7_75t_SL g8281 ( 
.A1(n_6600),
.A2(n_6518),
.B(n_7254),
.Y(n_8281)
);

BUFx12f_ASAP7_75t_L g8282 ( 
.A(n_7028),
.Y(n_8282)
);

AOI21xp5_ASAP7_75t_L g8283 ( 
.A1(n_7003),
.A2(n_7008),
.B(n_7007),
.Y(n_8283)
);

INVx2_ASAP7_75t_SL g8284 ( 
.A(n_7515),
.Y(n_8284)
);

OAI21x1_ASAP7_75t_SL g8285 ( 
.A1(n_7066),
.A2(n_6273),
.B(n_6561),
.Y(n_8285)
);

AND2x2_ASAP7_75t_L g8286 ( 
.A(n_6300),
.B(n_6509),
.Y(n_8286)
);

AO31x2_ASAP7_75t_L g8287 ( 
.A1(n_7608),
.A2(n_6526),
.A3(n_6542),
.B(n_6529),
.Y(n_8287)
);

AOI21xp5_ASAP7_75t_L g8288 ( 
.A1(n_7008),
.A2(n_7021),
.B(n_6601),
.Y(n_8288)
);

AOI221x1_ASAP7_75t_L g8289 ( 
.A1(n_6760),
.A2(n_6600),
.B1(n_6835),
.B2(n_6506),
.C(n_6389),
.Y(n_8289)
);

OAI21xp5_ASAP7_75t_L g8290 ( 
.A1(n_7426),
.A2(n_7343),
.B(n_6394),
.Y(n_8290)
);

AND2x2_ASAP7_75t_L g8291 ( 
.A(n_6509),
.B(n_6541),
.Y(n_8291)
);

AO32x2_ASAP7_75t_L g8292 ( 
.A1(n_7090),
.A2(n_7302),
.A3(n_7253),
.B1(n_7614),
.B2(n_7369),
.Y(n_8292)
);

O2A1O1Ixp5_ASAP7_75t_L g8293 ( 
.A1(n_6434),
.A2(n_6533),
.B(n_6455),
.C(n_6395),
.Y(n_8293)
);

NAND2xp5_ASAP7_75t_SL g8294 ( 
.A(n_7054),
.B(n_7056),
.Y(n_8294)
);

AOI221xp5_ASAP7_75t_L g8295 ( 
.A1(n_7368),
.A2(n_7336),
.B1(n_6811),
.B2(n_7445),
.C(n_7280),
.Y(n_8295)
);

BUFx6f_ASAP7_75t_L g8296 ( 
.A(n_7043),
.Y(n_8296)
);

NAND2xp5_ASAP7_75t_L g8297 ( 
.A(n_6876),
.B(n_6878),
.Y(n_8297)
);

NOR2x1_ASAP7_75t_R g8298 ( 
.A(n_6641),
.B(n_6829),
.Y(n_8298)
);

INVx3_ASAP7_75t_L g8299 ( 
.A(n_7412),
.Y(n_8299)
);

INVx5_ASAP7_75t_L g8300 ( 
.A(n_7183),
.Y(n_8300)
);

NAND2xp5_ASAP7_75t_L g8301 ( 
.A(n_6880),
.B(n_6890),
.Y(n_8301)
);

NAND2xp5_ASAP7_75t_L g8302 ( 
.A(n_6880),
.B(n_6890),
.Y(n_8302)
);

NAND2xp5_ASAP7_75t_L g8303 ( 
.A(n_6901),
.B(n_6904),
.Y(n_8303)
);

NAND2xp5_ASAP7_75t_L g8304 ( 
.A(n_6901),
.B(n_6904),
.Y(n_8304)
);

CKINVDCx5p33_ASAP7_75t_R g8305 ( 
.A(n_6577),
.Y(n_8305)
);

OR2x2_ASAP7_75t_L g8306 ( 
.A(n_7444),
.B(n_7472),
.Y(n_8306)
);

AO21x2_ASAP7_75t_L g8307 ( 
.A1(n_6290),
.A2(n_6307),
.B(n_6297),
.Y(n_8307)
);

NOR2xp33_ASAP7_75t_L g8308 ( 
.A(n_6907),
.B(n_6943),
.Y(n_8308)
);

NAND2xp5_ASAP7_75t_SL g8309 ( 
.A(n_7054),
.B(n_7056),
.Y(n_8309)
);

A2O1A1Ixp33_ASAP7_75t_L g8310 ( 
.A1(n_6395),
.A2(n_6394),
.B(n_6468),
.C(n_7612),
.Y(n_8310)
);

NAND2xp5_ASAP7_75t_L g8311 ( 
.A(n_6907),
.B(n_6943),
.Y(n_8311)
);

OAI22xp5_ASAP7_75t_L g8312 ( 
.A1(n_6946),
.A2(n_6947),
.B1(n_6987),
.B2(n_6986),
.Y(n_8312)
);

A2O1A1Ixp33_ASAP7_75t_L g8313 ( 
.A1(n_6468),
.A2(n_7612),
.B(n_7336),
.C(n_6402),
.Y(n_8313)
);

BUFx6f_ASAP7_75t_L g8314 ( 
.A(n_7043),
.Y(n_8314)
);

INVx3_ASAP7_75t_L g8315 ( 
.A(n_7412),
.Y(n_8315)
);

AOI21xp5_ASAP7_75t_L g8316 ( 
.A1(n_6596),
.A2(n_6606),
.B(n_6604),
.Y(n_8316)
);

NOR2xp33_ASAP7_75t_L g8317 ( 
.A(n_6946),
.B(n_6947),
.Y(n_8317)
);

NAND2xp5_ASAP7_75t_L g8318 ( 
.A(n_6986),
.B(n_6987),
.Y(n_8318)
);

OAI21xp5_ASAP7_75t_L g8319 ( 
.A1(n_7343),
.A2(n_6951),
.B(n_6524),
.Y(n_8319)
);

AOI21xp5_ASAP7_75t_L g8320 ( 
.A1(n_6604),
.A2(n_6606),
.B(n_7245),
.Y(n_8320)
);

AO21x2_ASAP7_75t_L g8321 ( 
.A1(n_6313),
.A2(n_6445),
.B(n_6444),
.Y(n_8321)
);

INVx2_ASAP7_75t_SL g8322 ( 
.A(n_7515),
.Y(n_8322)
);

AOI22xp33_ASAP7_75t_L g8323 ( 
.A1(n_6478),
.A2(n_6487),
.B1(n_6909),
.B2(n_6829),
.Y(n_8323)
);

AOI21xp5_ASAP7_75t_L g8324 ( 
.A1(n_7245),
.A2(n_7254),
.B(n_6346),
.Y(n_8324)
);

AOI22xp33_ASAP7_75t_L g8325 ( 
.A1(n_6478),
.A2(n_6909),
.B1(n_6829),
.B2(n_6442),
.Y(n_8325)
);

AOI21xp5_ASAP7_75t_L g8326 ( 
.A1(n_6334),
.A2(n_6346),
.B(n_6989),
.Y(n_8326)
);

OAI22xp5_ASAP7_75t_L g8327 ( 
.A1(n_6988),
.A2(n_7009),
.B1(n_6488),
.B2(n_7318),
.Y(n_8327)
);

NOR2x1_ASAP7_75t_L g8328 ( 
.A(n_6330),
.B(n_7591),
.Y(n_8328)
);

AOI21xp5_ASAP7_75t_L g8329 ( 
.A1(n_6334),
.A2(n_6989),
.B(n_6415),
.Y(n_8329)
);

NOR4xp25_ASAP7_75t_L g8330 ( 
.A(n_7269),
.B(n_6506),
.C(n_6423),
.D(n_6428),
.Y(n_8330)
);

NAND2xp5_ASAP7_75t_L g8331 ( 
.A(n_6988),
.B(n_7009),
.Y(n_8331)
);

NOR2xp33_ASAP7_75t_L g8332 ( 
.A(n_7140),
.B(n_7174),
.Y(n_8332)
);

OAI21x1_ASAP7_75t_L g8333 ( 
.A1(n_6839),
.A2(n_6847),
.B(n_7586),
.Y(n_8333)
);

NAND2xp5_ASAP7_75t_L g8334 ( 
.A(n_6462),
.B(n_7481),
.Y(n_8334)
);

OR2x2_ASAP7_75t_L g8335 ( 
.A(n_7472),
.B(n_7561),
.Y(n_8335)
);

NAND2xp5_ASAP7_75t_L g8336 ( 
.A(n_6462),
.B(n_7481),
.Y(n_8336)
);

AOI21xp5_ASAP7_75t_SL g8337 ( 
.A1(n_6571),
.A2(n_6590),
.B(n_6469),
.Y(n_8337)
);

CKINVDCx5p33_ASAP7_75t_R g8338 ( 
.A(n_6532),
.Y(n_8338)
);

AOI22xp5_ASAP7_75t_L g8339 ( 
.A1(n_6349),
.A2(n_6478),
.B1(n_6442),
.B2(n_7288),
.Y(n_8339)
);

NOR2xp67_ASAP7_75t_L g8340 ( 
.A(n_7530),
.B(n_7541),
.Y(n_8340)
);

AOI21x1_ASAP7_75t_L g8341 ( 
.A1(n_6445),
.A2(n_6460),
.B(n_6254),
.Y(n_8341)
);

INVxp67_ASAP7_75t_L g8342 ( 
.A(n_7476),
.Y(n_8342)
);

OAI21x1_ASAP7_75t_L g8343 ( 
.A1(n_6839),
.A2(n_6847),
.B(n_7592),
.Y(n_8343)
);

BUFx4f_ASAP7_75t_L g8344 ( 
.A(n_6531),
.Y(n_8344)
);

OAI21x1_ASAP7_75t_SL g8345 ( 
.A1(n_6273),
.A2(n_7638),
.B(n_6434),
.Y(n_8345)
);

OAI21x1_ASAP7_75t_SL g8346 ( 
.A1(n_6273),
.A2(n_7638),
.B(n_6434),
.Y(n_8346)
);

A2O1A1Ixp33_ASAP7_75t_L g8347 ( 
.A1(n_6468),
.A2(n_6402),
.B(n_7306),
.C(n_6488),
.Y(n_8347)
);

OAI21x1_ASAP7_75t_L g8348 ( 
.A1(n_6839),
.A2(n_7592),
.B(n_6424),
.Y(n_8348)
);

BUFx6f_ASAP7_75t_L g8349 ( 
.A(n_7061),
.Y(n_8349)
);

NAND2xp5_ASAP7_75t_SL g8350 ( 
.A(n_7058),
.B(n_7067),
.Y(n_8350)
);

NAND2xp5_ASAP7_75t_L g8351 ( 
.A(n_7481),
.B(n_7268),
.Y(n_8351)
);

OAI21x1_ASAP7_75t_L g8352 ( 
.A1(n_6424),
.A2(n_7030),
.B(n_7142),
.Y(n_8352)
);

CKINVDCx9p33_ASAP7_75t_R g8353 ( 
.A(n_7288),
.Y(n_8353)
);

NAND2xp5_ASAP7_75t_L g8354 ( 
.A(n_7481),
.B(n_7268),
.Y(n_8354)
);

OAI21x1_ASAP7_75t_L g8355 ( 
.A1(n_7030),
.A2(n_7142),
.B(n_6594),
.Y(n_8355)
);

NAND2xp5_ASAP7_75t_L g8356 ( 
.A(n_7481),
.B(n_7275),
.Y(n_8356)
);

NAND2xp5_ASAP7_75t_L g8357 ( 
.A(n_7481),
.B(n_7275),
.Y(n_8357)
);

AOI21xp5_ASAP7_75t_L g8358 ( 
.A1(n_6989),
.A2(n_6428),
.B(n_6406),
.Y(n_8358)
);

OAI21x1_ASAP7_75t_L g8359 ( 
.A1(n_7030),
.A2(n_6594),
.B(n_7034),
.Y(n_8359)
);

OAI21x1_ASAP7_75t_L g8360 ( 
.A1(n_6594),
.A2(n_7034),
.B(n_7203),
.Y(n_8360)
);

OAI21xp5_ASAP7_75t_SL g8361 ( 
.A1(n_6511),
.A2(n_7434),
.B(n_7329),
.Y(n_8361)
);

NAND2xp5_ASAP7_75t_L g8362 ( 
.A(n_7591),
.B(n_7607),
.Y(n_8362)
);

AND2x2_ASAP7_75t_L g8363 ( 
.A(n_6509),
.B(n_6541),
.Y(n_8363)
);

OAI22x1_ASAP7_75t_L g8364 ( 
.A1(n_6680),
.A2(n_6892),
.B1(n_6806),
.B2(n_7423),
.Y(n_8364)
);

AOI21xp5_ASAP7_75t_L g8365 ( 
.A1(n_6339),
.A2(n_6354),
.B(n_6306),
.Y(n_8365)
);

NAND2xp5_ASAP7_75t_L g8366 ( 
.A(n_7591),
.B(n_7607),
.Y(n_8366)
);

AOI21x1_ASAP7_75t_L g8367 ( 
.A1(n_6445),
.A2(n_6460),
.B(n_6254),
.Y(n_8367)
);

NAND2xp5_ASAP7_75t_SL g8368 ( 
.A(n_7058),
.B(n_7067),
.Y(n_8368)
);

OR2x6_ASAP7_75t_L g8369 ( 
.A(n_6623),
.B(n_7183),
.Y(n_8369)
);

AND2x6_ASAP7_75t_L g8370 ( 
.A(n_6284),
.B(n_6511),
.Y(n_8370)
);

AOI21xp5_ASAP7_75t_L g8371 ( 
.A1(n_6339),
.A2(n_6354),
.B(n_6306),
.Y(n_8371)
);

OAI21x1_ASAP7_75t_L g8372 ( 
.A1(n_7034),
.A2(n_7213),
.B(n_7203),
.Y(n_8372)
);

AOI21xp5_ASAP7_75t_L g8373 ( 
.A1(n_6305),
.A2(n_6318),
.B(n_6311),
.Y(n_8373)
);

INVx3_ASAP7_75t_SL g8374 ( 
.A(n_6291),
.Y(n_8374)
);

OAI21xp5_ASAP7_75t_L g8375 ( 
.A1(n_6951),
.A2(n_6452),
.B(n_6451),
.Y(n_8375)
);

OAI21x1_ASAP7_75t_L g8376 ( 
.A1(n_7034),
.A2(n_7213),
.B(n_6554),
.Y(n_8376)
);

AOI22xp5_ASAP7_75t_L g8377 ( 
.A1(n_6478),
.A2(n_7329),
.B1(n_6513),
.B2(n_6469),
.Y(n_8377)
);

BUFx3_ASAP7_75t_L g8378 ( 
.A(n_7449),
.Y(n_8378)
);

O2A1O1Ixp33_ASAP7_75t_L g8379 ( 
.A1(n_6811),
.A2(n_7174),
.B(n_7140),
.C(n_6389),
.Y(n_8379)
);

OAI21x1_ASAP7_75t_L g8380 ( 
.A1(n_6540),
.A2(n_6554),
.B(n_7061),
.Y(n_8380)
);

AOI21xp5_ASAP7_75t_L g8381 ( 
.A1(n_6305),
.A2(n_6318),
.B(n_6311),
.Y(n_8381)
);

AND2x2_ASAP7_75t_L g8382 ( 
.A(n_6541),
.B(n_6622),
.Y(n_8382)
);

NAND2xp5_ASAP7_75t_L g8383 ( 
.A(n_7607),
.B(n_7636),
.Y(n_8383)
);

AO31x2_ASAP7_75t_L g8384 ( 
.A1(n_6639),
.A2(n_6646),
.A3(n_6653),
.B(n_7559),
.Y(n_8384)
);

AOI21xp5_ASAP7_75t_L g8385 ( 
.A1(n_6363),
.A2(n_6373),
.B(n_6371),
.Y(n_8385)
);

NAND2xp5_ASAP7_75t_L g8386 ( 
.A(n_7636),
.B(n_7558),
.Y(n_8386)
);

NOR2xp67_ASAP7_75t_L g8387 ( 
.A(n_7530),
.B(n_7541),
.Y(n_8387)
);

A2O1A1Ixp33_ASAP7_75t_L g8388 ( 
.A1(n_6402),
.A2(n_7306),
.B(n_6590),
.C(n_6571),
.Y(n_8388)
);

NAND3x1_ASAP7_75t_L g8389 ( 
.A(n_6505),
.B(n_6494),
.C(n_7305),
.Y(n_8389)
);

NAND2xp5_ASAP7_75t_L g8390 ( 
.A(n_7636),
.B(n_7558),
.Y(n_8390)
);

OAI21xp5_ASAP7_75t_SL g8391 ( 
.A1(n_7434),
.A2(n_7329),
.B(n_6455),
.Y(n_8391)
);

OAI21x1_ASAP7_75t_L g8392 ( 
.A1(n_6540),
.A2(n_6554),
.B(n_7061),
.Y(n_8392)
);

A2O1A1Ixp33_ASAP7_75t_L g8393 ( 
.A1(n_7596),
.A2(n_7609),
.B(n_7312),
.C(n_7314),
.Y(n_8393)
);

AND2x2_ASAP7_75t_L g8394 ( 
.A(n_6541),
.B(n_6622),
.Y(n_8394)
);

NAND3xp33_ASAP7_75t_L g8395 ( 
.A(n_7341),
.B(n_7407),
.C(n_6369),
.Y(n_8395)
);

AO31x2_ASAP7_75t_L g8396 ( 
.A1(n_6639),
.A2(n_6646),
.A3(n_6653),
.B(n_7559),
.Y(n_8396)
);

AOI21xp5_ASAP7_75t_L g8397 ( 
.A1(n_6363),
.A2(n_6373),
.B(n_6371),
.Y(n_8397)
);

INVx3_ASAP7_75t_L g8398 ( 
.A(n_7238),
.Y(n_8398)
);

AO32x2_ASAP7_75t_L g8399 ( 
.A1(n_7090),
.A2(n_7302),
.A3(n_7253),
.B1(n_7614),
.B2(n_7369),
.Y(n_8399)
);

AOI21xp5_ASAP7_75t_L g8400 ( 
.A1(n_6584),
.A2(n_7568),
.B(n_7563),
.Y(n_8400)
);

BUFx3_ASAP7_75t_L g8401 ( 
.A(n_7449),
.Y(n_8401)
);

OAI21xp5_ASAP7_75t_L g8402 ( 
.A1(n_6451),
.A2(n_6452),
.B(n_7087),
.Y(n_8402)
);

AOI22xp5_ASAP7_75t_L g8403 ( 
.A1(n_6478),
.A2(n_6513),
.B1(n_6469),
.B2(n_6383),
.Y(n_8403)
);

OAI21xp5_ASAP7_75t_L g8404 ( 
.A1(n_7087),
.A2(n_6484),
.B(n_6504),
.Y(n_8404)
);

BUFx6f_ASAP7_75t_L g8405 ( 
.A(n_7183),
.Y(n_8405)
);

OAI21x1_ASAP7_75t_L g8406 ( 
.A1(n_6540),
.A2(n_6435),
.B(n_6261),
.Y(n_8406)
);

OA22x2_ASAP7_75t_L g8407 ( 
.A1(n_6811),
.A2(n_6383),
.B1(n_6321),
.B2(n_7654),
.Y(n_8407)
);

OAI21xp5_ASAP7_75t_L g8408 ( 
.A1(n_6484),
.A2(n_6504),
.B(n_7133),
.Y(n_8408)
);

OAI21x1_ASAP7_75t_L g8409 ( 
.A1(n_6435),
.A2(n_6261),
.B(n_6260),
.Y(n_8409)
);

INVx3_ASAP7_75t_L g8410 ( 
.A(n_7238),
.Y(n_8410)
);

AO31x2_ASAP7_75t_L g8411 ( 
.A1(n_6646),
.A2(n_6653),
.A3(n_7559),
.B(n_6321),
.Y(n_8411)
);

AOI21xp5_ASAP7_75t_L g8412 ( 
.A1(n_7563),
.A2(n_7574),
.B(n_7568),
.Y(n_8412)
);

AOI22xp5_ASAP7_75t_L g8413 ( 
.A1(n_6478),
.A2(n_6513),
.B1(n_6469),
.B2(n_6383),
.Y(n_8413)
);

A2O1A1Ixp33_ASAP7_75t_L g8414 ( 
.A1(n_7596),
.A2(n_7609),
.B(n_7312),
.C(n_7314),
.Y(n_8414)
);

INVx3_ASAP7_75t_L g8415 ( 
.A(n_7238),
.Y(n_8415)
);

CKINVDCx5p33_ASAP7_75t_R g8416 ( 
.A(n_7332),
.Y(n_8416)
);

AOI21xp5_ASAP7_75t_L g8417 ( 
.A1(n_7574),
.A2(n_7576),
.B(n_6409),
.Y(n_8417)
);

NAND3x1_ASAP7_75t_L g8418 ( 
.A(n_6494),
.B(n_7317),
.C(n_7305),
.Y(n_8418)
);

AOI21xp5_ASAP7_75t_L g8419 ( 
.A1(n_7576),
.A2(n_6409),
.B(n_6400),
.Y(n_8419)
);

INVx5_ASAP7_75t_L g8420 ( 
.A(n_7183),
.Y(n_8420)
);

BUFx3_ASAP7_75t_L g8421 ( 
.A(n_7449),
.Y(n_8421)
);

OAI21x1_ASAP7_75t_L g8422 ( 
.A1(n_6260),
.A2(n_6261),
.B(n_7069),
.Y(n_8422)
);

NOR2xp33_ASAP7_75t_L g8423 ( 
.A(n_7403),
.B(n_6615),
.Y(n_8423)
);

OAI21x1_ASAP7_75t_L g8424 ( 
.A1(n_6260),
.A2(n_6261),
.B(n_7069),
.Y(n_8424)
);

OAI22xp5_ASAP7_75t_L g8425 ( 
.A1(n_7318),
.A2(n_7681),
.B1(n_6615),
.B2(n_6310),
.Y(n_8425)
);

OAI21x1_ASAP7_75t_L g8426 ( 
.A1(n_6260),
.A2(n_7069),
.B(n_6254),
.Y(n_8426)
);

OAI22xp5_ASAP7_75t_L g8427 ( 
.A1(n_7318),
.A2(n_7681),
.B1(n_6615),
.B2(n_6356),
.Y(n_8427)
);

AOI21xp5_ASAP7_75t_L g8428 ( 
.A1(n_6400),
.A2(n_7355),
.B(n_7354),
.Y(n_8428)
);

NAND2x1p5_ASAP7_75t_L g8429 ( 
.A(n_7020),
.B(n_7308),
.Y(n_8429)
);

OAI21x1_ASAP7_75t_L g8430 ( 
.A1(n_7069),
.A2(n_6456),
.B(n_7238),
.Y(n_8430)
);

OAI21x1_ASAP7_75t_SL g8431 ( 
.A1(n_7638),
.A2(n_7419),
.B(n_6298),
.Y(n_8431)
);

OAI21xp5_ASAP7_75t_L g8432 ( 
.A1(n_7133),
.A2(n_6448),
.B(n_6330),
.Y(n_8432)
);

O2A1O1Ixp33_ASAP7_75t_SL g8433 ( 
.A1(n_7488),
.A2(n_7462),
.B(n_7440),
.C(n_7427),
.Y(n_8433)
);

OR2x2_ASAP7_75t_L g8434 ( 
.A(n_7472),
.B(n_7561),
.Y(n_8434)
);

NOR2x1_ASAP7_75t_L g8435 ( 
.A(n_7309),
.B(n_7394),
.Y(n_8435)
);

OAI22xp5_ASAP7_75t_L g8436 ( 
.A1(n_7318),
.A2(n_7681),
.B1(n_6356),
.B2(n_6396),
.Y(n_8436)
);

AOI22xp5_ASAP7_75t_L g8437 ( 
.A1(n_6478),
.A2(n_6513),
.B1(n_6469),
.B2(n_7457),
.Y(n_8437)
);

AOI21x1_ASAP7_75t_L g8438 ( 
.A1(n_6485),
.A2(n_6492),
.B(n_6489),
.Y(n_8438)
);

CKINVDCx20_ASAP7_75t_R g8439 ( 
.A(n_6648),
.Y(n_8439)
);

BUFx3_ASAP7_75t_L g8440 ( 
.A(n_7449),
.Y(n_8440)
);

NAND2xp5_ASAP7_75t_L g8441 ( 
.A(n_7584),
.B(n_7533),
.Y(n_8441)
);

BUFx3_ASAP7_75t_L g8442 ( 
.A(n_6772),
.Y(n_8442)
);

AND2x2_ASAP7_75t_L g8443 ( 
.A(n_6622),
.B(n_7566),
.Y(n_8443)
);

AOI31xp67_ASAP7_75t_L g8444 ( 
.A1(n_6320),
.A2(n_6337),
.A3(n_6348),
.B(n_6322),
.Y(n_8444)
);

AOI21xp5_ASAP7_75t_L g8445 ( 
.A1(n_7354),
.A2(n_7372),
.B(n_7355),
.Y(n_8445)
);

NAND2xp5_ASAP7_75t_SL g8446 ( 
.A(n_6495),
.B(n_7407),
.Y(n_8446)
);

AOI21xp5_ASAP7_75t_L g8447 ( 
.A1(n_7372),
.A2(n_7376),
.B(n_7375),
.Y(n_8447)
);

INVxp67_ASAP7_75t_L g8448 ( 
.A(n_7476),
.Y(n_8448)
);

INVx6_ASAP7_75t_L g8449 ( 
.A(n_6952),
.Y(n_8449)
);

OAI21x1_ASAP7_75t_L g8450 ( 
.A1(n_6456),
.A2(n_7240),
.B(n_6564),
.Y(n_8450)
);

AO31x2_ASAP7_75t_L g8451 ( 
.A1(n_6337),
.A2(n_6348),
.A3(n_6430),
.B(n_6366),
.Y(n_8451)
);

A2O1A1Ixp33_ASAP7_75t_L g8452 ( 
.A1(n_7317),
.A2(n_6298),
.B(n_6281),
.C(n_6520),
.Y(n_8452)
);

INVxp67_ASAP7_75t_L g8453 ( 
.A(n_7476),
.Y(n_8453)
);

AO22x2_ASAP7_75t_L g8454 ( 
.A1(n_7041),
.A2(n_7185),
.B1(n_6387),
.B2(n_6372),
.Y(n_8454)
);

AOI221x1_ASAP7_75t_L g8455 ( 
.A1(n_6760),
.A2(n_6835),
.B1(n_6369),
.B2(n_7411),
.C(n_7595),
.Y(n_8455)
);

AOI21xp5_ASAP7_75t_L g8456 ( 
.A1(n_7375),
.A2(n_7378),
.B(n_7376),
.Y(n_8456)
);

AOI21xp5_ASAP7_75t_SL g8457 ( 
.A1(n_6469),
.A2(n_6513),
.B(n_7440),
.Y(n_8457)
);

NOR2xp33_ASAP7_75t_SL g8458 ( 
.A(n_7190),
.B(n_6829),
.Y(n_8458)
);

A2O1A1Ixp33_ASAP7_75t_L g8459 ( 
.A1(n_6281),
.A2(n_6752),
.B(n_6985),
.C(n_6520),
.Y(n_8459)
);

INVx4_ASAP7_75t_L g8460 ( 
.A(n_6453),
.Y(n_8460)
);

INVx3_ASAP7_75t_L g8461 ( 
.A(n_7240),
.Y(n_8461)
);

NAND2xp5_ASAP7_75t_SL g8462 ( 
.A(n_6495),
.B(n_7407),
.Y(n_8462)
);

NAND2xp5_ASAP7_75t_SL g8463 ( 
.A(n_6495),
.B(n_7341),
.Y(n_8463)
);

NAND3x1_ASAP7_75t_L g8464 ( 
.A(n_7309),
.B(n_7391),
.C(n_6617),
.Y(n_8464)
);

AO21x2_ASAP7_75t_L g8465 ( 
.A1(n_6313),
.A2(n_6366),
.B(n_6348),
.Y(n_8465)
);

NAND3xp33_ASAP7_75t_SL g8466 ( 
.A(n_7093),
.B(n_7152),
.C(n_7136),
.Y(n_8466)
);

NAND2xp5_ASAP7_75t_L g8467 ( 
.A(n_7584),
.B(n_7533),
.Y(n_8467)
);

NOR2xp33_ASAP7_75t_L g8468 ( 
.A(n_7403),
.B(n_6340),
.Y(n_8468)
);

AOI21xp5_ASAP7_75t_L g8469 ( 
.A1(n_7378),
.A2(n_7393),
.B(n_7382),
.Y(n_8469)
);

O2A1O1Ixp33_ASAP7_75t_SL g8470 ( 
.A1(n_7462),
.A2(n_7427),
.B(n_6340),
.C(n_6579),
.Y(n_8470)
);

A2O1A1Ixp33_ASAP7_75t_L g8471 ( 
.A1(n_6520),
.A2(n_6985),
.B(n_7016),
.C(n_6752),
.Y(n_8471)
);

INVx5_ASAP7_75t_L g8472 ( 
.A(n_7183),
.Y(n_8472)
);

AOI22xp5_ASAP7_75t_L g8473 ( 
.A1(n_6513),
.A2(n_6469),
.B1(n_7493),
.B2(n_7457),
.Y(n_8473)
);

AOI21xp5_ASAP7_75t_L g8474 ( 
.A1(n_7382),
.A2(n_7405),
.B(n_7393),
.Y(n_8474)
);

AND2x2_ASAP7_75t_SL g8475 ( 
.A(n_7409),
.B(n_7423),
.Y(n_8475)
);

OAI21x1_ASAP7_75t_L g8476 ( 
.A1(n_7240),
.A2(n_6564),
.B(n_6430),
.Y(n_8476)
);

AOI21xp5_ASAP7_75t_L g8477 ( 
.A1(n_7405),
.A2(n_7417),
.B(n_7406),
.Y(n_8477)
);

AND2x2_ASAP7_75t_L g8478 ( 
.A(n_6622),
.B(n_7566),
.Y(n_8478)
);

NAND2xp5_ASAP7_75t_SL g8479 ( 
.A(n_6892),
.B(n_7394),
.Y(n_8479)
);

BUFx2_ASAP7_75t_L g8480 ( 
.A(n_7313),
.Y(n_8480)
);

NAND3xp33_ASAP7_75t_SL g8481 ( 
.A(n_7136),
.B(n_7152),
.C(n_6579),
.Y(n_8481)
);

NAND2xp5_ASAP7_75t_SL g8482 ( 
.A(n_7418),
.B(n_7391),
.Y(n_8482)
);

AO31x2_ASAP7_75t_L g8483 ( 
.A1(n_6366),
.A2(n_6476),
.A3(n_6496),
.B(n_6430),
.Y(n_8483)
);

BUFx3_ASAP7_75t_L g8484 ( 
.A(n_6772),
.Y(n_8484)
);

A2O1A1Ixp33_ASAP7_75t_L g8485 ( 
.A1(n_6520),
.A2(n_6985),
.B(n_7016),
.C(n_6752),
.Y(n_8485)
);

O2A1O1Ixp33_ASAP7_75t_SL g8486 ( 
.A1(n_6396),
.A2(n_6627),
.B(n_6684),
.C(n_6660),
.Y(n_8486)
);

OAI21xp5_ASAP7_75t_L g8487 ( 
.A1(n_6448),
.A2(n_6513),
.B(n_6482),
.Y(n_8487)
);

AOI21xp5_ASAP7_75t_L g8488 ( 
.A1(n_7406),
.A2(n_7425),
.B(n_7417),
.Y(n_8488)
);

OAI21x1_ASAP7_75t_L g8489 ( 
.A1(n_6564),
.A2(n_6496),
.B(n_7156),
.Y(n_8489)
);

OAI21x1_ASAP7_75t_L g8490 ( 
.A1(n_7156),
.A2(n_7220),
.B(n_7202),
.Y(n_8490)
);

OAI21x1_ASAP7_75t_L g8491 ( 
.A1(n_7156),
.A2(n_7220),
.B(n_7202),
.Y(n_8491)
);

A2O1A1Ixp33_ASAP7_75t_L g8492 ( 
.A1(n_6752),
.A2(n_7016),
.B(n_7153),
.C(n_6985),
.Y(n_8492)
);

NAND3xp33_ASAP7_75t_L g8493 ( 
.A(n_7361),
.B(n_7387),
.C(n_7640),
.Y(n_8493)
);

AOI21xp5_ASAP7_75t_L g8494 ( 
.A1(n_7425),
.A2(n_7435),
.B(n_7429),
.Y(n_8494)
);

AO21x2_ASAP7_75t_L g8495 ( 
.A1(n_6485),
.A2(n_6492),
.B(n_6489),
.Y(n_8495)
);

O2A1O1Ixp5_ASAP7_75t_L g8496 ( 
.A1(n_7265),
.A2(n_6482),
.B(n_7377),
.C(n_7297),
.Y(n_8496)
);

INVx6_ASAP7_75t_L g8497 ( 
.A(n_6952),
.Y(n_8497)
);

AOI21xp5_ASAP7_75t_SL g8498 ( 
.A1(n_6825),
.A2(n_6899),
.B(n_6826),
.Y(n_8498)
);

NAND2xp5_ASAP7_75t_L g8499 ( 
.A(n_7464),
.B(n_7473),
.Y(n_8499)
);

OAI21x1_ASAP7_75t_L g8500 ( 
.A1(n_7202),
.A2(n_7282),
.B(n_7220),
.Y(n_8500)
);

OA22x2_ASAP7_75t_L g8501 ( 
.A1(n_7654),
.A2(n_7493),
.B1(n_6746),
.B2(n_7041),
.Y(n_8501)
);

AOI21xp5_ASAP7_75t_L g8502 ( 
.A1(n_7429),
.A2(n_7436),
.B(n_7435),
.Y(n_8502)
);

AND2x2_ASAP7_75t_L g8503 ( 
.A(n_7566),
.B(n_7587),
.Y(n_8503)
);

INVx1_ASAP7_75t_SL g8504 ( 
.A(n_7198),
.Y(n_8504)
);

NAND2xp5_ASAP7_75t_L g8505 ( 
.A(n_7464),
.B(n_7473),
.Y(n_8505)
);

AOI221xp5_ASAP7_75t_SL g8506 ( 
.A1(n_7418),
.A2(n_6335),
.B1(n_6684),
.B2(n_6660),
.C(n_6627),
.Y(n_8506)
);

AOI21xp5_ASAP7_75t_L g8507 ( 
.A1(n_7436),
.A2(n_7439),
.B(n_7441),
.Y(n_8507)
);

AOI21x1_ASAP7_75t_L g8508 ( 
.A1(n_6485),
.A2(n_6492),
.B(n_6489),
.Y(n_8508)
);

NAND2x1p5_ASAP7_75t_L g8509 ( 
.A(n_7020),
.B(n_7308),
.Y(n_8509)
);

NAND2xp5_ASAP7_75t_L g8510 ( 
.A(n_7487),
.B(n_7494),
.Y(n_8510)
);

OAI22xp5_ASAP7_75t_L g8511 ( 
.A1(n_7681),
.A2(n_6848),
.B1(n_6920),
.B2(n_6722),
.Y(n_8511)
);

OAI22xp5_ASAP7_75t_L g8512 ( 
.A1(n_6722),
.A2(n_6920),
.B1(n_6848),
.B2(n_7016),
.Y(n_8512)
);

OA22x2_ASAP7_75t_L g8513 ( 
.A1(n_6746),
.A2(n_7677),
.B1(n_6609),
.B2(n_7349),
.Y(n_8513)
);

AOI21xp5_ASAP7_75t_SL g8514 ( 
.A1(n_6825),
.A2(n_6899),
.B(n_6826),
.Y(n_8514)
);

NOR2xp33_ASAP7_75t_L g8515 ( 
.A(n_7304),
.B(n_6335),
.Y(n_8515)
);

AOI21xp5_ASAP7_75t_L g8516 ( 
.A1(n_7439),
.A2(n_7441),
.B(n_7297),
.Y(n_8516)
);

INVx4_ASAP7_75t_L g8517 ( 
.A(n_6453),
.Y(n_8517)
);

AOI21x1_ASAP7_75t_L g8518 ( 
.A1(n_7327),
.A2(n_7047),
.B(n_7038),
.Y(n_8518)
);

O2A1O1Ixp33_ASAP7_75t_SL g8519 ( 
.A1(n_7524),
.A2(n_7550),
.B(n_7388),
.C(n_7184),
.Y(n_8519)
);

OR2x2_ASAP7_75t_L g8520 ( 
.A(n_7561),
.B(n_7092),
.Y(n_8520)
);

AOI21xp33_ASAP7_75t_L g8521 ( 
.A1(n_6522),
.A2(n_6536),
.B(n_6530),
.Y(n_8521)
);

NAND2xp5_ASAP7_75t_SL g8522 ( 
.A(n_7640),
.B(n_7153),
.Y(n_8522)
);

CKINVDCx5p33_ASAP7_75t_R g8523 ( 
.A(n_7332),
.Y(n_8523)
);

AO32x2_ASAP7_75t_L g8524 ( 
.A1(n_7369),
.A2(n_7614),
.A3(n_6483),
.B1(n_6573),
.B2(n_6384),
.Y(n_8524)
);

CKINVDCx5p33_ASAP7_75t_R g8525 ( 
.A(n_7370),
.Y(n_8525)
);

O2A1O1Ixp33_ASAP7_75t_SL g8526 ( 
.A1(n_7524),
.A2(n_7550),
.B(n_7388),
.C(n_7184),
.Y(n_8526)
);

OAI22x1_ASAP7_75t_L g8527 ( 
.A1(n_7409),
.A2(n_7480),
.B1(n_7519),
.B2(n_7423),
.Y(n_8527)
);

OAI21x1_ASAP7_75t_SL g8528 ( 
.A1(n_7419),
.A2(n_6609),
.B(n_7485),
.Y(n_8528)
);

NAND2xp5_ASAP7_75t_L g8529 ( 
.A(n_7487),
.B(n_7494),
.Y(n_8529)
);

AOI21xp5_ASAP7_75t_L g8530 ( 
.A1(n_7279),
.A2(n_7242),
.B(n_6453),
.Y(n_8530)
);

AOI21xp5_ASAP7_75t_L g8531 ( 
.A1(n_7279),
.A2(n_7242),
.B(n_6453),
.Y(n_8531)
);

OAI21x1_ASAP7_75t_L g8532 ( 
.A1(n_7282),
.A2(n_7299),
.B(n_7291),
.Y(n_8532)
);

AOI21xp5_ASAP7_75t_SL g8533 ( 
.A1(n_6825),
.A2(n_6899),
.B(n_6826),
.Y(n_8533)
);

AND2x2_ASAP7_75t_L g8534 ( 
.A(n_7566),
.B(n_7587),
.Y(n_8534)
);

NAND2xp5_ASAP7_75t_L g8535 ( 
.A(n_7496),
.B(n_7503),
.Y(n_8535)
);

NAND2xp5_ASAP7_75t_L g8536 ( 
.A(n_7496),
.B(n_7503),
.Y(n_8536)
);

BUFx2_ASAP7_75t_L g8537 ( 
.A(n_7313),
.Y(n_8537)
);

AOI21xp5_ASAP7_75t_L g8538 ( 
.A1(n_7242),
.A2(n_7337),
.B(n_7447),
.Y(n_8538)
);

AOI221x1_ASAP7_75t_L g8539 ( 
.A1(n_7682),
.A2(n_7501),
.B1(n_7513),
.B2(n_7508),
.C(n_6980),
.Y(n_8539)
);

NAND2xp5_ASAP7_75t_L g8540 ( 
.A(n_7504),
.B(n_7527),
.Y(n_8540)
);

AOI21xp5_ASAP7_75t_L g8541 ( 
.A1(n_7337),
.A2(n_7447),
.B(n_7265),
.Y(n_8541)
);

NAND2xp5_ASAP7_75t_SL g8542 ( 
.A(n_7153),
.B(n_7229),
.Y(n_8542)
);

AOI21xp5_ASAP7_75t_L g8543 ( 
.A1(n_7272),
.A2(n_7273),
.B(n_7583),
.Y(n_8543)
);

OAI21xp5_ASAP7_75t_L g8544 ( 
.A1(n_7112),
.A2(n_7114),
.B(n_7096),
.Y(n_8544)
);

NAND2xp5_ASAP7_75t_L g8545 ( 
.A(n_7504),
.B(n_7527),
.Y(n_8545)
);

NOR2xp33_ASAP7_75t_SL g8546 ( 
.A(n_6909),
.B(n_7383),
.Y(n_8546)
);

O2A1O1Ixp5_ASAP7_75t_L g8547 ( 
.A1(n_7377),
.A2(n_7500),
.B(n_7655),
.C(n_6980),
.Y(n_8547)
);

O2A1O1Ixp33_ASAP7_75t_L g8548 ( 
.A1(n_6530),
.A2(n_6549),
.B(n_6536),
.C(n_6609),
.Y(n_8548)
);

BUFx6f_ASAP7_75t_L g8549 ( 
.A(n_7020),
.Y(n_8549)
);

NAND2xp5_ASAP7_75t_L g8550 ( 
.A(n_7535),
.B(n_7575),
.Y(n_8550)
);

AOI22xp33_ASAP7_75t_L g8551 ( 
.A1(n_6909),
.A2(n_7383),
.B1(n_6617),
.B2(n_7209),
.Y(n_8551)
);

OAI21x1_ASAP7_75t_L g8552 ( 
.A1(n_7282),
.A2(n_7299),
.B(n_7291),
.Y(n_8552)
);

AOI21xp5_ASAP7_75t_L g8553 ( 
.A1(n_7272),
.A2(n_7273),
.B(n_7583),
.Y(n_8553)
);

AOI21xp5_ASAP7_75t_L g8554 ( 
.A1(n_7301),
.A2(n_7274),
.B(n_7505),
.Y(n_8554)
);

OAI21x1_ASAP7_75t_L g8555 ( 
.A1(n_7291),
.A2(n_7299),
.B(n_6345),
.Y(n_8555)
);

OAI21x1_ASAP7_75t_L g8556 ( 
.A1(n_6345),
.A2(n_7047),
.B(n_7038),
.Y(n_8556)
);

OAI21xp5_ASAP7_75t_L g8557 ( 
.A1(n_7112),
.A2(n_7114),
.B(n_7096),
.Y(n_8557)
);

CKINVDCx20_ASAP7_75t_R g8558 ( 
.A(n_7132),
.Y(n_8558)
);

AOI21xp33_ASAP7_75t_L g8559 ( 
.A1(n_6549),
.A2(n_6611),
.B(n_6408),
.Y(n_8559)
);

AOI221xp5_ASAP7_75t_L g8560 ( 
.A1(n_7185),
.A2(n_7538),
.B1(n_7485),
.B2(n_7571),
.C(n_7650),
.Y(n_8560)
);

A2O1A1Ixp33_ASAP7_75t_L g8561 ( 
.A1(n_7153),
.A2(n_7229),
.B(n_7298),
.C(n_7507),
.Y(n_8561)
);

OAI21x1_ASAP7_75t_L g8562 ( 
.A1(n_7038),
.A2(n_7047),
.B(n_7415),
.Y(n_8562)
);

NAND2xp5_ASAP7_75t_L g8563 ( 
.A(n_7535),
.B(n_7575),
.Y(n_8563)
);

NOR2xp33_ASAP7_75t_L g8564 ( 
.A(n_7304),
.B(n_7278),
.Y(n_8564)
);

NAND2xp5_ASAP7_75t_L g8565 ( 
.A(n_7579),
.B(n_7278),
.Y(n_8565)
);

AO31x2_ASAP7_75t_L g8566 ( 
.A1(n_7239),
.A2(n_7521),
.A3(n_7448),
.B(n_7471),
.Y(n_8566)
);

AO31x2_ASAP7_75t_L g8567 ( 
.A1(n_7442),
.A2(n_7471),
.A3(n_7482),
.B(n_7448),
.Y(n_8567)
);

OAI22xp5_ASAP7_75t_L g8568 ( 
.A1(n_7229),
.A2(n_6867),
.B1(n_6557),
.B2(n_6560),
.Y(n_8568)
);

O2A1O1Ixp5_ASAP7_75t_L g8569 ( 
.A1(n_7377),
.A2(n_7500),
.B(n_7655),
.C(n_7428),
.Y(n_8569)
);

A2O1A1Ixp33_ASAP7_75t_L g8570 ( 
.A1(n_7229),
.A2(n_7298),
.B(n_7507),
.C(n_7099),
.Y(n_8570)
);

NOR4xp25_ASAP7_75t_L g8571 ( 
.A(n_7349),
.B(n_7387),
.C(n_7361),
.D(n_6429),
.Y(n_8571)
);

OAI21x1_ASAP7_75t_L g8572 ( 
.A1(n_7415),
.A2(n_7420),
.B(n_7075),
.Y(n_8572)
);

AOI221x1_ASAP7_75t_L g8573 ( 
.A1(n_7508),
.A2(n_7301),
.B1(n_7349),
.B2(n_7538),
.C(n_7623),
.Y(n_8573)
);

OAI21xp33_ASAP7_75t_L g8574 ( 
.A1(n_7650),
.A2(n_7104),
.B(n_7099),
.Y(n_8574)
);

AO21x1_ASAP7_75t_L g8575 ( 
.A1(n_7159),
.A2(n_7266),
.B(n_6611),
.Y(n_8575)
);

OAI21xp5_ASAP7_75t_SL g8576 ( 
.A1(n_6617),
.A2(n_7677),
.B(n_7673),
.Y(n_8576)
);

AOI21xp5_ASAP7_75t_L g8577 ( 
.A1(n_7274),
.A2(n_7505),
.B(n_7020),
.Y(n_8577)
);

OAI21x1_ASAP7_75t_L g8578 ( 
.A1(n_7415),
.A2(n_7420),
.B(n_7075),
.Y(n_8578)
);

INVxp67_ASAP7_75t_SL g8579 ( 
.A(n_7247),
.Y(n_8579)
);

AOI21xp5_ASAP7_75t_L g8580 ( 
.A1(n_7348),
.A2(n_7360),
.B(n_7308),
.Y(n_8580)
);

BUFx6f_ASAP7_75t_L g8581 ( 
.A(n_7308),
.Y(n_8581)
);

OAI21x1_ASAP7_75t_L g8582 ( 
.A1(n_7420),
.A2(n_7075),
.B(n_6599),
.Y(n_8582)
);

AOI21xp5_ASAP7_75t_L g8583 ( 
.A1(n_7360),
.A2(n_7348),
.B(n_6303),
.Y(n_8583)
);

AOI21xp5_ASAP7_75t_L g8584 ( 
.A1(n_7360),
.A2(n_7348),
.B(n_6303),
.Y(n_8584)
);

AO31x2_ASAP7_75t_L g8585 ( 
.A1(n_7442),
.A2(n_7471),
.A3(n_7482),
.B(n_7448),
.Y(n_8585)
);

AND2x2_ASAP7_75t_L g8586 ( 
.A(n_7587),
.B(n_7561),
.Y(n_8586)
);

NOR2xp33_ASAP7_75t_L g8587 ( 
.A(n_6407),
.B(n_6429),
.Y(n_8587)
);

AOI21xp5_ASAP7_75t_L g8588 ( 
.A1(n_7348),
.A2(n_7360),
.B(n_6303),
.Y(n_8588)
);

OAI22xp5_ASAP7_75t_L g8589 ( 
.A1(n_6867),
.A2(n_6552),
.B1(n_6560),
.B2(n_6557),
.Y(n_8589)
);

AOI21xp5_ASAP7_75t_L g8590 ( 
.A1(n_7348),
.A2(n_7360),
.B(n_6303),
.Y(n_8590)
);

INVx1_ASAP7_75t_L g8591 ( 
.A(n_7319),
.Y(n_8591)
);

OAI22xp5_ASAP7_75t_L g8592 ( 
.A1(n_6563),
.A2(n_6566),
.B1(n_6568),
.B2(n_6567),
.Y(n_8592)
);

INVx1_ASAP7_75t_L g8593 ( 
.A(n_7319),
.Y(n_8593)
);

A2O1A1Ixp33_ASAP7_75t_L g8594 ( 
.A1(n_7104),
.A2(n_6611),
.B(n_7480),
.C(n_7409),
.Y(n_8594)
);

INVx1_ASAP7_75t_L g8595 ( 
.A(n_7319),
.Y(n_8595)
);

AOI21xp5_ASAP7_75t_L g8596 ( 
.A1(n_7348),
.A2(n_7360),
.B(n_6303),
.Y(n_8596)
);

AND2x2_ASAP7_75t_L g8597 ( 
.A(n_7587),
.B(n_7105),
.Y(n_8597)
);

OAI21xp5_ASAP7_75t_L g8598 ( 
.A1(n_6278),
.A2(n_6517),
.B(n_6508),
.Y(n_8598)
);

A2O1A1Ixp33_ASAP7_75t_L g8599 ( 
.A1(n_7480),
.A2(n_7519),
.B(n_7410),
.C(n_7075),
.Y(n_8599)
);

AOI21x1_ASAP7_75t_L g8600 ( 
.A1(n_7327),
.A2(n_7495),
.B(n_7470),
.Y(n_8600)
);

OAI21x1_ASAP7_75t_L g8601 ( 
.A1(n_6565),
.A2(n_6599),
.B(n_7095),
.Y(n_8601)
);

OAI21xp5_ASAP7_75t_L g8602 ( 
.A1(n_6278),
.A2(n_6517),
.B(n_6508),
.Y(n_8602)
);

AOI21xp5_ASAP7_75t_L g8603 ( 
.A1(n_7348),
.A2(n_7360),
.B(n_6303),
.Y(n_8603)
);

OAI21xp5_ASAP7_75t_L g8604 ( 
.A1(n_6278),
.A2(n_6517),
.B(n_6508),
.Y(n_8604)
);

OAI21xp5_ASAP7_75t_L g8605 ( 
.A1(n_6517),
.A2(n_6610),
.B(n_7433),
.Y(n_8605)
);

OAI21x1_ASAP7_75t_SL g8606 ( 
.A1(n_7485),
.A2(n_7571),
.B(n_6447),
.Y(n_8606)
);

BUFx2_ASAP7_75t_L g8607 ( 
.A(n_7313),
.Y(n_8607)
);

BUFx12f_ASAP7_75t_L g8608 ( 
.A(n_7045),
.Y(n_8608)
);

OAI21xp5_ASAP7_75t_L g8609 ( 
.A1(n_6610),
.A2(n_7433),
.B(n_7470),
.Y(n_8609)
);

OAI21x1_ASAP7_75t_L g8610 ( 
.A1(n_6565),
.A2(n_6599),
.B(n_7095),
.Y(n_8610)
);

NOR2xp67_ASAP7_75t_SL g8611 ( 
.A(n_7383),
.B(n_7045),
.Y(n_8611)
);

INVx1_ASAP7_75t_SL g8612 ( 
.A(n_7198),
.Y(n_8612)
);

NAND3xp33_ASAP7_75t_L g8613 ( 
.A(n_6407),
.B(n_6626),
.C(n_6582),
.Y(n_8613)
);

AOI221xp5_ASAP7_75t_SL g8614 ( 
.A1(n_6633),
.A2(n_7022),
.B1(n_6942),
.B2(n_6703),
.C(n_7262),
.Y(n_8614)
);

OAI22x1_ASAP7_75t_L g8615 ( 
.A1(n_7519),
.A2(n_7051),
.B1(n_7196),
.B2(n_6882),
.Y(n_8615)
);

OAI21x1_ASAP7_75t_L g8616 ( 
.A1(n_6565),
.A2(n_7498),
.B(n_7495),
.Y(n_8616)
);

AND2x4_ASAP7_75t_L g8617 ( 
.A(n_7232),
.B(n_7348),
.Y(n_8617)
);

INVxp67_ASAP7_75t_L g8618 ( 
.A(n_7571),
.Y(n_8618)
);

NAND2xp5_ASAP7_75t_SL g8619 ( 
.A(n_7661),
.B(n_7673),
.Y(n_8619)
);

OR2x2_ASAP7_75t_L g8620 ( 
.A(n_7092),
.B(n_7127),
.Y(n_8620)
);

AOI21xp5_ASAP7_75t_L g8621 ( 
.A1(n_7348),
.A2(n_7360),
.B(n_6357),
.Y(n_8621)
);

OAI21xp5_ASAP7_75t_L g8622 ( 
.A1(n_6610),
.A2(n_7498),
.B(n_6353),
.Y(n_8622)
);

INVx2_ASAP7_75t_SL g8623 ( 
.A(n_7469),
.Y(n_8623)
);

AOI21xp5_ASAP7_75t_L g8624 ( 
.A1(n_7348),
.A2(n_7360),
.B(n_6357),
.Y(n_8624)
);

BUFx6f_ASAP7_75t_L g8625 ( 
.A(n_7360),
.Y(n_8625)
);

AOI22xp5_ASAP7_75t_L g8626 ( 
.A1(n_7383),
.A2(n_7209),
.B1(n_7045),
.B2(n_6408),
.Y(n_8626)
);

AOI21xp5_ASAP7_75t_L g8627 ( 
.A1(n_6357),
.A2(n_6384),
.B(n_6287),
.Y(n_8627)
);

AOI21xp5_ASAP7_75t_L g8628 ( 
.A1(n_6357),
.A2(n_6384),
.B(n_6287),
.Y(n_8628)
);

OAI22xp5_ASAP7_75t_L g8629 ( 
.A1(n_6586),
.A2(n_6591),
.B1(n_7661),
.B2(n_7062),
.Y(n_8629)
);

AOI21xp5_ASAP7_75t_L g8630 ( 
.A1(n_6357),
.A2(n_6384),
.B(n_6287),
.Y(n_8630)
);

OAI21x1_ASAP7_75t_L g8631 ( 
.A1(n_7126),
.A2(n_7129),
.B(n_6382),
.Y(n_8631)
);

OR2x2_ASAP7_75t_L g8632 ( 
.A(n_7092),
.B(n_7127),
.Y(n_8632)
);

A2O1A1Ixp33_ASAP7_75t_L g8633 ( 
.A1(n_7410),
.A2(n_7656),
.B(n_6610),
.C(n_7052),
.Y(n_8633)
);

CKINVDCx5p33_ASAP7_75t_R g8634 ( 
.A(n_7370),
.Y(n_8634)
);

OAI21xp5_ASAP7_75t_L g8635 ( 
.A1(n_6353),
.A2(n_6296),
.B(n_6293),
.Y(n_8635)
);

INVx3_ASAP7_75t_SL g8636 ( 
.A(n_6291),
.Y(n_8636)
);

OAI21x1_ASAP7_75t_L g8637 ( 
.A1(n_7126),
.A2(n_7129),
.B(n_6382),
.Y(n_8637)
);

AND2x2_ASAP7_75t_L g8638 ( 
.A(n_7105),
.B(n_6661),
.Y(n_8638)
);

INVx1_ASAP7_75t_SL g8639 ( 
.A(n_7221),
.Y(n_8639)
);

NOR4xp25_ASAP7_75t_L g8640 ( 
.A(n_6626),
.B(n_6591),
.C(n_7062),
.D(n_7644),
.Y(n_8640)
);

OAI22xp5_ASAP7_75t_L g8641 ( 
.A1(n_7289),
.A2(n_7295),
.B1(n_7296),
.B2(n_7438),
.Y(n_8641)
);

OA21x2_ASAP7_75t_L g8642 ( 
.A1(n_7363),
.A2(n_7365),
.B(n_7129),
.Y(n_8642)
);

OAI22xp5_ASAP7_75t_L g8643 ( 
.A1(n_7289),
.A2(n_7295),
.B1(n_7296),
.B2(n_7438),
.Y(n_8643)
);

INVx2_ASAP7_75t_L g8644 ( 
.A(n_7468),
.Y(n_8644)
);

CKINVDCx11_ASAP7_75t_R g8645 ( 
.A(n_7045),
.Y(n_8645)
);

NAND2xp5_ASAP7_75t_L g8646 ( 
.A(n_7627),
.B(n_7629),
.Y(n_8646)
);

CKINVDCx20_ASAP7_75t_R g8647 ( 
.A(n_7132),
.Y(n_8647)
);

CKINVDCx11_ASAP7_75t_R g8648 ( 
.A(n_7209),
.Y(n_8648)
);

OAI22x1_ASAP7_75t_L g8649 ( 
.A1(n_6882),
.A2(n_7196),
.B1(n_7340),
.B2(n_7051),
.Y(n_8649)
);

CKINVDCx5p33_ASAP7_75t_R g8650 ( 
.A(n_7404),
.Y(n_8650)
);

OAI21x1_ASAP7_75t_L g8651 ( 
.A1(n_7126),
.A2(n_7129),
.B(n_6382),
.Y(n_8651)
);

AO21x1_ASAP7_75t_L g8652 ( 
.A1(n_7159),
.A2(n_7266),
.B(n_7310),
.Y(n_8652)
);

INVx1_ASAP7_75t_SL g8653 ( 
.A(n_7221),
.Y(n_8653)
);

OAI21x1_ASAP7_75t_L g8654 ( 
.A1(n_7126),
.A2(n_6376),
.B(n_7363),
.Y(n_8654)
);

OAI21x1_ASAP7_75t_L g8655 ( 
.A1(n_6376),
.A2(n_7365),
.B(n_7363),
.Y(n_8655)
);

AOI21xp5_ASAP7_75t_L g8656 ( 
.A1(n_6357),
.A2(n_6483),
.B(n_6287),
.Y(n_8656)
);

OAI22xp5_ASAP7_75t_L g8657 ( 
.A1(n_7443),
.A2(n_7455),
.B1(n_7458),
.B2(n_7644),
.Y(n_8657)
);

OAI21x1_ASAP7_75t_L g8658 ( 
.A1(n_6376),
.A2(n_7365),
.B(n_7252),
.Y(n_8658)
);

A2O1A1Ixp33_ASAP7_75t_L g8659 ( 
.A1(n_7656),
.A2(n_7052),
.B(n_7604),
.C(n_6762),
.Y(n_8659)
);

INVx3_ASAP7_75t_SL g8660 ( 
.A(n_6291),
.Y(n_8660)
);

O2A1O1Ixp5_ASAP7_75t_L g8661 ( 
.A1(n_6772),
.A2(n_7428),
.B(n_7327),
.C(n_7585),
.Y(n_8661)
);

O2A1O1Ixp33_ASAP7_75t_L g8662 ( 
.A1(n_7185),
.A2(n_6447),
.B(n_6302),
.C(n_6433),
.Y(n_8662)
);

NOR2xp33_ASAP7_75t_R g8663 ( 
.A(n_6612),
.B(n_7404),
.Y(n_8663)
);

OAI21x1_ASAP7_75t_L g8664 ( 
.A1(n_7247),
.A2(n_7259),
.B(n_7252),
.Y(n_8664)
);

AOI21xp5_ASAP7_75t_L g8665 ( 
.A1(n_6483),
.A2(n_6707),
.B(n_6573),
.Y(n_8665)
);

OAI21xp33_ASAP7_75t_L g8666 ( 
.A1(n_7627),
.A2(n_7634),
.B(n_7629),
.Y(n_8666)
);

NAND2xp5_ASAP7_75t_L g8667 ( 
.A(n_7634),
.B(n_7635),
.Y(n_8667)
);

OAI21xp5_ASAP7_75t_L g8668 ( 
.A1(n_6353),
.A2(n_6299),
.B(n_6296),
.Y(n_8668)
);

A2O1A1Ixp33_ASAP7_75t_L g8669 ( 
.A1(n_7656),
.A2(n_7052),
.B(n_7604),
.C(n_6762),
.Y(n_8669)
);

AOI21xp5_ASAP7_75t_L g8670 ( 
.A1(n_6483),
.A2(n_6707),
.B(n_6573),
.Y(n_8670)
);

CKINVDCx5p33_ASAP7_75t_R g8671 ( 
.A(n_7484),
.Y(n_8671)
);

OAI21x1_ASAP7_75t_L g8672 ( 
.A1(n_7247),
.A2(n_7259),
.B(n_7252),
.Y(n_8672)
);

A2O1A1Ixp33_ASAP7_75t_L g8673 ( 
.A1(n_7656),
.A2(n_7052),
.B(n_6762),
.C(n_6923),
.Y(n_8673)
);

BUFx2_ASAP7_75t_L g8674 ( 
.A(n_7313),
.Y(n_8674)
);

INVx6_ASAP7_75t_L g8675 ( 
.A(n_7581),
.Y(n_8675)
);

NAND2xp5_ASAP7_75t_L g8676 ( 
.A(n_7635),
.B(n_7641),
.Y(n_8676)
);

OAI22xp5_ASAP7_75t_L g8677 ( 
.A1(n_7443),
.A2(n_7455),
.B1(n_7458),
.B2(n_7461),
.Y(n_8677)
);

OAI21x1_ASAP7_75t_L g8678 ( 
.A1(n_7247),
.A2(n_7259),
.B(n_7252),
.Y(n_8678)
);

O2A1O1Ixp5_ASAP7_75t_L g8679 ( 
.A1(n_7428),
.A2(n_7605),
.B(n_7617),
.C(n_7424),
.Y(n_8679)
);

OAI21xp5_ASAP7_75t_L g8680 ( 
.A1(n_6353),
.A2(n_6296),
.B(n_6293),
.Y(n_8680)
);

AND2x2_ASAP7_75t_L g8681 ( 
.A(n_7105),
.B(n_6661),
.Y(n_8681)
);

NAND2xp5_ASAP7_75t_L g8682 ( 
.A(n_7641),
.B(n_7645),
.Y(n_8682)
);

INVx3_ASAP7_75t_L g8683 ( 
.A(n_7413),
.Y(n_8683)
);

INVx3_ASAP7_75t_L g8684 ( 
.A(n_7413),
.Y(n_8684)
);

CKINVDCx5p33_ASAP7_75t_R g8685 ( 
.A(n_7484),
.Y(n_8685)
);

A2O1A1Ixp33_ASAP7_75t_L g8686 ( 
.A1(n_7052),
.A2(n_6762),
.B(n_6344),
.C(n_7621),
.Y(n_8686)
);

AND2x2_ASAP7_75t_L g8687 ( 
.A(n_7105),
.B(n_6661),
.Y(n_8687)
);

NAND2xp33_ASAP7_75t_L g8688 ( 
.A(n_7525),
.B(n_6629),
.Y(n_8688)
);

AO32x2_ASAP7_75t_L g8689 ( 
.A1(n_7614),
.A2(n_6887),
.A3(n_6916),
.B1(n_6707),
.B2(n_6573),
.Y(n_8689)
);

OAI21x1_ASAP7_75t_L g8690 ( 
.A1(n_7259),
.A2(n_7277),
.B(n_7264),
.Y(n_8690)
);

AOI21x1_ASAP7_75t_L g8691 ( 
.A1(n_7451),
.A2(n_7351),
.B(n_7246),
.Y(n_8691)
);

AOI21x1_ASAP7_75t_L g8692 ( 
.A1(n_7451),
.A2(n_7351),
.B(n_7246),
.Y(n_8692)
);

A2O1A1Ixp33_ASAP7_75t_L g8693 ( 
.A1(n_7052),
.A2(n_6762),
.B(n_6344),
.C(n_7621),
.Y(n_8693)
);

AND2x2_ASAP7_75t_L g8694 ( 
.A(n_6661),
.B(n_6664),
.Y(n_8694)
);

OAI22xp5_ASAP7_75t_L g8695 ( 
.A1(n_7461),
.A2(n_7645),
.B1(n_7209),
.B2(n_7466),
.Y(n_8695)
);

OAI21x1_ASAP7_75t_L g8696 ( 
.A1(n_7264),
.A2(n_7287),
.B(n_7277),
.Y(n_8696)
);

AOI21xp5_ASAP7_75t_L g8697 ( 
.A1(n_6707),
.A2(n_6916),
.B(n_6887),
.Y(n_8697)
);

O2A1O1Ixp5_ASAP7_75t_L g8698 ( 
.A1(n_7605),
.A2(n_7617),
.B(n_7424),
.C(n_6607),
.Y(n_8698)
);

NAND2x1p5_ASAP7_75t_L g8699 ( 
.A(n_6291),
.B(n_6312),
.Y(n_8699)
);

AO31x2_ASAP7_75t_L g8700 ( 
.A1(n_6667),
.A2(n_6714),
.A3(n_6715),
.B(n_6702),
.Y(n_8700)
);

BUFx6f_ASAP7_75t_L g8701 ( 
.A(n_6259),
.Y(n_8701)
);

AOI21xp5_ASAP7_75t_L g8702 ( 
.A1(n_6887),
.A2(n_6916),
.B(n_7510),
.Y(n_8702)
);

O2A1O1Ixp33_ASAP7_75t_L g8703 ( 
.A1(n_6447),
.A2(n_6302),
.B(n_6433),
.C(n_6255),
.Y(n_8703)
);

INVx2_ASAP7_75t_L g8704 ( 
.A(n_7468),
.Y(n_8704)
);

A2O1A1Ixp33_ASAP7_75t_L g8705 ( 
.A1(n_7052),
.A2(n_6762),
.B(n_7621),
.C(n_7657),
.Y(n_8705)
);

CKINVDCx20_ASAP7_75t_R g8706 ( 
.A(n_7525),
.Y(n_8706)
);

OAI21x1_ASAP7_75t_L g8707 ( 
.A1(n_7264),
.A2(n_7287),
.B(n_7277),
.Y(n_8707)
);

NAND2xp5_ASAP7_75t_SL g8708 ( 
.A(n_7678),
.B(n_7683),
.Y(n_8708)
);

AOI21xp5_ASAP7_75t_L g8709 ( 
.A1(n_6887),
.A2(n_6916),
.B(n_7603),
.Y(n_8709)
);

BUFx6f_ASAP7_75t_L g8710 ( 
.A(n_6259),
.Y(n_8710)
);

AO31x2_ASAP7_75t_L g8711 ( 
.A1(n_6667),
.A2(n_6714),
.A3(n_6715),
.B(n_6702),
.Y(n_8711)
);

AOI21xp5_ASAP7_75t_L g8712 ( 
.A1(n_7611),
.A2(n_7309),
.B(n_6531),
.Y(n_8712)
);

AO31x2_ASAP7_75t_L g8713 ( 
.A1(n_6715),
.A2(n_6724),
.A3(n_6742),
.B(n_6725),
.Y(n_8713)
);

NAND3xp33_ASAP7_75t_L g8714 ( 
.A(n_7483),
.B(n_6703),
.C(n_6633),
.Y(n_8714)
);

INVxp67_ASAP7_75t_SL g8715 ( 
.A(n_7264),
.Y(n_8715)
);

AND2x4_ASAP7_75t_L g8716 ( 
.A(n_6580),
.B(n_6607),
.Y(n_8716)
);

NAND3xp33_ASAP7_75t_L g8717 ( 
.A(n_7483),
.B(n_7022),
.C(n_6942),
.Y(n_8717)
);

AND2x2_ASAP7_75t_L g8718 ( 
.A(n_6664),
.B(n_6701),
.Y(n_8718)
);

OAI21x1_ASAP7_75t_L g8719 ( 
.A1(n_7277),
.A2(n_7292),
.B(n_7287),
.Y(n_8719)
);

CKINVDCx20_ASAP7_75t_R g8720 ( 
.A(n_6629),
.Y(n_8720)
);

OAI21x1_ASAP7_75t_L g8721 ( 
.A1(n_7287),
.A2(n_7293),
.B(n_7292),
.Y(n_8721)
);

AOI21xp33_ASAP7_75t_L g8722 ( 
.A1(n_6408),
.A2(n_6405),
.B(n_6397),
.Y(n_8722)
);

OAI21x1_ASAP7_75t_L g8723 ( 
.A1(n_7292),
.A2(n_7293),
.B(n_7490),
.Y(n_8723)
);

OAI21x1_ASAP7_75t_L g8724 ( 
.A1(n_7292),
.A2(n_7293),
.B(n_7490),
.Y(n_8724)
);

CKINVDCx5p33_ASAP7_75t_R g8725 ( 
.A(n_6838),
.Y(n_8725)
);

O2A1O1Ixp5_ASAP7_75t_L g8726 ( 
.A1(n_7424),
.A2(n_6607),
.B(n_6644),
.C(n_6580),
.Y(n_8726)
);

AOI221x1_ASAP7_75t_L g8727 ( 
.A1(n_7623),
.A2(n_7625),
.B1(n_7658),
.B2(n_7653),
.C(n_7632),
.Y(n_8727)
);

OAI21x1_ASAP7_75t_SL g8728 ( 
.A1(n_7664),
.A2(n_7668),
.B(n_7322),
.Y(n_8728)
);

INVx2_ASAP7_75t_L g8729 ( 
.A(n_7468),
.Y(n_8729)
);

AOI21xp5_ASAP7_75t_L g8730 ( 
.A1(n_6531),
.A2(n_7490),
.B(n_6312),
.Y(n_8730)
);

OAI21xp5_ASAP7_75t_L g8731 ( 
.A1(n_6293),
.A2(n_6299),
.B(n_6296),
.Y(n_8731)
);

AOI221x1_ASAP7_75t_L g8732 ( 
.A1(n_7623),
.A2(n_7625),
.B1(n_7658),
.B2(n_7653),
.C(n_7632),
.Y(n_8732)
);

NAND2xp5_ASAP7_75t_L g8733 ( 
.A(n_7652),
.B(n_7310),
.Y(n_8733)
);

BUFx3_ASAP7_75t_L g8734 ( 
.A(n_6732),
.Y(n_8734)
);

NAND3xp33_ASAP7_75t_L g8735 ( 
.A(n_7322),
.B(n_7342),
.C(n_7326),
.Y(n_8735)
);

AOI21xp5_ASAP7_75t_L g8736 ( 
.A1(n_6531),
.A2(n_7490),
.B(n_6312),
.Y(n_8736)
);

NAND2xp33_ASAP7_75t_R g8737 ( 
.A(n_7610),
.B(n_7631),
.Y(n_8737)
);

BUFx6f_ASAP7_75t_L g8738 ( 
.A(n_6259),
.Y(n_8738)
);

AOI21x1_ASAP7_75t_L g8739 ( 
.A1(n_7451),
.A2(n_7351),
.B(n_7246),
.Y(n_8739)
);

AND2x4_ASAP7_75t_L g8740 ( 
.A(n_6580),
.B(n_6607),
.Y(n_8740)
);

AOI21x1_ASAP7_75t_L g8741 ( 
.A1(n_7246),
.A2(n_7351),
.B(n_7398),
.Y(n_8741)
);

BUFx12f_ASAP7_75t_L g8742 ( 
.A(n_6838),
.Y(n_8742)
);

NAND2xp5_ASAP7_75t_L g8743 ( 
.A(n_7652),
.B(n_7326),
.Y(n_8743)
);

AND2x4_ASAP7_75t_L g8744 ( 
.A(n_6580),
.B(n_6607),
.Y(n_8744)
);

BUFx3_ASAP7_75t_L g8745 ( 
.A(n_6732),
.Y(n_8745)
);

AOI211x1_ASAP7_75t_L g8746 ( 
.A1(n_7598),
.A2(n_7345),
.B(n_7357),
.C(n_7678),
.Y(n_8746)
);

NAND2xp5_ASAP7_75t_L g8747 ( 
.A(n_7652),
.B(n_7342),
.Y(n_8747)
);

OAI21x1_ASAP7_75t_L g8748 ( 
.A1(n_7293),
.A2(n_7490),
.B(n_6325),
.Y(n_8748)
);

INVx4_ASAP7_75t_L g8749 ( 
.A(n_6832),
.Y(n_8749)
);

AOI21xp5_ASAP7_75t_L g8750 ( 
.A1(n_6291),
.A2(n_6324),
.B(n_6312),
.Y(n_8750)
);

AOI211x1_ASAP7_75t_L g8751 ( 
.A1(n_7598),
.A2(n_7357),
.B(n_7345),
.C(n_7683),
.Y(n_8751)
);

AOI22xp5_ASAP7_75t_L g8752 ( 
.A1(n_6408),
.A2(n_6284),
.B1(n_7033),
.B2(n_6551),
.Y(n_8752)
);

A2O1A1Ixp33_ASAP7_75t_L g8753 ( 
.A1(n_7052),
.A2(n_6762),
.B(n_7621),
.C(n_7657),
.Y(n_8753)
);

NAND3xp33_ASAP7_75t_L g8754 ( 
.A(n_6255),
.B(n_6486),
.C(n_7072),
.Y(n_8754)
);

AND2x2_ASAP7_75t_L g8755 ( 
.A(n_6664),
.B(n_6701),
.Y(n_8755)
);

AND2x2_ASAP7_75t_L g8756 ( 
.A(n_6664),
.B(n_6701),
.Y(n_8756)
);

CKINVDCx5p33_ASAP7_75t_R g8757 ( 
.A(n_6840),
.Y(n_8757)
);

O2A1O1Ixp5_ASAP7_75t_L g8758 ( 
.A1(n_6580),
.A2(n_6644),
.B(n_6713),
.C(n_6607),
.Y(n_8758)
);

AND2x2_ASAP7_75t_L g8759 ( 
.A(n_6701),
.B(n_6721),
.Y(n_8759)
);

BUFx2_ASAP7_75t_L g8760 ( 
.A(n_7313),
.Y(n_8760)
);

A2O1A1Ixp33_ASAP7_75t_L g8761 ( 
.A1(n_7052),
.A2(n_6762),
.B(n_7657),
.C(n_7340),
.Y(n_8761)
);

NOR2xp33_ASAP7_75t_SL g8762 ( 
.A(n_7033),
.B(n_7460),
.Y(n_8762)
);

AO31x2_ASAP7_75t_L g8763 ( 
.A1(n_6724),
.A2(n_6725),
.A3(n_6786),
.B(n_6742),
.Y(n_8763)
);

BUFx2_ASAP7_75t_L g8764 ( 
.A(n_7313),
.Y(n_8764)
);

AO21x1_ASAP7_75t_L g8765 ( 
.A1(n_6724),
.A2(n_6742),
.B(n_6725),
.Y(n_8765)
);

A2O1A1Ixp33_ASAP7_75t_L g8766 ( 
.A1(n_6762),
.A2(n_7657),
.B(n_7092),
.C(n_7672),
.Y(n_8766)
);

INVx5_ASAP7_75t_L g8767 ( 
.A(n_6732),
.Y(n_8767)
);

AND2x2_ASAP7_75t_SL g8768 ( 
.A(n_6644),
.B(n_6713),
.Y(n_8768)
);

A2O1A1Ixp33_ASAP7_75t_L g8769 ( 
.A1(n_7092),
.A2(n_7672),
.B(n_7679),
.C(n_7676),
.Y(n_8769)
);

NAND3xp33_ASAP7_75t_SL g8770 ( 
.A(n_6840),
.B(n_7668),
.C(n_7664),
.Y(n_8770)
);

AOI21xp5_ASAP7_75t_L g8771 ( 
.A1(n_6291),
.A2(n_6324),
.B(n_6312),
.Y(n_8771)
);

AOI21xp5_ASAP7_75t_L g8772 ( 
.A1(n_6312),
.A2(n_6419),
.B(n_6324),
.Y(n_8772)
);

AOI21xp5_ASAP7_75t_L g8773 ( 
.A1(n_6324),
.A2(n_6426),
.B(n_6419),
.Y(n_8773)
);

BUFx2_ASAP7_75t_L g8774 ( 
.A(n_7313),
.Y(n_8774)
);

OAI22xp5_ASAP7_75t_L g8775 ( 
.A1(n_7463),
.A2(n_7474),
.B1(n_7477),
.B2(n_7466),
.Y(n_8775)
);

OAI21x1_ASAP7_75t_SL g8776 ( 
.A1(n_7033),
.A2(n_7398),
.B(n_6713),
.Y(n_8776)
);

A2O1A1Ixp33_ASAP7_75t_L g8777 ( 
.A1(n_7092),
.A2(n_7676),
.B(n_7679),
.C(n_7672),
.Y(n_8777)
);

AOI21xp5_ASAP7_75t_L g8778 ( 
.A1(n_6324),
.A2(n_6426),
.B(n_6419),
.Y(n_8778)
);

AOI221xp5_ASAP7_75t_SL g8779 ( 
.A1(n_7072),
.A2(n_7262),
.B1(n_7148),
.B2(n_7121),
.C(n_7516),
.Y(n_8779)
);

BUFx2_ASAP7_75t_L g8780 ( 
.A(n_7313),
.Y(n_8780)
);

AOI221xp5_ASAP7_75t_L g8781 ( 
.A1(n_7379),
.A2(n_7390),
.B1(n_7397),
.B2(n_7389),
.C(n_7385),
.Y(n_8781)
);

A2O1A1Ixp33_ASAP7_75t_L g8782 ( 
.A1(n_7092),
.A2(n_7676),
.B(n_7679),
.C(n_7672),
.Y(n_8782)
);

AOI221xp5_ASAP7_75t_SL g8783 ( 
.A1(n_7121),
.A2(n_7148),
.B1(n_7567),
.B2(n_7599),
.C(n_7516),
.Y(n_8783)
);

OAI21xp5_ASAP7_75t_L g8784 ( 
.A1(n_6293),
.A2(n_6299),
.B(n_6414),
.Y(n_8784)
);

OAI21xp5_ASAP7_75t_L g8785 ( 
.A1(n_6299),
.A2(n_6420),
.B(n_6414),
.Y(n_8785)
);

NAND2xp5_ASAP7_75t_L g8786 ( 
.A(n_7652),
.B(n_7628),
.Y(n_8786)
);

OAI21xp5_ASAP7_75t_L g8787 ( 
.A1(n_6414),
.A2(n_6432),
.B(n_6420),
.Y(n_8787)
);

NAND2xp5_ASAP7_75t_L g8788 ( 
.A(n_7628),
.B(n_7633),
.Y(n_8788)
);

AOI21x1_ASAP7_75t_SL g8789 ( 
.A1(n_6551),
.A2(n_6486),
.B(n_6387),
.Y(n_8789)
);

NAND2xp5_ASAP7_75t_L g8790 ( 
.A(n_7628),
.B(n_7633),
.Y(n_8790)
);

NAND2xp5_ASAP7_75t_L g8791 ( 
.A(n_7628),
.B(n_7633),
.Y(n_8791)
);

INVx2_ASAP7_75t_L g8792 ( 
.A(n_7468),
.Y(n_8792)
);

OAI22xp5_ASAP7_75t_L g8793 ( 
.A1(n_7463),
.A2(n_7477),
.B1(n_7486),
.B2(n_7474),
.Y(n_8793)
);

NAND2xp5_ASAP7_75t_L g8794 ( 
.A(n_7633),
.B(n_7637),
.Y(n_8794)
);

OAI22xp5_ASAP7_75t_L g8795 ( 
.A1(n_7486),
.A2(n_7518),
.B1(n_7520),
.B2(n_7492),
.Y(n_8795)
);

CKINVDCx20_ASAP7_75t_R g8796 ( 
.A(n_7446),
.Y(n_8796)
);

AOI21x1_ASAP7_75t_L g8797 ( 
.A1(n_7351),
.A2(n_7398),
.B(n_6510),
.Y(n_8797)
);

NAND2xp5_ASAP7_75t_L g8798 ( 
.A(n_7637),
.B(n_7643),
.Y(n_8798)
);

BUFx2_ASAP7_75t_L g8799 ( 
.A(n_7313),
.Y(n_8799)
);

AOI21xp5_ASAP7_75t_L g8800 ( 
.A1(n_6324),
.A2(n_6426),
.B(n_6419),
.Y(n_8800)
);

NAND3xp33_ASAP7_75t_L g8801 ( 
.A(n_7624),
.B(n_7400),
.C(n_7674),
.Y(n_8801)
);

AOI21xp5_ASAP7_75t_L g8802 ( 
.A1(n_6419),
.A2(n_6461),
.B(n_6426),
.Y(n_8802)
);

NAND2xp5_ASAP7_75t_L g8803 ( 
.A(n_7637),
.B(n_7643),
.Y(n_8803)
);

NAND3x1_ASAP7_75t_L g8804 ( 
.A(n_6274),
.B(n_6538),
.C(n_6399),
.Y(n_8804)
);

AOI21xp5_ASAP7_75t_L g8805 ( 
.A1(n_6419),
.A2(n_6461),
.B(n_6426),
.Y(n_8805)
);

NAND2xp5_ASAP7_75t_L g8806 ( 
.A(n_7637),
.B(n_7643),
.Y(n_8806)
);

OAI21xp5_ASAP7_75t_L g8807 ( 
.A1(n_6414),
.A2(n_6432),
.B(n_6420),
.Y(n_8807)
);

OAI22xp5_ASAP7_75t_L g8808 ( 
.A1(n_7492),
.A2(n_7520),
.B1(n_7518),
.B2(n_6397),
.Y(n_8808)
);

OAI21xp5_ASAP7_75t_L g8809 ( 
.A1(n_6420),
.A2(n_6446),
.B(n_6432),
.Y(n_8809)
);

OA21x2_ASAP7_75t_L g8810 ( 
.A1(n_7367),
.A2(n_7374),
.B(n_7414),
.Y(n_8810)
);

NAND2xp5_ASAP7_75t_L g8811 ( 
.A(n_7643),
.B(n_7651),
.Y(n_8811)
);

NAND2xp5_ASAP7_75t_L g8812 ( 
.A(n_7651),
.B(n_7600),
.Y(n_8812)
);

NAND2xp5_ASAP7_75t_L g8813 ( 
.A(n_7651),
.B(n_7600),
.Y(n_8813)
);

CKINVDCx6p67_ASAP7_75t_R g8814 ( 
.A(n_7622),
.Y(n_8814)
);

BUFx3_ASAP7_75t_L g8815 ( 
.A(n_6732),
.Y(n_8815)
);

OR2x2_ASAP7_75t_L g8816 ( 
.A(n_7092),
.B(n_7333),
.Y(n_8816)
);

AO22x2_ASAP7_75t_L g8817 ( 
.A1(n_6372),
.A2(n_6387),
.B1(n_6284),
.B2(n_6551),
.Y(n_8817)
);

OAI22xp5_ASAP7_75t_L g8818 ( 
.A1(n_6397),
.A2(n_6405),
.B1(n_7622),
.B2(n_7366),
.Y(n_8818)
);

AO31x2_ASAP7_75t_L g8819 ( 
.A1(n_6786),
.A2(n_6799),
.A3(n_6865),
.B(n_6789),
.Y(n_8819)
);

AOI22xp5_ASAP7_75t_L g8820 ( 
.A1(n_6408),
.A2(n_6284),
.B1(n_7033),
.B2(n_6551),
.Y(n_8820)
);

BUFx3_ASAP7_75t_L g8821 ( 
.A(n_6732),
.Y(n_8821)
);

INVxp67_ASAP7_75t_L g8822 ( 
.A(n_7624),
.Y(n_8822)
);

NAND4xp25_ASAP7_75t_L g8823 ( 
.A(n_6405),
.B(n_7366),
.C(n_7362),
.D(n_7619),
.Y(n_8823)
);

AND2x2_ASAP7_75t_L g8824 ( 
.A(n_6721),
.B(n_6778),
.Y(n_8824)
);

NAND2xp5_ASAP7_75t_L g8825 ( 
.A(n_7651),
.B(n_7600),
.Y(n_8825)
);

BUFx3_ASAP7_75t_L g8826 ( 
.A(n_6732),
.Y(n_8826)
);

A2O1A1Ixp33_ASAP7_75t_L g8827 ( 
.A1(n_7092),
.A2(n_7679),
.B(n_7676),
.C(n_6372),
.Y(n_8827)
);

NAND2x1_ASAP7_75t_L g8828 ( 
.A(n_7536),
.B(n_7545),
.Y(n_8828)
);

AOI21xp5_ASAP7_75t_L g8829 ( 
.A1(n_6426),
.A2(n_6477),
.B(n_6461),
.Y(n_8829)
);

NOR2x1_ASAP7_75t_SL g8830 ( 
.A(n_7536),
.B(n_7545),
.Y(n_8830)
);

AOI21xp5_ASAP7_75t_L g8831 ( 
.A1(n_6461),
.A2(n_6477),
.B(n_7536),
.Y(n_8831)
);

AOI21x1_ASAP7_75t_L g8832 ( 
.A1(n_7351),
.A2(n_6510),
.B(n_7517),
.Y(n_8832)
);

INVx2_ASAP7_75t_L g8833 ( 
.A(n_7522),
.Y(n_8833)
);

A2O1A1Ixp33_ASAP7_75t_L g8834 ( 
.A1(n_6372),
.A2(n_6387),
.B(n_6744),
.C(n_6377),
.Y(n_8834)
);

NAND2xp5_ASAP7_75t_SL g8835 ( 
.A(n_6387),
.B(n_6259),
.Y(n_8835)
);

AOI21xp5_ASAP7_75t_L g8836 ( 
.A1(n_6461),
.A2(n_6477),
.B(n_7536),
.Y(n_8836)
);

NAND2x1_ASAP7_75t_L g8837 ( 
.A(n_7536),
.B(n_7545),
.Y(n_8837)
);

NAND2xp5_ASAP7_75t_L g8838 ( 
.A(n_7600),
.B(n_7619),
.Y(n_8838)
);

O2A1O1Ixp5_ASAP7_75t_SL g8839 ( 
.A1(n_6786),
.A2(n_6799),
.B(n_6865),
.C(n_6789),
.Y(n_8839)
);

A2O1A1Ixp33_ASAP7_75t_L g8840 ( 
.A1(n_6387),
.A2(n_6744),
.B(n_6377),
.C(n_6365),
.Y(n_8840)
);

OAI22xp5_ASAP7_75t_L g8841 ( 
.A1(n_7622),
.A2(n_7362),
.B1(n_7333),
.B2(n_7379),
.Y(n_8841)
);

AOI21xp5_ASAP7_75t_L g8842 ( 
.A1(n_6461),
.A2(n_6477),
.B(n_7536),
.Y(n_8842)
);

AOI21xp5_ASAP7_75t_L g8843 ( 
.A1(n_6477),
.A2(n_7545),
.B(n_7536),
.Y(n_8843)
);

OAI21xp5_ASAP7_75t_L g8844 ( 
.A1(n_6432),
.A2(n_6457),
.B(n_6446),
.Y(n_8844)
);

AND2x2_ASAP7_75t_L g8845 ( 
.A(n_6721),
.B(n_6778),
.Y(n_8845)
);

AOI22xp5_ASAP7_75t_L g8846 ( 
.A1(n_6408),
.A2(n_7033),
.B1(n_6551),
.B2(n_6826),
.Y(n_8846)
);

OAI21x1_ASAP7_75t_L g8847 ( 
.A1(n_6341),
.A2(n_6343),
.B(n_6365),
.Y(n_8847)
);

NAND2xp5_ASAP7_75t_L g8848 ( 
.A(n_7564),
.B(n_7385),
.Y(n_8848)
);

AOI21xp5_ASAP7_75t_L g8849 ( 
.A1(n_6477),
.A2(n_7545),
.B(n_7351),
.Y(n_8849)
);

INVx3_ASAP7_75t_L g8850 ( 
.A(n_7414),
.Y(n_8850)
);

AOI21xp5_ASAP7_75t_L g8851 ( 
.A1(n_7545),
.A2(n_7400),
.B(n_6808),
.Y(n_8851)
);

NAND2xp5_ASAP7_75t_L g8852 ( 
.A(n_7564),
.B(n_7389),
.Y(n_8852)
);

AO32x2_ASAP7_75t_L g8853 ( 
.A1(n_7338),
.A2(n_7347),
.A3(n_7531),
.B1(n_7460),
.B2(n_6644),
.Y(n_8853)
);

AND2x2_ASAP7_75t_L g8854 ( 
.A(n_6721),
.B(n_6778),
.Y(n_8854)
);

OR2x2_ASAP7_75t_L g8855 ( 
.A(n_7333),
.B(n_7564),
.Y(n_8855)
);

OAI21x1_ASAP7_75t_L g8856 ( 
.A1(n_6341),
.A2(n_6343),
.B(n_6365),
.Y(n_8856)
);

O2A1O1Ixp5_ASAP7_75t_L g8857 ( 
.A1(n_6644),
.A2(n_6713),
.B(n_7674),
.C(n_7347),
.Y(n_8857)
);

AOI22xp5_ASAP7_75t_L g8858 ( 
.A1(n_7033),
.A2(n_6551),
.B1(n_6826),
.B2(n_6825),
.Y(n_8858)
);

AND2x2_ASAP7_75t_L g8859 ( 
.A(n_6778),
.B(n_6783),
.Y(n_8859)
);

AND2x4_ASAP7_75t_L g8860 ( 
.A(n_6713),
.B(n_7545),
.Y(n_8860)
);

O2A1O1Ixp33_ASAP7_75t_L g8861 ( 
.A1(n_7601),
.A2(n_7632),
.B(n_7653),
.C(n_7625),
.Y(n_8861)
);

OA21x2_ASAP7_75t_L g8862 ( 
.A1(n_7367),
.A2(n_7374),
.B(n_6343),
.Y(n_8862)
);

OAI21x1_ASAP7_75t_L g8863 ( 
.A1(n_6341),
.A2(n_6343),
.B(n_6377),
.Y(n_8863)
);

OAI21x1_ASAP7_75t_L g8864 ( 
.A1(n_7367),
.A2(n_7374),
.B(n_7147),
.Y(n_8864)
);

OAI21x1_ASAP7_75t_L g8865 ( 
.A1(n_7367),
.A2(n_7374),
.B(n_7147),
.Y(n_8865)
);

NAND2xp5_ASAP7_75t_L g8866 ( 
.A(n_7564),
.B(n_7390),
.Y(n_8866)
);

INVx5_ASAP7_75t_L g8867 ( 
.A(n_6259),
.Y(n_8867)
);

AOI21xp5_ASAP7_75t_L g8868 ( 
.A1(n_7400),
.A2(n_6808),
.B(n_6784),
.Y(n_8868)
);

AOI21xp5_ASAP7_75t_L g8869 ( 
.A1(n_7400),
.A2(n_6808),
.B(n_6784),
.Y(n_8869)
);

AO31x2_ASAP7_75t_L g8870 ( 
.A1(n_6789),
.A2(n_6865),
.A3(n_6895),
.B(n_6799),
.Y(n_8870)
);

A2O1A1Ixp33_ASAP7_75t_L g8871 ( 
.A1(n_6744),
.A2(n_6411),
.B(n_7662),
.C(n_7646),
.Y(n_8871)
);

OAI21xp33_ASAP7_75t_L g8872 ( 
.A1(n_7397),
.A2(n_7416),
.B(n_7401),
.Y(n_8872)
);

OAI21x1_ASAP7_75t_L g8873 ( 
.A1(n_7145),
.A2(n_7147),
.B(n_6412),
.Y(n_8873)
);

BUFx2_ASAP7_75t_L g8874 ( 
.A(n_7300),
.Y(n_8874)
);

AO21x1_ASAP7_75t_L g8875 ( 
.A1(n_6895),
.A2(n_6914),
.B(n_6906),
.Y(n_8875)
);

NAND2x1_ASAP7_75t_L g8876 ( 
.A(n_6825),
.B(n_6826),
.Y(n_8876)
);

AOI21xp5_ASAP7_75t_L g8877 ( 
.A1(n_7400),
.A2(n_6808),
.B(n_6784),
.Y(n_8877)
);

INVx6_ASAP7_75t_L g8878 ( 
.A(n_7581),
.Y(n_8878)
);

AOI21xp5_ASAP7_75t_L g8879 ( 
.A1(n_7400),
.A2(n_6808),
.B(n_6784),
.Y(n_8879)
);

AND2x2_ASAP7_75t_L g8880 ( 
.A(n_6783),
.B(n_6816),
.Y(n_8880)
);

CKINVDCx20_ASAP7_75t_R g8881 ( 
.A(n_7446),
.Y(n_8881)
);

OAI21x1_ASAP7_75t_L g8882 ( 
.A1(n_7145),
.A2(n_7147),
.B(n_6412),
.Y(n_8882)
);

OAI21x1_ASAP7_75t_L g8883 ( 
.A1(n_7145),
.A2(n_6412),
.B(n_6398),
.Y(n_8883)
);

NOR2xp67_ASAP7_75t_L g8884 ( 
.A(n_6274),
.B(n_6399),
.Y(n_8884)
);

NOR2xp33_ASAP7_75t_L g8885 ( 
.A(n_7665),
.B(n_7356),
.Y(n_8885)
);

AOI21xp5_ASAP7_75t_L g8886 ( 
.A1(n_7400),
.A2(n_6850),
.B(n_6784),
.Y(n_8886)
);

AOI31xp67_ASAP7_75t_L g8887 ( 
.A1(n_7647),
.A2(n_6750),
.A3(n_6759),
.B(n_6716),
.Y(n_8887)
);

AOI22xp5_ASAP7_75t_L g8888 ( 
.A1(n_6825),
.A2(n_6826),
.B1(n_6899),
.B2(n_6338),
.Y(n_8888)
);

OAI21xp5_ASAP7_75t_L g8889 ( 
.A1(n_6446),
.A2(n_6471),
.B(n_6457),
.Y(n_8889)
);

OAI21xp5_ASAP7_75t_L g8890 ( 
.A1(n_6446),
.A2(n_6471),
.B(n_6457),
.Y(n_8890)
);

NOR2xp67_ASAP7_75t_L g8891 ( 
.A(n_6274),
.B(n_6399),
.Y(n_8891)
);

AOI21xp5_ASAP7_75t_L g8892 ( 
.A1(n_6850),
.A2(n_6919),
.B(n_6852),
.Y(n_8892)
);

NOR2xp33_ASAP7_75t_L g8893 ( 
.A(n_7665),
.B(n_7356),
.Y(n_8893)
);

AOI22xp33_ASAP7_75t_SL g8894 ( 
.A1(n_6558),
.A2(n_6683),
.B1(n_6756),
.B2(n_6744),
.Y(n_8894)
);

NAND2x1p5_ASAP7_75t_L g8895 ( 
.A(n_7338),
.B(n_7347),
.Y(n_8895)
);

OAI21x1_ASAP7_75t_L g8896 ( 
.A1(n_7145),
.A2(n_6412),
.B(n_6398),
.Y(n_8896)
);

NAND2xp5_ASAP7_75t_L g8897 ( 
.A(n_7421),
.B(n_7565),
.Y(n_8897)
);

OAI21x1_ASAP7_75t_L g8898 ( 
.A1(n_6398),
.A2(n_6413),
.B(n_7155),
.Y(n_8898)
);

NAND3x1_ASAP7_75t_L g8899 ( 
.A(n_6274),
.B(n_6538),
.C(n_6399),
.Y(n_8899)
);

OAI21xp33_ASAP7_75t_L g8900 ( 
.A1(n_7421),
.A2(n_7620),
.B(n_7601),
.Y(n_8900)
);

OAI21x1_ASAP7_75t_L g8901 ( 
.A1(n_6398),
.A2(n_6413),
.B(n_7155),
.Y(n_8901)
);

NAND2xp5_ASAP7_75t_SL g8902 ( 
.A(n_6388),
.B(n_6516),
.Y(n_8902)
);

AO31x2_ASAP7_75t_L g8903 ( 
.A1(n_6895),
.A2(n_6914),
.A3(n_6921),
.B(n_6906),
.Y(n_8903)
);

BUFx3_ASAP7_75t_L g8904 ( 
.A(n_7300),
.Y(n_8904)
);

OAI21x1_ASAP7_75t_L g8905 ( 
.A1(n_6413),
.A2(n_7158),
.B(n_7155),
.Y(n_8905)
);

NAND2xp5_ASAP7_75t_L g8906 ( 
.A(n_7565),
.B(n_7580),
.Y(n_8906)
);

NAND2xp5_ASAP7_75t_L g8907 ( 
.A(n_7565),
.B(n_7580),
.Y(n_8907)
);

NAND2xp5_ASAP7_75t_L g8908 ( 
.A(n_7565),
.B(n_7580),
.Y(n_8908)
);

OAI21xp5_ASAP7_75t_L g8909 ( 
.A1(n_6457),
.A2(n_6473),
.B(n_6471),
.Y(n_8909)
);

OAI21xp5_ASAP7_75t_L g8910 ( 
.A1(n_6471),
.A2(n_6474),
.B(n_6473),
.Y(n_8910)
);

OR2x2_ASAP7_75t_L g8911 ( 
.A(n_7116),
.B(n_6744),
.Y(n_8911)
);

OAI22xp5_ASAP7_75t_L g8912 ( 
.A1(n_7622),
.A2(n_7620),
.B1(n_7599),
.B2(n_7567),
.Y(n_8912)
);

AO31x2_ASAP7_75t_L g8913 ( 
.A1(n_6906),
.A2(n_6921),
.A3(n_6924),
.B(n_6914),
.Y(n_8913)
);

NAND2x1p5_ASAP7_75t_L g8914 ( 
.A(n_7338),
.B(n_7347),
.Y(n_8914)
);

AOI21xp5_ASAP7_75t_L g8915 ( 
.A1(n_6850),
.A2(n_6919),
.B(n_6852),
.Y(n_8915)
);

AO31x2_ASAP7_75t_L g8916 ( 
.A1(n_6921),
.A2(n_6927),
.A3(n_6937),
.B(n_6924),
.Y(n_8916)
);

NAND2xp5_ASAP7_75t_L g8917 ( 
.A(n_7580),
.B(n_7589),
.Y(n_8917)
);

OAI21x1_ASAP7_75t_L g8918 ( 
.A1(n_6413),
.A2(n_7158),
.B(n_7155),
.Y(n_8918)
);

AOI221x1_ASAP7_75t_L g8919 ( 
.A1(n_7658),
.A2(n_7666),
.B1(n_7680),
.B2(n_7669),
.C(n_7663),
.Y(n_8919)
);

AO31x2_ASAP7_75t_L g8920 ( 
.A1(n_6924),
.A2(n_6937),
.A3(n_6953),
.B(n_6927),
.Y(n_8920)
);

NAND2xp5_ASAP7_75t_L g8921 ( 
.A(n_7589),
.B(n_7594),
.Y(n_8921)
);

OAI21x1_ASAP7_75t_L g8922 ( 
.A1(n_7158),
.A2(n_7172),
.B(n_7170),
.Y(n_8922)
);

OAI21x1_ASAP7_75t_L g8923 ( 
.A1(n_7158),
.A2(n_7172),
.B(n_7170),
.Y(n_8923)
);

AOI21xp5_ASAP7_75t_L g8924 ( 
.A1(n_6850),
.A2(n_6919),
.B(n_6852),
.Y(n_8924)
);

NOR2xp33_ASAP7_75t_L g8925 ( 
.A(n_7665),
.B(n_7386),
.Y(n_8925)
);

NAND2xp5_ASAP7_75t_L g8926 ( 
.A(n_7589),
.B(n_7594),
.Y(n_8926)
);

NAND2xp5_ASAP7_75t_L g8927 ( 
.A(n_7589),
.B(n_7594),
.Y(n_8927)
);

CKINVDCx20_ASAP7_75t_R g8928 ( 
.A(n_7446),
.Y(n_8928)
);

INVx2_ASAP7_75t_L g8929 ( 
.A(n_7522),
.Y(n_8929)
);

AO31x2_ASAP7_75t_L g8930 ( 
.A1(n_6927),
.A2(n_6953),
.A3(n_6963),
.B(n_6937),
.Y(n_8930)
);

OR2x2_ASAP7_75t_L g8931 ( 
.A(n_7116),
.B(n_6744),
.Y(n_8931)
);

NOR2xp67_ASAP7_75t_L g8932 ( 
.A(n_6274),
.B(n_6399),
.Y(n_8932)
);

NAND3xp33_ASAP7_75t_L g8933 ( 
.A(n_6953),
.B(n_6972),
.C(n_6963),
.Y(n_8933)
);

AOI22xp33_ASAP7_75t_L g8934 ( 
.A1(n_6558),
.A2(n_6683),
.B1(n_6826),
.B2(n_6825),
.Y(n_8934)
);

O2A1O1Ixp33_ASAP7_75t_L g8935 ( 
.A1(n_7659),
.A2(n_7663),
.B(n_7622),
.C(n_7666),
.Y(n_8935)
);

NAND2xp5_ASAP7_75t_L g8936 ( 
.A(n_7594),
.B(n_7602),
.Y(n_8936)
);

NAND2xp5_ASAP7_75t_L g8937 ( 
.A(n_7602),
.B(n_7606),
.Y(n_8937)
);

OAI21x1_ASAP7_75t_L g8938 ( 
.A1(n_7170),
.A2(n_7173),
.B(n_7172),
.Y(n_8938)
);

O2A1O1Ixp33_ASAP7_75t_L g8939 ( 
.A1(n_7659),
.A2(n_7669),
.B(n_7680),
.C(n_7647),
.Y(n_8939)
);

NAND2xp5_ASAP7_75t_L g8940 ( 
.A(n_7602),
.B(n_7606),
.Y(n_8940)
);

AOI21x1_ASAP7_75t_L g8941 ( 
.A1(n_7517),
.A2(n_7547),
.B(n_7542),
.Y(n_8941)
);

NOR2xp33_ASAP7_75t_L g8942 ( 
.A(n_7386),
.B(n_7422),
.Y(n_8942)
);

OR2x6_ASAP7_75t_L g8943 ( 
.A(n_6825),
.B(n_6899),
.Y(n_8943)
);

A2O1A1Ixp33_ASAP7_75t_L g8944 ( 
.A1(n_6744),
.A2(n_6411),
.B(n_7662),
.C(n_7646),
.Y(n_8944)
);

OAI21x1_ASAP7_75t_L g8945 ( 
.A1(n_7170),
.A2(n_7173),
.B(n_7172),
.Y(n_8945)
);

NAND3xp33_ASAP7_75t_SL g8946 ( 
.A(n_6850),
.B(n_6919),
.C(n_6852),
.Y(n_8946)
);

OAI21x1_ASAP7_75t_L g8947 ( 
.A1(n_7173),
.A2(n_7182),
.B(n_7176),
.Y(n_8947)
);

INVx2_ASAP7_75t_L g8948 ( 
.A(n_7522),
.Y(n_8948)
);

AOI21xp5_ASAP7_75t_L g8949 ( 
.A1(n_6852),
.A2(n_7023),
.B(n_6919),
.Y(n_8949)
);

OAI21x1_ASAP7_75t_L g8950 ( 
.A1(n_7173),
.A2(n_7182),
.B(n_7176),
.Y(n_8950)
);

NOR2xp67_ASAP7_75t_L g8951 ( 
.A(n_6274),
.B(n_6399),
.Y(n_8951)
);

NAND2xp5_ASAP7_75t_L g8952 ( 
.A(n_7602),
.B(n_7606),
.Y(n_8952)
);

NAND2xp5_ASAP7_75t_L g8953 ( 
.A(n_7602),
.B(n_7606),
.Y(n_8953)
);

OAI21x1_ASAP7_75t_L g8954 ( 
.A1(n_7176),
.A2(n_7205),
.B(n_7182),
.Y(n_8954)
);

INVxp67_ASAP7_75t_SL g8955 ( 
.A(n_7381),
.Y(n_8955)
);

OAI21x1_ASAP7_75t_L g8956 ( 
.A1(n_7176),
.A2(n_7205),
.B(n_7182),
.Y(n_8956)
);

NAND2xp5_ASAP7_75t_SL g8957 ( 
.A(n_6388),
.B(n_6516),
.Y(n_8957)
);

NAND3x1_ASAP7_75t_L g8958 ( 
.A(n_6538),
.B(n_6597),
.C(n_6585),
.Y(n_8958)
);

AOI21xp5_ASAP7_75t_L g8959 ( 
.A1(n_7023),
.A2(n_7201),
.B(n_7084),
.Y(n_8959)
);

NAND2xp5_ASAP7_75t_L g8960 ( 
.A(n_7602),
.B(n_7615),
.Y(n_8960)
);

OAI22xp5_ASAP7_75t_L g8961 ( 
.A1(n_6899),
.A2(n_7570),
.B1(n_7578),
.B2(n_7555),
.Y(n_8961)
);

CKINVDCx5p33_ASAP7_75t_R g8962 ( 
.A(n_7446),
.Y(n_8962)
);

A2O1A1Ixp33_ASAP7_75t_L g8963 ( 
.A1(n_6744),
.A2(n_6411),
.B(n_6474),
.C(n_6473),
.Y(n_8963)
);

OAI21x1_ASAP7_75t_L g8964 ( 
.A1(n_7205),
.A2(n_7219),
.B(n_7212),
.Y(n_8964)
);

OAI21x1_ASAP7_75t_L g8965 ( 
.A1(n_7205),
.A2(n_7219),
.B(n_7212),
.Y(n_8965)
);

AOI21xp5_ASAP7_75t_L g8966 ( 
.A1(n_7023),
.A2(n_7201),
.B(n_7084),
.Y(n_8966)
);

NAND2xp5_ASAP7_75t_SL g8967 ( 
.A(n_6388),
.B(n_6516),
.Y(n_8967)
);

OAI22x1_ASAP7_75t_L g8968 ( 
.A1(n_7610),
.A2(n_7631),
.B1(n_7011),
.B2(n_7049),
.Y(n_8968)
);

NAND2xp5_ASAP7_75t_L g8969 ( 
.A(n_7602),
.B(n_7615),
.Y(n_8969)
);

OAI21x1_ASAP7_75t_L g8970 ( 
.A1(n_7212),
.A2(n_7223),
.B(n_7219),
.Y(n_8970)
);

INVx2_ASAP7_75t_L g8971 ( 
.A(n_7522),
.Y(n_8971)
);

AOI22xp5_ASAP7_75t_L g8972 ( 
.A1(n_6899),
.A2(n_6338),
.B1(n_6512),
.B2(n_6507),
.Y(n_8972)
);

NAND3xp33_ASAP7_75t_L g8973 ( 
.A(n_6983),
.B(n_7049),
.C(n_7011),
.Y(n_8973)
);

NAND2xp5_ASAP7_75t_L g8974 ( 
.A(n_7602),
.B(n_7615),
.Y(n_8974)
);

NOR2xp33_ASAP7_75t_L g8975 ( 
.A(n_7874),
.B(n_7809),
.Y(n_8975)
);

NAND3xp33_ASAP7_75t_L g8976 ( 
.A(n_7786),
.B(n_7071),
.C(n_7063),
.Y(n_8976)
);

BUFx2_ASAP7_75t_L g8977 ( 
.A(n_8853),
.Y(n_8977)
);

OAI21x1_ASAP7_75t_L g8978 ( 
.A1(n_7844),
.A2(n_7873),
.B(n_8348),
.Y(n_8978)
);

INVx1_ASAP7_75t_L g8979 ( 
.A(n_8700),
.Y(n_8979)
);

AO21x1_ASAP7_75t_L g8980 ( 
.A1(n_7832),
.A2(n_7071),
.B(n_7063),
.Y(n_8980)
);

INVx2_ASAP7_75t_SL g8981 ( 
.A(n_8867),
.Y(n_8981)
);

INVxp67_ASAP7_75t_SL g8982 ( 
.A(n_8652),
.Y(n_8982)
);

OAI21x1_ASAP7_75t_L g8983 ( 
.A1(n_7873),
.A2(n_7582),
.B(n_7103),
.Y(n_8983)
);

NAND3xp33_ASAP7_75t_L g8984 ( 
.A(n_7786),
.B(n_7073),
.C(n_7071),
.Y(n_8984)
);

INVx2_ASAP7_75t_L g8985 ( 
.A(n_8887),
.Y(n_8985)
);

INVx2_ASAP7_75t_L g8986 ( 
.A(n_8887),
.Y(n_8986)
);

INVx1_ASAP7_75t_L g8987 ( 
.A(n_8700),
.Y(n_8987)
);

OR2x6_ASAP7_75t_L g8988 ( 
.A(n_8498),
.B(n_6899),
.Y(n_8988)
);

INVx1_ASAP7_75t_L g8989 ( 
.A(n_8700),
.Y(n_8989)
);

AO21x2_ASAP7_75t_L g8990 ( 
.A1(n_7975),
.A2(n_7384),
.B(n_7102),
.Y(n_8990)
);

OAI21x1_ASAP7_75t_L g8991 ( 
.A1(n_7873),
.A2(n_8348),
.B(n_8033),
.Y(n_8991)
);

AOI22x1_ASAP7_75t_L g8992 ( 
.A1(n_8006),
.A2(n_7084),
.B1(n_7201),
.B2(n_7023),
.Y(n_8992)
);

INVx1_ASAP7_75t_L g8993 ( 
.A(n_8700),
.Y(n_8993)
);

XNOR2xp5_ASAP7_75t_L g8994 ( 
.A(n_7891),
.B(n_7422),
.Y(n_8994)
);

NAND3xp33_ASAP7_75t_L g8995 ( 
.A(n_7742),
.B(n_7102),
.C(n_7073),
.Y(n_8995)
);

INVx1_ASAP7_75t_L g8996 ( 
.A(n_8700),
.Y(n_8996)
);

AND2x4_ASAP7_75t_L g8997 ( 
.A(n_8867),
.B(n_7469),
.Y(n_8997)
);

AO31x2_ASAP7_75t_L g8998 ( 
.A1(n_7991),
.A2(n_7102),
.A3(n_7115),
.B(n_7073),
.Y(n_8998)
);

AO21x2_ASAP7_75t_L g8999 ( 
.A1(n_7975),
.A2(n_7384),
.B(n_7137),
.Y(n_8999)
);

INVx1_ASAP7_75t_L g9000 ( 
.A(n_8700),
.Y(n_9000)
);

INVx1_ASAP7_75t_SL g9001 ( 
.A(n_8642),
.Y(n_9001)
);

OAI21x1_ASAP7_75t_L g9002 ( 
.A1(n_8010),
.A2(n_8030),
.B(n_8352),
.Y(n_9002)
);

AO21x1_ASAP7_75t_L g9003 ( 
.A1(n_7832),
.A2(n_8011),
.B(n_8069),
.Y(n_9003)
);

BUFx3_ASAP7_75t_L g9004 ( 
.A(n_8098),
.Y(n_9004)
);

INVx6_ASAP7_75t_L g9005 ( 
.A(n_7735),
.Y(n_9005)
);

INVx2_ASAP7_75t_L g9006 ( 
.A(n_8887),
.Y(n_9006)
);

OAI22xp33_ASAP7_75t_L g9007 ( 
.A1(n_7716),
.A2(n_7549),
.B1(n_7531),
.B2(n_7460),
.Y(n_9007)
);

BUFx2_ASAP7_75t_L g9008 ( 
.A(n_8853),
.Y(n_9008)
);

AOI22xp33_ASAP7_75t_L g9009 ( 
.A1(n_7809),
.A2(n_6683),
.B1(n_6558),
.B2(n_6970),
.Y(n_9009)
);

NOR2xp33_ASAP7_75t_SL g9010 ( 
.A(n_8006),
.B(n_6756),
.Y(n_9010)
);

INVxp67_ASAP7_75t_SL g9011 ( 
.A(n_8652),
.Y(n_9011)
);

AO21x1_ASAP7_75t_L g9012 ( 
.A1(n_8011),
.A2(n_7137),
.B(n_7115),
.Y(n_9012)
);

BUFx2_ASAP7_75t_L g9013 ( 
.A(n_8853),
.Y(n_9013)
);

CKINVDCx20_ASAP7_75t_R g9014 ( 
.A(n_7966),
.Y(n_9014)
);

OAI21x1_ASAP7_75t_SL g9015 ( 
.A1(n_7739),
.A2(n_7531),
.B(n_7460),
.Y(n_9015)
);

OR2x2_ASAP7_75t_L g9016 ( 
.A(n_8520),
.B(n_6735),
.Y(n_9016)
);

BUFx3_ASAP7_75t_L g9017 ( 
.A(n_8098),
.Y(n_9017)
);

AND2x2_ASAP7_75t_L g9018 ( 
.A(n_8586),
.B(n_6783),
.Y(n_9018)
);

INVx3_ASAP7_75t_L g9019 ( 
.A(n_8617),
.Y(n_9019)
);

INVx1_ASAP7_75t_L g9020 ( 
.A(n_8700),
.Y(n_9020)
);

AOI21x1_ASAP7_75t_L g9021 ( 
.A1(n_7708),
.A2(n_7542),
.B(n_7517),
.Y(n_9021)
);

NAND2xp5_ASAP7_75t_L g9022 ( 
.A(n_7734),
.B(n_7813),
.Y(n_9022)
);

INVx1_ASAP7_75t_L g9023 ( 
.A(n_8700),
.Y(n_9023)
);

AO21x2_ASAP7_75t_L g9024 ( 
.A1(n_8004),
.A2(n_7146),
.B(n_7115),
.Y(n_9024)
);

CKINVDCx6p67_ASAP7_75t_R g9025 ( 
.A(n_8022),
.Y(n_9025)
);

NAND2xp5_ASAP7_75t_L g9026 ( 
.A(n_7734),
.B(n_7116),
.Y(n_9026)
);

NAND2x1p5_ASAP7_75t_L g9027 ( 
.A(n_7686),
.B(n_7338),
.Y(n_9027)
);

HB1xp67_ASAP7_75t_L g9028 ( 
.A(n_8700),
.Y(n_9028)
);

AOI21xp5_ASAP7_75t_L g9029 ( 
.A1(n_7796),
.A2(n_7084),
.B(n_7023),
.Y(n_9029)
);

AOI22xp33_ASAP7_75t_L g9030 ( 
.A1(n_7809),
.A2(n_6683),
.B1(n_6558),
.B2(n_6970),
.Y(n_9030)
);

AOI21xp5_ASAP7_75t_L g9031 ( 
.A1(n_7796),
.A2(n_7201),
.B(n_7084),
.Y(n_9031)
);

OAI21xp5_ASAP7_75t_L g9032 ( 
.A1(n_7781),
.A2(n_7830),
.B(n_7773),
.Y(n_9032)
);

INVx1_ASAP7_75t_L g9033 ( 
.A(n_8711),
.Y(n_9033)
);

AOI21x1_ASAP7_75t_L g9034 ( 
.A1(n_7708),
.A2(n_7547),
.B(n_7542),
.Y(n_9034)
);

BUFx3_ASAP7_75t_L g9035 ( 
.A(n_8098),
.Y(n_9035)
);

NAND2xp5_ASAP7_75t_SL g9036 ( 
.A(n_7863),
.B(n_6388),
.Y(n_9036)
);

A2O1A1Ixp33_ASAP7_75t_L g9037 ( 
.A1(n_7716),
.A2(n_6411),
.B(n_7116),
.C(n_6683),
.Y(n_9037)
);

AOI21xp33_ASAP7_75t_L g9038 ( 
.A1(n_7889),
.A2(n_7160),
.B(n_7146),
.Y(n_9038)
);

INVx1_ASAP7_75t_L g9039 ( 
.A(n_8711),
.Y(n_9039)
);

INVx3_ASAP7_75t_L g9040 ( 
.A(n_8617),
.Y(n_9040)
);

INVx1_ASAP7_75t_L g9041 ( 
.A(n_8711),
.Y(n_9041)
);

INVx2_ASAP7_75t_L g9042 ( 
.A(n_7702),
.Y(n_9042)
);

INVx2_ASAP7_75t_L g9043 ( 
.A(n_7702),
.Y(n_9043)
);

BUFx3_ASAP7_75t_L g9044 ( 
.A(n_8158),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_8711),
.Y(n_9045)
);

AND2x2_ASAP7_75t_L g9046 ( 
.A(n_8586),
.B(n_7784),
.Y(n_9046)
);

AND2x4_ASAP7_75t_L g9047 ( 
.A(n_8867),
.B(n_7469),
.Y(n_9047)
);

AND2x4_ASAP7_75t_L g9048 ( 
.A(n_8867),
.B(n_7469),
.Y(n_9048)
);

AOI21xp5_ASAP7_75t_L g9049 ( 
.A1(n_7802),
.A2(n_7230),
.B(n_7201),
.Y(n_9049)
);

NOR2xp33_ASAP7_75t_L g9050 ( 
.A(n_7874),
.B(n_6902),
.Y(n_9050)
);

INVx4_ASAP7_75t_L g9051 ( 
.A(n_7971),
.Y(n_9051)
);

INVx2_ASAP7_75t_L g9052 ( 
.A(n_7702),
.Y(n_9052)
);

INVx1_ASAP7_75t_L g9053 ( 
.A(n_8711),
.Y(n_9053)
);

INVx3_ASAP7_75t_L g9054 ( 
.A(n_8617),
.Y(n_9054)
);

INVx1_ASAP7_75t_L g9055 ( 
.A(n_8711),
.Y(n_9055)
);

CKINVDCx5p33_ASAP7_75t_R g9056 ( 
.A(n_7966),
.Y(n_9056)
);

OAI21xp5_ASAP7_75t_L g9057 ( 
.A1(n_7781),
.A2(n_6481),
.B(n_6474),
.Y(n_9057)
);

OR3x4_ASAP7_75t_SL g9058 ( 
.A(n_8046),
.B(n_7675),
.C(n_6411),
.Y(n_9058)
);

NOR2x1_ASAP7_75t_R g9059 ( 
.A(n_8022),
.B(n_7460),
.Y(n_9059)
);

BUFx6f_ASAP7_75t_L g9060 ( 
.A(n_8549),
.Y(n_9060)
);

AOI22xp5_ASAP7_75t_L g9061 ( 
.A1(n_7908),
.A2(n_7553),
.B1(n_7573),
.B2(n_6756),
.Y(n_9061)
);

OAI21xp5_ASAP7_75t_L g9062 ( 
.A1(n_7830),
.A2(n_6481),
.B(n_7502),
.Y(n_9062)
);

NOR2x1_ASAP7_75t_R g9063 ( 
.A(n_8022),
.B(n_7460),
.Y(n_9063)
);

AOI22x1_ASAP7_75t_L g9064 ( 
.A1(n_7928),
.A2(n_7271),
.B1(n_7285),
.B2(n_7230),
.Y(n_9064)
);

NAND2x1p5_ASAP7_75t_L g9065 ( 
.A(n_7686),
.B(n_7714),
.Y(n_9065)
);

AND2x4_ASAP7_75t_L g9066 ( 
.A(n_8867),
.B(n_7715),
.Y(n_9066)
);

AO21x2_ASAP7_75t_L g9067 ( 
.A1(n_7778),
.A2(n_7186),
.B(n_7177),
.Y(n_9067)
);

BUFx3_ASAP7_75t_L g9068 ( 
.A(n_8158),
.Y(n_9068)
);

OAI21x1_ASAP7_75t_L g9069 ( 
.A1(n_8077),
.A2(n_8089),
.B(n_8097),
.Y(n_9069)
);

INVx1_ASAP7_75t_L g9070 ( 
.A(n_8711),
.Y(n_9070)
);

INVx2_ASAP7_75t_L g9071 ( 
.A(n_7702),
.Y(n_9071)
);

INVx3_ASAP7_75t_L g9072 ( 
.A(n_8617),
.Y(n_9072)
);

BUFx8_ASAP7_75t_L g9073 ( 
.A(n_8022),
.Y(n_9073)
);

NAND2x1_ASAP7_75t_L g9074 ( 
.A(n_8137),
.B(n_7588),
.Y(n_9074)
);

BUFx2_ASAP7_75t_L g9075 ( 
.A(n_8853),
.Y(n_9075)
);

AOI22xp33_ASAP7_75t_SL g9076 ( 
.A1(n_7805),
.A2(n_6756),
.B1(n_6411),
.B2(n_6683),
.Y(n_9076)
);

BUFx6f_ASAP7_75t_L g9077 ( 
.A(n_8549),
.Y(n_9077)
);

BUFx2_ASAP7_75t_L g9078 ( 
.A(n_8853),
.Y(n_9078)
);

OA21x2_ASAP7_75t_L g9079 ( 
.A1(n_8455),
.A2(n_7509),
.B(n_7506),
.Y(n_9079)
);

OAI21x1_ASAP7_75t_L g9080 ( 
.A1(n_8089),
.A2(n_8097),
.B(n_8144),
.Y(n_9080)
);

INVx1_ASAP7_75t_L g9081 ( 
.A(n_8711),
.Y(n_9081)
);

BUFx4f_ASAP7_75t_L g9082 ( 
.A(n_7971),
.Y(n_9082)
);

OAI21x1_ASAP7_75t_SL g9083 ( 
.A1(n_7739),
.A2(n_7531),
.B(n_7570),
.Y(n_9083)
);

INVx2_ASAP7_75t_SL g9084 ( 
.A(n_8867),
.Y(n_9084)
);

AOI22xp33_ASAP7_75t_L g9085 ( 
.A1(n_7805),
.A2(n_6683),
.B1(n_6558),
.B2(n_6970),
.Y(n_9085)
);

BUFx3_ASAP7_75t_L g9086 ( 
.A(n_8158),
.Y(n_9086)
);

BUFx2_ASAP7_75t_R g9087 ( 
.A(n_8090),
.Y(n_9087)
);

AOI21x1_ASAP7_75t_L g9088 ( 
.A1(n_7708),
.A2(n_8518),
.B(n_7913),
.Y(n_9088)
);

AND2x4_ASAP7_75t_L g9089 ( 
.A(n_8867),
.B(n_7469),
.Y(n_9089)
);

BUFx3_ASAP7_75t_L g9090 ( 
.A(n_8181),
.Y(n_9090)
);

BUFx2_ASAP7_75t_L g9091 ( 
.A(n_8853),
.Y(n_9091)
);

NAND2x1_ASAP7_75t_L g9092 ( 
.A(n_8149),
.B(n_7588),
.Y(n_9092)
);

BUFx2_ASAP7_75t_L g9093 ( 
.A(n_8853),
.Y(n_9093)
);

BUFx4f_ASAP7_75t_L g9094 ( 
.A(n_7971),
.Y(n_9094)
);

OAI21xp5_ASAP7_75t_L g9095 ( 
.A1(n_7773),
.A2(n_6481),
.B(n_7523),
.Y(n_9095)
);

INVx1_ASAP7_75t_L g9096 ( 
.A(n_8711),
.Y(n_9096)
);

BUFx3_ASAP7_75t_L g9097 ( 
.A(n_8181),
.Y(n_9097)
);

OR2x2_ASAP7_75t_L g9098 ( 
.A(n_8520),
.B(n_6735),
.Y(n_9098)
);

CKINVDCx6p67_ASAP7_75t_R g9099 ( 
.A(n_8025),
.Y(n_9099)
);

INVx1_ASAP7_75t_L g9100 ( 
.A(n_8713),
.Y(n_9100)
);

OA21x2_ASAP7_75t_L g9101 ( 
.A1(n_8455),
.A2(n_7529),
.B(n_7523),
.Y(n_9101)
);

INVx3_ASAP7_75t_L g9102 ( 
.A(n_8617),
.Y(n_9102)
);

INVx1_ASAP7_75t_L g9103 ( 
.A(n_8713),
.Y(n_9103)
);

AND2x2_ASAP7_75t_L g9104 ( 
.A(n_8586),
.B(n_6783),
.Y(n_9104)
);

AND2x2_ASAP7_75t_L g9105 ( 
.A(n_8586),
.B(n_6816),
.Y(n_9105)
);

AOI22xp33_ASAP7_75t_L g9106 ( 
.A1(n_7924),
.A2(n_6683),
.B1(n_6558),
.B2(n_6970),
.Y(n_9106)
);

INVx2_ASAP7_75t_L g9107 ( 
.A(n_7775),
.Y(n_9107)
);

INVx1_ASAP7_75t_SL g9108 ( 
.A(n_8642),
.Y(n_9108)
);

AND2x4_ASAP7_75t_L g9109 ( 
.A(n_8867),
.B(n_7489),
.Y(n_9109)
);

OA21x2_ASAP7_75t_L g9110 ( 
.A1(n_8455),
.A2(n_8539),
.B(n_7802),
.Y(n_9110)
);

NOR2xp33_ASAP7_75t_L g9111 ( 
.A(n_7799),
.B(n_6902),
.Y(n_9111)
);

AND2x2_ASAP7_75t_L g9112 ( 
.A(n_7784),
.B(n_6816),
.Y(n_9112)
);

AND2x4_ASAP7_75t_L g9113 ( 
.A(n_8867),
.B(n_7489),
.Y(n_9113)
);

INVx2_ASAP7_75t_L g9114 ( 
.A(n_7775),
.Y(n_9114)
);

OAI21xp5_ASAP7_75t_L g9115 ( 
.A1(n_7950),
.A2(n_7544),
.B(n_7540),
.Y(n_9115)
);

OAI21xp5_ASAP7_75t_L g9116 ( 
.A1(n_7950),
.A2(n_7544),
.B(n_7540),
.Y(n_9116)
);

OR2x2_ASAP7_75t_L g9117 ( 
.A(n_8520),
.B(n_8411),
.Y(n_9117)
);

NAND2xp5_ASAP7_75t_L g9118 ( 
.A(n_7813),
.B(n_7116),
.Y(n_9118)
);

A2O1A1Ixp33_ASAP7_75t_L g9119 ( 
.A1(n_7716),
.A2(n_7712),
.B(n_7806),
.C(n_7882),
.Y(n_9119)
);

INVx2_ASAP7_75t_L g9120 ( 
.A(n_7775),
.Y(n_9120)
);

AND2x2_ASAP7_75t_L g9121 ( 
.A(n_7784),
.B(n_6816),
.Y(n_9121)
);

NAND2xp5_ASAP7_75t_L g9122 ( 
.A(n_7725),
.B(n_7116),
.Y(n_9122)
);

OA21x2_ASAP7_75t_L g9123 ( 
.A1(n_8539),
.A2(n_7544),
.B(n_7540),
.Y(n_9123)
);

AOI21xp33_ASAP7_75t_L g9124 ( 
.A1(n_7889),
.A2(n_7251),
.B(n_7227),
.Y(n_9124)
);

BUFx3_ASAP7_75t_L g9125 ( 
.A(n_8181),
.Y(n_9125)
);

AND2x2_ASAP7_75t_L g9126 ( 
.A(n_7784),
.B(n_6860),
.Y(n_9126)
);

AOI22xp33_ASAP7_75t_L g9127 ( 
.A1(n_7924),
.A2(n_6558),
.B1(n_6970),
.B2(n_7630),
.Y(n_9127)
);

INVx1_ASAP7_75t_L g9128 ( 
.A(n_8713),
.Y(n_9128)
);

AND2x4_ASAP7_75t_L g9129 ( 
.A(n_8867),
.B(n_7489),
.Y(n_9129)
);

AOI21x1_ASAP7_75t_L g9130 ( 
.A1(n_8518),
.A2(n_7551),
.B(n_7547),
.Y(n_9130)
);

BUFx8_ASAP7_75t_L g9131 ( 
.A(n_8025),
.Y(n_9131)
);

INVx1_ASAP7_75t_L g9132 ( 
.A(n_8713),
.Y(n_9132)
);

INVx1_ASAP7_75t_L g9133 ( 
.A(n_8713),
.Y(n_9133)
);

BUFx2_ASAP7_75t_R g9134 ( 
.A(n_8090),
.Y(n_9134)
);

OAI21x1_ASAP7_75t_L g9135 ( 
.A1(n_8150),
.A2(n_8372),
.B(n_8333),
.Y(n_9135)
);

OAI21x1_ASAP7_75t_L g9136 ( 
.A1(n_8150),
.A2(n_8372),
.B(n_8333),
.Y(n_9136)
);

NOR2xp33_ASAP7_75t_L g9137 ( 
.A(n_7799),
.B(n_7927),
.Y(n_9137)
);

INVx2_ASAP7_75t_L g9138 ( 
.A(n_7775),
.Y(n_9138)
);

NAND3xp33_ASAP7_75t_L g9139 ( 
.A(n_7789),
.B(n_7257),
.C(n_7255),
.Y(n_9139)
);

OAI21xp5_ASAP7_75t_L g9140 ( 
.A1(n_7961),
.A2(n_7618),
.B(n_7615),
.Y(n_9140)
);

BUFx6f_ASAP7_75t_L g9141 ( 
.A(n_8549),
.Y(n_9141)
);

NAND2xp5_ASAP7_75t_L g9142 ( 
.A(n_7725),
.B(n_7116),
.Y(n_9142)
);

CKINVDCx11_ASAP7_75t_R g9143 ( 
.A(n_8025),
.Y(n_9143)
);

HB1xp67_ASAP7_75t_L g9144 ( 
.A(n_8713),
.Y(n_9144)
);

AOI22x1_ASAP7_75t_L g9145 ( 
.A1(n_7928),
.A2(n_7271),
.B1(n_7285),
.B2(n_7230),
.Y(n_9145)
);

AND2x4_ASAP7_75t_L g9146 ( 
.A(n_7715),
.B(n_7489),
.Y(n_9146)
);

INVx1_ASAP7_75t_L g9147 ( 
.A(n_8713),
.Y(n_9147)
);

BUFx12f_ASAP7_75t_L g9148 ( 
.A(n_8025),
.Y(n_9148)
);

CKINVDCx20_ASAP7_75t_R g9149 ( 
.A(n_7974),
.Y(n_9149)
);

NAND2xp5_ASAP7_75t_L g9150 ( 
.A(n_7743),
.B(n_7116),
.Y(n_9150)
);

INVx2_ASAP7_75t_L g9151 ( 
.A(n_7787),
.Y(n_9151)
);

AOI22xp33_ASAP7_75t_L g9152 ( 
.A1(n_7712),
.A2(n_6558),
.B1(n_6970),
.B2(n_7630),
.Y(n_9152)
);

AND2x2_ASAP7_75t_L g9153 ( 
.A(n_7793),
.B(n_6860),
.Y(n_9153)
);

AOI21x1_ASAP7_75t_L g9154 ( 
.A1(n_8518),
.A2(n_7572),
.B(n_7551),
.Y(n_9154)
);

INVx1_ASAP7_75t_L g9155 ( 
.A(n_8713),
.Y(n_9155)
);

NAND2x1p5_ASAP7_75t_L g9156 ( 
.A(n_7686),
.B(n_7714),
.Y(n_9156)
);

NAND2xp5_ASAP7_75t_L g9157 ( 
.A(n_7743),
.B(n_7116),
.Y(n_9157)
);

BUFx3_ASAP7_75t_L g9158 ( 
.A(n_7881),
.Y(n_9158)
);

NOR2xp67_ASAP7_75t_L g9159 ( 
.A(n_7686),
.B(n_7380),
.Y(n_9159)
);

INVx2_ASAP7_75t_L g9160 ( 
.A(n_7787),
.Y(n_9160)
);

BUFx12f_ASAP7_75t_L g9161 ( 
.A(n_8059),
.Y(n_9161)
);

INVx1_ASAP7_75t_L g9162 ( 
.A(n_8713),
.Y(n_9162)
);

AND2x2_ASAP7_75t_L g9163 ( 
.A(n_7793),
.B(n_6860),
.Y(n_9163)
);

AND2x2_ASAP7_75t_L g9164 ( 
.A(n_7793),
.B(n_6860),
.Y(n_9164)
);

INVx1_ASAP7_75t_L g9165 ( 
.A(n_8763),
.Y(n_9165)
);

INVx2_ASAP7_75t_L g9166 ( 
.A(n_7787),
.Y(n_9166)
);

BUFx3_ASAP7_75t_L g9167 ( 
.A(n_7881),
.Y(n_9167)
);

NOR2xp33_ASAP7_75t_L g9168 ( 
.A(n_7799),
.B(n_6902),
.Y(n_9168)
);

BUFx3_ASAP7_75t_L g9169 ( 
.A(n_7881),
.Y(n_9169)
);

INVx2_ASAP7_75t_L g9170 ( 
.A(n_7787),
.Y(n_9170)
);

AND2x2_ASAP7_75t_L g9171 ( 
.A(n_7793),
.B(n_7848),
.Y(n_9171)
);

INVx3_ASAP7_75t_L g9172 ( 
.A(n_8617),
.Y(n_9172)
);

INVx1_ASAP7_75t_L g9173 ( 
.A(n_8763),
.Y(n_9173)
);

NAND2x1_ASAP7_75t_L g9174 ( 
.A(n_8149),
.B(n_7588),
.Y(n_9174)
);

BUFx10_ASAP7_75t_L g9175 ( 
.A(n_8105),
.Y(n_9175)
);

INVx1_ASAP7_75t_L g9176 ( 
.A(n_8763),
.Y(n_9176)
);

NAND2xp5_ASAP7_75t_SL g9177 ( 
.A(n_7863),
.B(n_6388),
.Y(n_9177)
);

INVx3_ASAP7_75t_SL g9178 ( 
.A(n_8069),
.Y(n_9178)
);

NOR2xp33_ASAP7_75t_L g9179 ( 
.A(n_7927),
.B(n_6902),
.Y(n_9179)
);

NAND3xp33_ASAP7_75t_L g9180 ( 
.A(n_7789),
.B(n_7257),
.C(n_7255),
.Y(n_9180)
);

HB1xp67_ASAP7_75t_L g9181 ( 
.A(n_8763),
.Y(n_9181)
);

AND2x4_ASAP7_75t_L g9182 ( 
.A(n_7715),
.B(n_7489),
.Y(n_9182)
);

AND2x4_ASAP7_75t_L g9183 ( 
.A(n_7715),
.B(n_7489),
.Y(n_9183)
);

NOR2xp33_ASAP7_75t_L g9184 ( 
.A(n_7927),
.B(n_6941),
.Y(n_9184)
);

BUFx12f_ASAP7_75t_L g9185 ( 
.A(n_8059),
.Y(n_9185)
);

INVx3_ASAP7_75t_L g9186 ( 
.A(n_7815),
.Y(n_9186)
);

OAI21xp5_ASAP7_75t_L g9187 ( 
.A1(n_7961),
.A2(n_7618),
.B(n_7316),
.Y(n_9187)
);

OAI21x1_ASAP7_75t_L g9188 ( 
.A1(n_8343),
.A2(n_8003),
.B(n_8360),
.Y(n_9188)
);

BUFx2_ASAP7_75t_L g9189 ( 
.A(n_8853),
.Y(n_9189)
);

OR2x2_ASAP7_75t_L g9190 ( 
.A(n_8411),
.B(n_7986),
.Y(n_9190)
);

NAND2xp5_ASAP7_75t_L g9191 ( 
.A(n_7767),
.B(n_6262),
.Y(n_9191)
);

NAND2xp5_ASAP7_75t_L g9192 ( 
.A(n_7767),
.B(n_6262),
.Y(n_9192)
);

INVx1_ASAP7_75t_L g9193 ( 
.A(n_8763),
.Y(n_9193)
);

INVx1_ASAP7_75t_L g9194 ( 
.A(n_8763),
.Y(n_9194)
);

HB1xp67_ASAP7_75t_L g9195 ( 
.A(n_8763),
.Y(n_9195)
);

NAND3xp33_ASAP7_75t_L g9196 ( 
.A(n_7758),
.B(n_7281),
.C(n_7261),
.Y(n_9196)
);

INVx1_ASAP7_75t_L g9197 ( 
.A(n_8763),
.Y(n_9197)
);

AND2x4_ASAP7_75t_L g9198 ( 
.A(n_7815),
.B(n_7489),
.Y(n_9198)
);

AOI22x1_ASAP7_75t_L g9199 ( 
.A1(n_7933),
.A2(n_7347),
.B1(n_7338),
.B2(n_7531),
.Y(n_9199)
);

INVxp67_ASAP7_75t_L g9200 ( 
.A(n_8328),
.Y(n_9200)
);

CKINVDCx16_ASAP7_75t_R g9201 ( 
.A(n_8125),
.Y(n_9201)
);

AOI22xp5_ASAP7_75t_L g9202 ( 
.A1(n_7908),
.A2(n_7573),
.B1(n_7553),
.B2(n_6338),
.Y(n_9202)
);

OAI21x1_ASAP7_75t_L g9203 ( 
.A1(n_8360),
.A2(n_8355),
.B(n_7780),
.Y(n_9203)
);

BUFx3_ASAP7_75t_L g9204 ( 
.A(n_7912),
.Y(n_9204)
);

AO31x2_ASAP7_75t_L g9205 ( 
.A1(n_7777),
.A2(n_7294),
.A3(n_7290),
.B(n_7281),
.Y(n_9205)
);

NOR2xp33_ASAP7_75t_L g9206 ( 
.A(n_7934),
.B(n_7726),
.Y(n_9206)
);

INVx1_ASAP7_75t_L g9207 ( 
.A(n_8763),
.Y(n_9207)
);

CKINVDCx8_ASAP7_75t_R g9208 ( 
.A(n_8105),
.Y(n_9208)
);

AND2x2_ASAP7_75t_L g9209 ( 
.A(n_7848),
.B(n_6864),
.Y(n_9209)
);

INVx4_ASAP7_75t_L g9210 ( 
.A(n_7971),
.Y(n_9210)
);

NOR2xp67_ASAP7_75t_L g9211 ( 
.A(n_7686),
.B(n_7380),
.Y(n_9211)
);

OR3x4_ASAP7_75t_SL g9212 ( 
.A(n_8046),
.B(n_7675),
.C(n_6411),
.Y(n_9212)
);

OAI21x1_ASAP7_75t_L g9213 ( 
.A1(n_8360),
.A2(n_8355),
.B(n_7780),
.Y(n_9213)
);

INVx3_ASAP7_75t_L g9214 ( 
.A(n_7815),
.Y(n_9214)
);

INVx1_ASAP7_75t_L g9215 ( 
.A(n_8819),
.Y(n_9215)
);

INVx1_ASAP7_75t_L g9216 ( 
.A(n_8819),
.Y(n_9216)
);

AND2x4_ASAP7_75t_L g9217 ( 
.A(n_7815),
.B(n_7489),
.Y(n_9217)
);

NAND2xp5_ASAP7_75t_L g9218 ( 
.A(n_7769),
.B(n_6262),
.Y(n_9218)
);

CKINVDCx5p33_ASAP7_75t_R g9219 ( 
.A(n_7929),
.Y(n_9219)
);

NAND2xp5_ASAP7_75t_SL g9220 ( 
.A(n_7846),
.B(n_6388),
.Y(n_9220)
);

INVx1_ASAP7_75t_L g9221 ( 
.A(n_8819),
.Y(n_9221)
);

AND2x4_ASAP7_75t_L g9222 ( 
.A(n_7821),
.B(n_7489),
.Y(n_9222)
);

OAI21xp5_ASAP7_75t_L g9223 ( 
.A1(n_7824),
.A2(n_7618),
.B(n_7325),
.Y(n_9223)
);

AND2x2_ASAP7_75t_L g9224 ( 
.A(n_7848),
.B(n_6864),
.Y(n_9224)
);

CKINVDCx20_ASAP7_75t_R g9225 ( 
.A(n_7974),
.Y(n_9225)
);

OAI21x1_ASAP7_75t_L g9226 ( 
.A1(n_7780),
.A2(n_7938),
.B(n_7936),
.Y(n_9226)
);

INVx1_ASAP7_75t_L g9227 ( 
.A(n_8819),
.Y(n_9227)
);

OAI21xp5_ASAP7_75t_L g9228 ( 
.A1(n_7824),
.A2(n_7618),
.B(n_7335),
.Y(n_9228)
);

INVx5_ASAP7_75t_L g9229 ( 
.A(n_8549),
.Y(n_9229)
);

OR2x2_ASAP7_75t_L g9230 ( 
.A(n_8411),
.B(n_6735),
.Y(n_9230)
);

OR2x2_ASAP7_75t_L g9231 ( 
.A(n_8411),
.B(n_6735),
.Y(n_9231)
);

NOR2xp33_ASAP7_75t_L g9232 ( 
.A(n_7934),
.B(n_6941),
.Y(n_9232)
);

OAI21x1_ASAP7_75t_SL g9233 ( 
.A1(n_7739),
.A2(n_7753),
.B(n_7817),
.Y(n_9233)
);

INVx1_ASAP7_75t_L g9234 ( 
.A(n_8819),
.Y(n_9234)
);

INVx1_ASAP7_75t_L g9235 ( 
.A(n_8819),
.Y(n_9235)
);

CKINVDCx5p33_ASAP7_75t_R g9236 ( 
.A(n_7929),
.Y(n_9236)
);

BUFx3_ASAP7_75t_L g9237 ( 
.A(n_7912),
.Y(n_9237)
);

INVx1_ASAP7_75t_L g9238 ( 
.A(n_8819),
.Y(n_9238)
);

AO21x2_ASAP7_75t_L g9239 ( 
.A1(n_7973),
.A2(n_7294),
.B(n_7284),
.Y(n_9239)
);

INVx4_ASAP7_75t_L g9240 ( 
.A(n_7971),
.Y(n_9240)
);

AND2x4_ASAP7_75t_L g9241 ( 
.A(n_7821),
.B(n_7590),
.Y(n_9241)
);

AOI22xp33_ASAP7_75t_L g9242 ( 
.A1(n_7758),
.A2(n_7649),
.B1(n_7630),
.B2(n_7531),
.Y(n_9242)
);

INVx4_ASAP7_75t_L g9243 ( 
.A(n_7971),
.Y(n_9243)
);

OR2x2_ASAP7_75t_L g9244 ( 
.A(n_8411),
.B(n_6735),
.Y(n_9244)
);

INVx3_ASAP7_75t_L g9245 ( 
.A(n_7821),
.Y(n_9245)
);

A2O1A1Ixp33_ASAP7_75t_SL g9246 ( 
.A1(n_7933),
.A2(n_7670),
.B(n_7539),
.C(n_7497),
.Y(n_9246)
);

OAI21x1_ASAP7_75t_SL g9247 ( 
.A1(n_7753),
.A2(n_7593),
.B(n_7578),
.Y(n_9247)
);

NOR2xp33_ASAP7_75t_SL g9248 ( 
.A(n_8023),
.B(n_7338),
.Y(n_9248)
);

NAND2x1_ASAP7_75t_L g9249 ( 
.A(n_8149),
.B(n_8345),
.Y(n_9249)
);

AOI21xp5_ASAP7_75t_L g9250 ( 
.A1(n_7828),
.A2(n_6556),
.B(n_6516),
.Y(n_9250)
);

AND2x6_ASAP7_75t_L g9251 ( 
.A(n_7752),
.B(n_7630),
.Y(n_9251)
);

HB1xp67_ASAP7_75t_L g9252 ( 
.A(n_8819),
.Y(n_9252)
);

AOI21xp5_ASAP7_75t_L g9253 ( 
.A1(n_7828),
.A2(n_6556),
.B(n_6516),
.Y(n_9253)
);

NAND3xp33_ASAP7_75t_L g9254 ( 
.A(n_7968),
.B(n_7294),
.C(n_7578),
.Y(n_9254)
);

CKINVDCx8_ASAP7_75t_R g9255 ( 
.A(n_8105),
.Y(n_9255)
);

BUFx3_ASAP7_75t_L g9256 ( 
.A(n_7912),
.Y(n_9256)
);

INVx1_ASAP7_75t_L g9257 ( 
.A(n_8819),
.Y(n_9257)
);

NAND3xp33_ASAP7_75t_L g9258 ( 
.A(n_7968),
.B(n_7597),
.C(n_7593),
.Y(n_9258)
);

OAI21xp5_ASAP7_75t_L g9259 ( 
.A1(n_7885),
.A2(n_7358),
.B(n_7572),
.Y(n_9259)
);

AOI22xp33_ASAP7_75t_L g9260 ( 
.A1(n_7726),
.A2(n_7649),
.B1(n_7630),
.B2(n_7588),
.Y(n_9260)
);

NAND2x1p5_ASAP7_75t_L g9261 ( 
.A(n_7686),
.B(n_7714),
.Y(n_9261)
);

OAI221xp5_ASAP7_75t_SL g9262 ( 
.A1(n_7841),
.A2(n_6262),
.B1(n_7588),
.B2(n_7626),
.C(n_6272),
.Y(n_9262)
);

AOI21xp5_ASAP7_75t_L g9263 ( 
.A1(n_7973),
.A2(n_6556),
.B(n_6516),
.Y(n_9263)
);

AND2x2_ASAP7_75t_L g9264 ( 
.A(n_7848),
.B(n_6864),
.Y(n_9264)
);

AND2x4_ASAP7_75t_L g9265 ( 
.A(n_7821),
.B(n_7590),
.Y(n_9265)
);

NAND2x1p5_ASAP7_75t_L g9266 ( 
.A(n_7686),
.B(n_7714),
.Y(n_9266)
);

BUFx3_ASAP7_75t_L g9267 ( 
.A(n_8008),
.Y(n_9267)
);

AO21x2_ASAP7_75t_L g9268 ( 
.A1(n_8102),
.A2(n_7597),
.B(n_7593),
.Y(n_9268)
);

CKINVDCx5p33_ASAP7_75t_R g9269 ( 
.A(n_7962),
.Y(n_9269)
);

INVx2_ASAP7_75t_L g9270 ( 
.A(n_7814),
.Y(n_9270)
);

INVx3_ASAP7_75t_L g9271 ( 
.A(n_7886),
.Y(n_9271)
);

BUFx2_ASAP7_75t_SL g9272 ( 
.A(n_7847),
.Y(n_9272)
);

AOI21x1_ASAP7_75t_L g9273 ( 
.A1(n_7913),
.A2(n_7610),
.B(n_7588),
.Y(n_9273)
);

INVx2_ASAP7_75t_L g9274 ( 
.A(n_7814),
.Y(n_9274)
);

HB1xp67_ASAP7_75t_L g9275 ( 
.A(n_8870),
.Y(n_9275)
);

INVx1_ASAP7_75t_L g9276 ( 
.A(n_8870),
.Y(n_9276)
);

AOI22xp5_ASAP7_75t_L g9277 ( 
.A1(n_7747),
.A2(n_7882),
.B1(n_7770),
.B2(n_7806),
.Y(n_9277)
);

INVx2_ASAP7_75t_L g9278 ( 
.A(n_7814),
.Y(n_9278)
);

NAND2xp5_ASAP7_75t_L g9279 ( 
.A(n_7769),
.B(n_6262),
.Y(n_9279)
);

NAND2xp5_ASAP7_75t_L g9280 ( 
.A(n_7783),
.B(n_6262),
.Y(n_9280)
);

INVx1_ASAP7_75t_L g9281 ( 
.A(n_8870),
.Y(n_9281)
);

INVx3_ASAP7_75t_L g9282 ( 
.A(n_7886),
.Y(n_9282)
);

OA21x2_ASAP7_75t_L g9283 ( 
.A1(n_7819),
.A2(n_8655),
.B(n_7964),
.Y(n_9283)
);

INVx1_ASAP7_75t_L g9284 ( 
.A(n_8870),
.Y(n_9284)
);

AOI22xp33_ASAP7_75t_L g9285 ( 
.A1(n_7747),
.A2(n_7649),
.B1(n_7630),
.B2(n_7588),
.Y(n_9285)
);

INVx1_ASAP7_75t_L g9286 ( 
.A(n_8870),
.Y(n_9286)
);

CKINVDCx6p67_ASAP7_75t_R g9287 ( 
.A(n_8059),
.Y(n_9287)
);

AO21x2_ASAP7_75t_L g9288 ( 
.A1(n_8102),
.A2(n_6750),
.B(n_6716),
.Y(n_9288)
);

NAND2x1p5_ASAP7_75t_L g9289 ( 
.A(n_7686),
.B(n_7347),
.Y(n_9289)
);

HB1xp67_ASAP7_75t_L g9290 ( 
.A(n_8870),
.Y(n_9290)
);

NAND2xp5_ASAP7_75t_L g9291 ( 
.A(n_7783),
.B(n_6262),
.Y(n_9291)
);

INVx1_ASAP7_75t_L g9292 ( 
.A(n_8870),
.Y(n_9292)
);

NAND2x1p5_ASAP7_75t_L g9293 ( 
.A(n_7686),
.B(n_6516),
.Y(n_9293)
);

INVx1_ASAP7_75t_SL g9294 ( 
.A(n_8642),
.Y(n_9294)
);

BUFx2_ASAP7_75t_L g9295 ( 
.A(n_8853),
.Y(n_9295)
);

BUFx2_ASAP7_75t_SL g9296 ( 
.A(n_7847),
.Y(n_9296)
);

BUFx3_ASAP7_75t_L g9297 ( 
.A(n_8008),
.Y(n_9297)
);

NAND2xp5_ASAP7_75t_L g9298 ( 
.A(n_8351),
.B(n_6262),
.Y(n_9298)
);

INVx2_ASAP7_75t_L g9299 ( 
.A(n_7814),
.Y(n_9299)
);

NAND2x1p5_ASAP7_75t_L g9300 ( 
.A(n_7714),
.B(n_6516),
.Y(n_9300)
);

INVx3_ASAP7_75t_L g9301 ( 
.A(n_7886),
.Y(n_9301)
);

INVx2_ASAP7_75t_L g9302 ( 
.A(n_8566),
.Y(n_9302)
);

INVx1_ASAP7_75t_L g9303 ( 
.A(n_8870),
.Y(n_9303)
);

OAI21x1_ASAP7_75t_SL g9304 ( 
.A1(n_7753),
.A2(n_7528),
.B(n_7526),
.Y(n_9304)
);

INVx1_ASAP7_75t_L g9305 ( 
.A(n_8870),
.Y(n_9305)
);

INVx1_ASAP7_75t_L g9306 ( 
.A(n_8903),
.Y(n_9306)
);

INVx1_ASAP7_75t_L g9307 ( 
.A(n_8903),
.Y(n_9307)
);

OR2x2_ASAP7_75t_L g9308 ( 
.A(n_8411),
.B(n_6735),
.Y(n_9308)
);

INVx1_ASAP7_75t_L g9309 ( 
.A(n_8903),
.Y(n_9309)
);

AO21x2_ASAP7_75t_L g9310 ( 
.A1(n_8106),
.A2(n_6765),
.B(n_6759),
.Y(n_9310)
);

AND2x4_ASAP7_75t_L g9311 ( 
.A(n_7886),
.B(n_7590),
.Y(n_9311)
);

AND2x4_ASAP7_75t_L g9312 ( 
.A(n_8132),
.B(n_7590),
.Y(n_9312)
);

INVx1_ASAP7_75t_L g9313 ( 
.A(n_8903),
.Y(n_9313)
);

AO21x2_ASAP7_75t_L g9314 ( 
.A1(n_8106),
.A2(n_6765),
.B(n_6759),
.Y(n_9314)
);

HB1xp67_ASAP7_75t_L g9315 ( 
.A(n_8903),
.Y(n_9315)
);

INVx2_ASAP7_75t_L g9316 ( 
.A(n_8566),
.Y(n_9316)
);

INVx1_ASAP7_75t_L g9317 ( 
.A(n_8903),
.Y(n_9317)
);

OAI21x1_ASAP7_75t_L g9318 ( 
.A1(n_8406),
.A2(n_8610),
.B(n_8601),
.Y(n_9318)
);

AO21x1_ASAP7_75t_L g9319 ( 
.A1(n_8091),
.A2(n_7528),
.B(n_7526),
.Y(n_9319)
);

AND2x2_ASAP7_75t_L g9320 ( 
.A(n_7892),
.B(n_7774),
.Y(n_9320)
);

AOI22x1_ASAP7_75t_L g9321 ( 
.A1(n_7811),
.A2(n_6828),
.B1(n_6776),
.B2(n_6731),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_8903),
.Y(n_9322)
);

OA21x2_ASAP7_75t_L g9323 ( 
.A1(n_8655),
.A2(n_6769),
.B(n_6765),
.Y(n_9323)
);

INVx1_ASAP7_75t_L g9324 ( 
.A(n_8903),
.Y(n_9324)
);

AOI22xp33_ASAP7_75t_SL g9325 ( 
.A1(n_7843),
.A2(n_6960),
.B1(n_6677),
.B2(n_7453),
.Y(n_9325)
);

AND2x4_ASAP7_75t_L g9326 ( 
.A(n_8132),
.B(n_7590),
.Y(n_9326)
);

OAI33xp33_ASAP7_75t_L g9327 ( 
.A1(n_7879),
.A2(n_7557),
.A3(n_7554),
.B1(n_7552),
.B2(n_7546),
.B3(n_7543),
.Y(n_9327)
);

BUFx12f_ASAP7_75t_L g9328 ( 
.A(n_8059),
.Y(n_9328)
);

INVx1_ASAP7_75t_SL g9329 ( 
.A(n_8642),
.Y(n_9329)
);

INVxp67_ASAP7_75t_L g9330 ( 
.A(n_8328),
.Y(n_9330)
);

NAND2xp5_ASAP7_75t_L g9331 ( 
.A(n_8351),
.B(n_6262),
.Y(n_9331)
);

INVx1_ASAP7_75t_SL g9332 ( 
.A(n_8642),
.Y(n_9332)
);

OR2x6_ASAP7_75t_L g9333 ( 
.A(n_8514),
.B(n_7588),
.Y(n_9333)
);

AOI21xp5_ASAP7_75t_L g9334 ( 
.A1(n_8005),
.A2(n_6556),
.B(n_6516),
.Y(n_9334)
);

NAND2x1_ASAP7_75t_L g9335 ( 
.A(n_8345),
.B(n_8346),
.Y(n_9335)
);

OA21x2_ASAP7_75t_L g9336 ( 
.A1(n_8655),
.A2(n_6775),
.B(n_6769),
.Y(n_9336)
);

OA21x2_ASAP7_75t_L g9337 ( 
.A1(n_8655),
.A2(n_6775),
.B(n_6769),
.Y(n_9337)
);

INVx1_ASAP7_75t_L g9338 ( 
.A(n_8903),
.Y(n_9338)
);

NAND2x1p5_ASAP7_75t_L g9339 ( 
.A(n_7714),
.B(n_6556),
.Y(n_9339)
);

INVx1_ASAP7_75t_L g9340 ( 
.A(n_8913),
.Y(n_9340)
);

NAND2xp5_ASAP7_75t_L g9341 ( 
.A(n_8354),
.B(n_6272),
.Y(n_9341)
);

INVx1_ASAP7_75t_L g9342 ( 
.A(n_8913),
.Y(n_9342)
);

AND2x2_ASAP7_75t_L g9343 ( 
.A(n_7892),
.B(n_6864),
.Y(n_9343)
);

AOI21xp5_ASAP7_75t_L g9344 ( 
.A1(n_8005),
.A2(n_6640),
.B(n_6556),
.Y(n_9344)
);

INVx3_ASAP7_75t_L g9345 ( 
.A(n_8132),
.Y(n_9345)
);

BUFx2_ASAP7_75t_L g9346 ( 
.A(n_8524),
.Y(n_9346)
);

OAI21x1_ASAP7_75t_SL g9347 ( 
.A1(n_7817),
.A2(n_7543),
.B(n_7537),
.Y(n_9347)
);

INVx2_ASAP7_75t_L g9348 ( 
.A(n_8566),
.Y(n_9348)
);

OAI22xp5_ASAP7_75t_L g9349 ( 
.A1(n_7816),
.A2(n_7569),
.B1(n_7549),
.B2(n_7649),
.Y(n_9349)
);

BUFx3_ASAP7_75t_L g9350 ( 
.A(n_8008),
.Y(n_9350)
);

NOR2xp67_ASAP7_75t_L g9351 ( 
.A(n_7714),
.B(n_7810),
.Y(n_9351)
);

INVx1_ASAP7_75t_L g9352 ( 
.A(n_8913),
.Y(n_9352)
);

CKINVDCx5p33_ASAP7_75t_R g9353 ( 
.A(n_7962),
.Y(n_9353)
);

INVx4_ASAP7_75t_L g9354 ( 
.A(n_7971),
.Y(n_9354)
);

INVx2_ASAP7_75t_L g9355 ( 
.A(n_8566),
.Y(n_9355)
);

INVx2_ASAP7_75t_L g9356 ( 
.A(n_8566),
.Y(n_9356)
);

INVx1_ASAP7_75t_L g9357 ( 
.A(n_8913),
.Y(n_9357)
);

NAND2x1p5_ASAP7_75t_L g9358 ( 
.A(n_7714),
.B(n_6556),
.Y(n_9358)
);

NAND2xp5_ASAP7_75t_L g9359 ( 
.A(n_8354),
.B(n_6272),
.Y(n_9359)
);

INVx1_ASAP7_75t_L g9360 ( 
.A(n_8913),
.Y(n_9360)
);

BUFx6f_ASAP7_75t_L g9361 ( 
.A(n_8549),
.Y(n_9361)
);

OAI21xp5_ASAP7_75t_L g9362 ( 
.A1(n_7885),
.A2(n_7626),
.B(n_7546),
.Y(n_9362)
);

INVx1_ASAP7_75t_L g9363 ( 
.A(n_8913),
.Y(n_9363)
);

AND2x2_ASAP7_75t_L g9364 ( 
.A(n_7892),
.B(n_6941),
.Y(n_9364)
);

O2A1O1Ixp33_ASAP7_75t_L g9365 ( 
.A1(n_7768),
.A2(n_7626),
.B(n_7537),
.C(n_7557),
.Y(n_9365)
);

INVx2_ASAP7_75t_L g9366 ( 
.A(n_8566),
.Y(n_9366)
);

BUFx4f_ASAP7_75t_SL g9367 ( 
.A(n_8254),
.Y(n_9367)
);

OAI21x1_ASAP7_75t_SL g9368 ( 
.A1(n_7817),
.A2(n_7554),
.B(n_7552),
.Y(n_9368)
);

INVxp33_ASAP7_75t_L g9369 ( 
.A(n_7889),
.Y(n_9369)
);

OA21x2_ASAP7_75t_L g9370 ( 
.A1(n_7856),
.A2(n_8414),
.B(n_8393),
.Y(n_9370)
);

INVx1_ASAP7_75t_L g9371 ( 
.A(n_8913),
.Y(n_9371)
);

OAI21xp5_ASAP7_75t_L g9372 ( 
.A1(n_7846),
.A2(n_7626),
.B(n_7029),
.Y(n_9372)
);

OAI21x1_ASAP7_75t_L g9373 ( 
.A1(n_7905),
.A2(n_7906),
.B(n_7926),
.Y(n_9373)
);

NOR2xp33_ASAP7_75t_L g9374 ( 
.A(n_7923),
.B(n_6941),
.Y(n_9374)
);

INVx1_ASAP7_75t_L g9375 ( 
.A(n_8913),
.Y(n_9375)
);

AND2x2_ASAP7_75t_L g9376 ( 
.A(n_7892),
.B(n_6994),
.Y(n_9376)
);

OR2x6_ASAP7_75t_L g9377 ( 
.A(n_8533),
.B(n_7626),
.Y(n_9377)
);

NAND2x1p5_ASAP7_75t_L g9378 ( 
.A(n_7714),
.B(n_6556),
.Y(n_9378)
);

AOI21xp5_ASAP7_75t_L g9379 ( 
.A1(n_7887),
.A2(n_6960),
.B(n_6731),
.Y(n_9379)
);

AOI21xp5_ASAP7_75t_L g9380 ( 
.A1(n_7887),
.A2(n_6960),
.B(n_6731),
.Y(n_9380)
);

BUFx3_ASAP7_75t_L g9381 ( 
.A(n_8159),
.Y(n_9381)
);

BUFx3_ASAP7_75t_L g9382 ( 
.A(n_8159),
.Y(n_9382)
);

INVx1_ASAP7_75t_L g9383 ( 
.A(n_8913),
.Y(n_9383)
);

NOR2xp33_ASAP7_75t_L g9384 ( 
.A(n_7923),
.B(n_6994),
.Y(n_9384)
);

AO21x2_ASAP7_75t_L g9385 ( 
.A1(n_7958),
.A2(n_7967),
.B(n_8110),
.Y(n_9385)
);

NOR2xp67_ASAP7_75t_L g9386 ( 
.A(n_7714),
.B(n_7670),
.Y(n_9386)
);

INVx1_ASAP7_75t_SL g9387 ( 
.A(n_8642),
.Y(n_9387)
);

BUFx12f_ASAP7_75t_L g9388 ( 
.A(n_8645),
.Y(n_9388)
);

NOR2xp33_ASAP7_75t_L g9389 ( 
.A(n_7947),
.B(n_6994),
.Y(n_9389)
);

BUFx3_ASAP7_75t_L g9390 ( 
.A(n_8159),
.Y(n_9390)
);

BUFx6f_ASAP7_75t_L g9391 ( 
.A(n_8549),
.Y(n_9391)
);

CKINVDCx16_ASAP7_75t_R g9392 ( 
.A(n_8125),
.Y(n_9392)
);

AND2x2_ASAP7_75t_L g9393 ( 
.A(n_7774),
.B(n_6994),
.Y(n_9393)
);

NAND2xp5_ASAP7_75t_L g9394 ( 
.A(n_8356),
.B(n_6272),
.Y(n_9394)
);

NOR2xp33_ASAP7_75t_L g9395 ( 
.A(n_7947),
.B(n_7027),
.Y(n_9395)
);

BUFx3_ASAP7_75t_L g9396 ( 
.A(n_8159),
.Y(n_9396)
);

OR2x2_ASAP7_75t_L g9397 ( 
.A(n_8411),
.B(n_6735),
.Y(n_9397)
);

OAI21x1_ASAP7_75t_L g9398 ( 
.A1(n_7932),
.A2(n_8066),
.B(n_8409),
.Y(n_9398)
);

CKINVDCx16_ASAP7_75t_R g9399 ( 
.A(n_8131),
.Y(n_9399)
);

AND2x4_ASAP7_75t_L g9400 ( 
.A(n_8209),
.B(n_7590),
.Y(n_9400)
);

CKINVDCx5p33_ASAP7_75t_R g9401 ( 
.A(n_8213),
.Y(n_9401)
);

NOR2x1_ASAP7_75t_SL g9402 ( 
.A(n_7971),
.B(n_7626),
.Y(n_9402)
);

BUFx2_ASAP7_75t_L g9403 ( 
.A(n_8524),
.Y(n_9403)
);

INVx1_ASAP7_75t_SL g9404 ( 
.A(n_8642),
.Y(n_9404)
);

INVx1_ASAP7_75t_L g9405 ( 
.A(n_8916),
.Y(n_9405)
);

AOI22x1_ASAP7_75t_L g9406 ( 
.A1(n_7811),
.A2(n_6556),
.B1(n_6731),
.B2(n_7453),
.Y(n_9406)
);

AOI22x1_ASAP7_75t_L g9407 ( 
.A1(n_7811),
.A2(n_7843),
.B1(n_7902),
.B2(n_8081),
.Y(n_9407)
);

NOR2xp33_ASAP7_75t_L g9408 ( 
.A(n_7947),
.B(n_7027),
.Y(n_9408)
);

AOI21xp5_ASAP7_75t_L g9409 ( 
.A1(n_7838),
.A2(n_6700),
.B(n_6938),
.Y(n_9409)
);

INVx1_ASAP7_75t_L g9410 ( 
.A(n_8916),
.Y(n_9410)
);

INVx2_ASAP7_75t_SL g9411 ( 
.A(n_8767),
.Y(n_9411)
);

AO21x2_ASAP7_75t_L g9412 ( 
.A1(n_8110),
.A2(n_6964),
.B(n_6831),
.Y(n_9412)
);

OAI21xp5_ASAP7_75t_L g9413 ( 
.A1(n_7795),
.A2(n_7626),
.B(n_7208),
.Y(n_9413)
);

AO21x1_ASAP7_75t_L g9414 ( 
.A1(n_8091),
.A2(n_7194),
.B(n_7029),
.Y(n_9414)
);

O2A1O1Ixp33_ASAP7_75t_L g9415 ( 
.A1(n_7768),
.A2(n_7626),
.B(n_7346),
.C(n_7339),
.Y(n_9415)
);

AOI21xp5_ASAP7_75t_L g9416 ( 
.A1(n_7838),
.A2(n_6969),
.B(n_6960),
.Y(n_9416)
);

OAI21x1_ASAP7_75t_L g9417 ( 
.A1(n_8099),
.A2(n_8108),
.B(n_8101),
.Y(n_9417)
);

NAND2xp5_ASAP7_75t_L g9418 ( 
.A(n_8356),
.B(n_6272),
.Y(n_9418)
);

HB1xp67_ASAP7_75t_L g9419 ( 
.A(n_8916),
.Y(n_9419)
);

INVx1_ASAP7_75t_L g9420 ( 
.A(n_8916),
.Y(n_9420)
);

INVx1_ASAP7_75t_L g9421 ( 
.A(n_8916),
.Y(n_9421)
);

CKINVDCx11_ASAP7_75t_R g9422 ( 
.A(n_8254),
.Y(n_9422)
);

CKINVDCx20_ASAP7_75t_R g9423 ( 
.A(n_8251),
.Y(n_9423)
);

INVxp67_ASAP7_75t_SL g9424 ( 
.A(n_8652),
.Y(n_9424)
);

NAND3xp33_ASAP7_75t_L g9425 ( 
.A(n_7816),
.B(n_6969),
.C(n_7359),
.Y(n_9425)
);

NAND2xp5_ASAP7_75t_L g9426 ( 
.A(n_8357),
.B(n_6272),
.Y(n_9426)
);

HB1xp67_ASAP7_75t_L g9427 ( 
.A(n_8916),
.Y(n_9427)
);

BUFx2_ASAP7_75t_R g9428 ( 
.A(n_8090),
.Y(n_9428)
);

INVx1_ASAP7_75t_L g9429 ( 
.A(n_8916),
.Y(n_9429)
);

INVx1_ASAP7_75t_L g9430 ( 
.A(n_8916),
.Y(n_9430)
);

OAI21xp5_ASAP7_75t_L g9431 ( 
.A1(n_7795),
.A2(n_7194),
.B(n_7208),
.Y(n_9431)
);

NAND2xp5_ASAP7_75t_L g9432 ( 
.A(n_8357),
.B(n_7812),
.Y(n_9432)
);

AOI22xp33_ASAP7_75t_L g9433 ( 
.A1(n_7978),
.A2(n_7649),
.B1(n_7549),
.B2(n_6960),
.Y(n_9433)
);

OAI21x1_ASAP7_75t_L g9434 ( 
.A1(n_8099),
.A2(n_8108),
.B(n_8101),
.Y(n_9434)
);

OA21x2_ASAP7_75t_L g9435 ( 
.A1(n_8490),
.A2(n_6900),
.B(n_6843),
.Y(n_9435)
);

INVx1_ASAP7_75t_L g9436 ( 
.A(n_8916),
.Y(n_9436)
);

NAND2xp5_ASAP7_75t_L g9437 ( 
.A(n_7812),
.B(n_6272),
.Y(n_9437)
);

INVx1_ASAP7_75t_L g9438 ( 
.A(n_8920),
.Y(n_9438)
);

OA21x2_ASAP7_75t_L g9439 ( 
.A1(n_8490),
.A2(n_6868),
.B(n_6900),
.Y(n_9439)
);

NOR2x1_ASAP7_75t_R g9440 ( 
.A(n_8645),
.B(n_6640),
.Y(n_9440)
);

INVx8_ASAP7_75t_L g9441 ( 
.A(n_8943),
.Y(n_9441)
);

AND2x4_ASAP7_75t_L g9442 ( 
.A(n_8209),
.B(n_8378),
.Y(n_9442)
);

AOI22x1_ASAP7_75t_L g9443 ( 
.A1(n_7811),
.A2(n_7107),
.B1(n_6700),
.B2(n_6776),
.Y(n_9443)
);

OR2x6_ASAP7_75t_L g9444 ( 
.A(n_8457),
.B(n_6640),
.Y(n_9444)
);

INVx3_ASAP7_75t_L g9445 ( 
.A(n_8209),
.Y(n_9445)
);

AOI221xp5_ASAP7_75t_L g9446 ( 
.A1(n_7816),
.A2(n_6776),
.B1(n_6969),
.B2(n_6960),
.C(n_7233),
.Y(n_9446)
);

OA21x2_ASAP7_75t_L g9447 ( 
.A1(n_8490),
.A2(n_6868),
.B(n_6900),
.Y(n_9447)
);

NOR2xp67_ASAP7_75t_L g9448 ( 
.A(n_7810),
.B(n_7861),
.Y(n_9448)
);

AO21x2_ASAP7_75t_L g9449 ( 
.A1(n_8963),
.A2(n_6905),
.B(n_7053),
.Y(n_9449)
);

INVx1_ASAP7_75t_L g9450 ( 
.A(n_8920),
.Y(n_9450)
);

BUFx2_ASAP7_75t_L g9451 ( 
.A(n_8524),
.Y(n_9451)
);

INVx3_ASAP7_75t_L g9452 ( 
.A(n_8378),
.Y(n_9452)
);

BUFx3_ASAP7_75t_L g9453 ( 
.A(n_8378),
.Y(n_9453)
);

NAND2x1p5_ASAP7_75t_L g9454 ( 
.A(n_7810),
.B(n_6640),
.Y(n_9454)
);

BUFx6f_ASAP7_75t_L g9455 ( 
.A(n_8549),
.Y(n_9455)
);

BUFx6f_ASAP7_75t_L g9456 ( 
.A(n_8549),
.Y(n_9456)
);

NAND2xp5_ASAP7_75t_L g9457 ( 
.A(n_8196),
.B(n_6272),
.Y(n_9457)
);

NOR2xp33_ASAP7_75t_L g9458 ( 
.A(n_8017),
.B(n_7027),
.Y(n_9458)
);

NAND2xp5_ASAP7_75t_L g9459 ( 
.A(n_8196),
.B(n_6272),
.Y(n_9459)
);

BUFx3_ASAP7_75t_L g9460 ( 
.A(n_8401),
.Y(n_9460)
);

BUFx3_ASAP7_75t_L g9461 ( 
.A(n_8401),
.Y(n_9461)
);

OA21x2_ASAP7_75t_L g9462 ( 
.A1(n_8490),
.A2(n_6964),
.B(n_7053),
.Y(n_9462)
);

INVx1_ASAP7_75t_L g9463 ( 
.A(n_8920),
.Y(n_9463)
);

NAND2x1p5_ASAP7_75t_L g9464 ( 
.A(n_7810),
.B(n_6640),
.Y(n_9464)
);

INVx1_ASAP7_75t_L g9465 ( 
.A(n_8920),
.Y(n_9465)
);

AND2x4_ASAP7_75t_L g9466 ( 
.A(n_8401),
.B(n_7270),
.Y(n_9466)
);

NAND3xp33_ASAP7_75t_L g9467 ( 
.A(n_7806),
.B(n_7324),
.C(n_6938),
.Y(n_9467)
);

BUFx6f_ASAP7_75t_L g9468 ( 
.A(n_8549),
.Y(n_9468)
);

NAND2xp5_ASAP7_75t_L g9469 ( 
.A(n_8221),
.B(n_6618),
.Y(n_9469)
);

AO21x2_ASAP7_75t_L g9470 ( 
.A1(n_8963),
.A2(n_6868),
.B(n_6905),
.Y(n_9470)
);

OAI21x1_ASAP7_75t_L g9471 ( 
.A1(n_8115),
.A2(n_8123),
.B(n_8117),
.Y(n_9471)
);

BUFx3_ASAP7_75t_L g9472 ( 
.A(n_8401),
.Y(n_9472)
);

OAI21xp5_ASAP7_75t_L g9473 ( 
.A1(n_7987),
.A2(n_7800),
.B(n_7910),
.Y(n_9473)
);

NAND2xp5_ASAP7_75t_L g9474 ( 
.A(n_8221),
.B(n_6618),
.Y(n_9474)
);

OAI21xp5_ASAP7_75t_L g9475 ( 
.A1(n_7987),
.A2(n_6767),
.B(n_7432),
.Y(n_9475)
);

BUFx6f_ASAP7_75t_L g9476 ( 
.A(n_8581),
.Y(n_9476)
);

CKINVDCx5p33_ASAP7_75t_R g9477 ( 
.A(n_8213),
.Y(n_9477)
);

OA21x2_ASAP7_75t_L g9478 ( 
.A1(n_8491),
.A2(n_6905),
.B(n_6930),
.Y(n_9478)
);

INVx1_ASAP7_75t_L g9479 ( 
.A(n_8920),
.Y(n_9479)
);

INVx1_ASAP7_75t_L g9480 ( 
.A(n_8920),
.Y(n_9480)
);

INVx1_ASAP7_75t_L g9481 ( 
.A(n_8920),
.Y(n_9481)
);

INVx2_ASAP7_75t_SL g9482 ( 
.A(n_8767),
.Y(n_9482)
);

INVx1_ASAP7_75t_L g9483 ( 
.A(n_8920),
.Y(n_9483)
);

OA21x2_ASAP7_75t_L g9484 ( 
.A1(n_8491),
.A2(n_6973),
.B(n_6964),
.Y(n_9484)
);

HB1xp67_ASAP7_75t_L g9485 ( 
.A(n_8920),
.Y(n_9485)
);

INVxp67_ASAP7_75t_SL g9486 ( 
.A(n_8765),
.Y(n_9486)
);

BUFx2_ASAP7_75t_L g9487 ( 
.A(n_8524),
.Y(n_9487)
);

OAI21xp5_ASAP7_75t_L g9488 ( 
.A1(n_7800),
.A2(n_7459),
.B(n_7208),
.Y(n_9488)
);

BUFx12f_ASAP7_75t_L g9489 ( 
.A(n_8648),
.Y(n_9489)
);

INVx3_ASAP7_75t_L g9490 ( 
.A(n_8421),
.Y(n_9490)
);

INVx1_ASAP7_75t_L g9491 ( 
.A(n_8930),
.Y(n_9491)
);

AND2x2_ASAP7_75t_L g9492 ( 
.A(n_7774),
.B(n_7027),
.Y(n_9492)
);

INVx1_ASAP7_75t_SL g9493 ( 
.A(n_8810),
.Y(n_9493)
);

INVx1_ASAP7_75t_L g9494 ( 
.A(n_8930),
.Y(n_9494)
);

BUFx4f_ASAP7_75t_L g9495 ( 
.A(n_7971),
.Y(n_9495)
);

OA21x2_ASAP7_75t_L g9496 ( 
.A1(n_8491),
.A2(n_7042),
.B(n_7215),
.Y(n_9496)
);

BUFx2_ASAP7_75t_R g9497 ( 
.A(n_8090),
.Y(n_9497)
);

NOR2xp33_ASAP7_75t_L g9498 ( 
.A(n_8017),
.B(n_7042),
.Y(n_9498)
);

AND2x2_ASAP7_75t_L g9499 ( 
.A(n_7774),
.B(n_7042),
.Y(n_9499)
);

INVx1_ASAP7_75t_L g9500 ( 
.A(n_8930),
.Y(n_9500)
);

OAI21xp5_ASAP7_75t_L g9501 ( 
.A1(n_7910),
.A2(n_7459),
.B(n_7208),
.Y(n_9501)
);

OAI21xp5_ASAP7_75t_L g9502 ( 
.A1(n_7978),
.A2(n_7459),
.B(n_7208),
.Y(n_9502)
);

NOR2xp33_ASAP7_75t_SL g9503 ( 
.A(n_8023),
.B(n_6288),
.Y(n_9503)
);

OAI21x1_ASAP7_75t_SL g9504 ( 
.A1(n_7728),
.A2(n_6832),
.B(n_6493),
.Y(n_9504)
);

OAI21x1_ASAP7_75t_SL g9505 ( 
.A1(n_7728),
.A2(n_6832),
.B(n_6493),
.Y(n_9505)
);

NAND2xp5_ASAP7_75t_L g9506 ( 
.A(n_7854),
.B(n_6618),
.Y(n_9506)
);

CKINVDCx5p33_ASAP7_75t_R g9507 ( 
.A(n_8663),
.Y(n_9507)
);

AND2x2_ASAP7_75t_L g9508 ( 
.A(n_8759),
.B(n_8824),
.Y(n_9508)
);

BUFx4f_ASAP7_75t_SL g9509 ( 
.A(n_8439),
.Y(n_9509)
);

AND2x4_ASAP7_75t_L g9510 ( 
.A(n_8421),
.B(n_6640),
.Y(n_9510)
);

BUFx2_ASAP7_75t_R g9511 ( 
.A(n_8090),
.Y(n_9511)
);

AO21x2_ASAP7_75t_L g9512 ( 
.A1(n_7972),
.A2(n_7215),
.B(n_7511),
.Y(n_9512)
);

OA21x2_ASAP7_75t_L g9513 ( 
.A1(n_8491),
.A2(n_7042),
.B(n_7211),
.Y(n_9513)
);

AND2x2_ASAP7_75t_L g9514 ( 
.A(n_8759),
.B(n_6735),
.Y(n_9514)
);

AOI22xp5_ASAP7_75t_L g9515 ( 
.A1(n_7770),
.A2(n_6338),
.B1(n_7649),
.B2(n_6570),
.Y(n_9515)
);

INVx1_ASAP7_75t_L g9516 ( 
.A(n_8930),
.Y(n_9516)
);

OAI21x1_ASAP7_75t_SL g9517 ( 
.A1(n_7728),
.A2(n_6832),
.B(n_6288),
.Y(n_9517)
);

AO21x2_ASAP7_75t_L g9518 ( 
.A1(n_7972),
.A2(n_7211),
.B(n_7512),
.Y(n_9518)
);

BUFx2_ASAP7_75t_L g9519 ( 
.A(n_8524),
.Y(n_9519)
);

AND2x4_ASAP7_75t_L g9520 ( 
.A(n_8421),
.B(n_6640),
.Y(n_9520)
);

INVx1_ASAP7_75t_L g9521 ( 
.A(n_8930),
.Y(n_9521)
);

OAI21x1_ASAP7_75t_L g9522 ( 
.A1(n_8450),
.A2(n_8128),
.B(n_8376),
.Y(n_9522)
);

AND2x2_ASAP7_75t_L g9523 ( 
.A(n_8759),
.B(n_6735),
.Y(n_9523)
);

AOI21xp33_ASAP7_75t_L g9524 ( 
.A1(n_7865),
.A2(n_7211),
.B(n_7532),
.Y(n_9524)
);

INVx1_ASAP7_75t_L g9525 ( 
.A(n_8930),
.Y(n_9525)
);

BUFx3_ASAP7_75t_L g9526 ( 
.A(n_8421),
.Y(n_9526)
);

INVx1_ASAP7_75t_L g9527 ( 
.A(n_8930),
.Y(n_9527)
);

NAND3xp33_ASAP7_75t_L g9528 ( 
.A(n_7841),
.B(n_7891),
.C(n_7797),
.Y(n_9528)
);

BUFx3_ASAP7_75t_L g9529 ( 
.A(n_8440),
.Y(n_9529)
);

NOR2xp33_ASAP7_75t_L g9530 ( 
.A(n_7797),
.B(n_7380),
.Y(n_9530)
);

OAI21xp5_ASAP7_75t_L g9531 ( 
.A1(n_7871),
.A2(n_7459),
.B(n_7208),
.Y(n_9531)
);

INVx1_ASAP7_75t_L g9532 ( 
.A(n_8930),
.Y(n_9532)
);

OAI21x1_ASAP7_75t_SL g9533 ( 
.A1(n_8830),
.A2(n_6832),
.B(n_6288),
.Y(n_9533)
);

NOR2xp33_ASAP7_75t_L g9534 ( 
.A(n_7797),
.B(n_7402),
.Y(n_9534)
);

NAND2x1p5_ASAP7_75t_L g9535 ( 
.A(n_7810),
.B(n_6640),
.Y(n_9535)
);

NOR2xp33_ASAP7_75t_L g9536 ( 
.A(n_7833),
.B(n_7402),
.Y(n_9536)
);

NOR2xp67_ASAP7_75t_L g9537 ( 
.A(n_7810),
.B(n_7402),
.Y(n_9537)
);

AND2x2_ASAP7_75t_L g9538 ( 
.A(n_8759),
.B(n_7569),
.Y(n_9538)
);

INVxp67_ASAP7_75t_SL g9539 ( 
.A(n_8765),
.Y(n_9539)
);

NAND2x1p5_ASAP7_75t_L g9540 ( 
.A(n_7810),
.B(n_6640),
.Y(n_9540)
);

OR2x2_ASAP7_75t_L g9541 ( 
.A(n_8411),
.B(n_6618),
.Y(n_9541)
);

BUFx4f_ASAP7_75t_L g9542 ( 
.A(n_8070),
.Y(n_9542)
);

INVx3_ASAP7_75t_L g9543 ( 
.A(n_8440),
.Y(n_9543)
);

NOR2xp33_ASAP7_75t_L g9544 ( 
.A(n_7833),
.B(n_8135),
.Y(n_9544)
);

NOR2xp33_ASAP7_75t_L g9545 ( 
.A(n_7833),
.B(n_7402),
.Y(n_9545)
);

AOI21xp5_ASAP7_75t_L g9546 ( 
.A1(n_8164),
.A2(n_6969),
.B(n_6776),
.Y(n_9546)
);

AND2x2_ASAP7_75t_L g9547 ( 
.A(n_8824),
.B(n_7569),
.Y(n_9547)
);

OA21x2_ASAP7_75t_L g9548 ( 
.A1(n_8500),
.A2(n_7211),
.B(n_7392),
.Y(n_9548)
);

INVx2_ASAP7_75t_SL g9549 ( 
.A(n_8767),
.Y(n_9549)
);

BUFx3_ASAP7_75t_L g9550 ( 
.A(n_8440),
.Y(n_9550)
);

AOI21x1_ASAP7_75t_L g9551 ( 
.A1(n_7913),
.A2(n_7511),
.B(n_7475),
.Y(n_9551)
);

AO21x1_ASAP7_75t_L g9552 ( 
.A1(n_8121),
.A2(n_7431),
.B(n_7350),
.Y(n_9552)
);

INVx3_ASAP7_75t_L g9553 ( 
.A(n_8440),
.Y(n_9553)
);

OAI22xp5_ASAP7_75t_L g9554 ( 
.A1(n_7909),
.A2(n_7569),
.B1(n_7549),
.B2(n_7437),
.Y(n_9554)
);

BUFx2_ASAP7_75t_R g9555 ( 
.A(n_7693),
.Y(n_9555)
);

INVxp67_ASAP7_75t_L g9556 ( 
.A(n_8328),
.Y(n_9556)
);

OAI21x1_ASAP7_75t_L g9557 ( 
.A1(n_8376),
.A2(n_8161),
.B(n_8359),
.Y(n_9557)
);

OAI21x1_ASAP7_75t_SL g9558 ( 
.A1(n_8830),
.A2(n_6832),
.B(n_6493),
.Y(n_9558)
);

INVx1_ASAP7_75t_L g9559 ( 
.A(n_8242),
.Y(n_9559)
);

OAI21xp5_ASAP7_75t_L g9560 ( 
.A1(n_7871),
.A2(n_8002),
.B(n_7951),
.Y(n_9560)
);

BUFx3_ASAP7_75t_L g9561 ( 
.A(n_8345),
.Y(n_9561)
);

INVx1_ASAP7_75t_L g9562 ( 
.A(n_8242),
.Y(n_9562)
);

AOI22x1_ASAP7_75t_L g9563 ( 
.A1(n_7902),
.A2(n_7233),
.B1(n_6938),
.B2(n_6960),
.Y(n_9563)
);

HB1xp67_ASAP7_75t_L g9564 ( 
.A(n_8242),
.Y(n_9564)
);

NAND2xp5_ASAP7_75t_L g9565 ( 
.A(n_7854),
.B(n_6618),
.Y(n_9565)
);

BUFx6f_ASAP7_75t_L g9566 ( 
.A(n_8581),
.Y(n_9566)
);

AND2x2_ASAP7_75t_L g9567 ( 
.A(n_8824),
.B(n_7569),
.Y(n_9567)
);

INVx2_ASAP7_75t_SL g9568 ( 
.A(n_8767),
.Y(n_9568)
);

AO21x2_ASAP7_75t_L g9569 ( 
.A1(n_8014),
.A2(n_7392),
.B(n_7352),
.Y(n_9569)
);

AOI21xp5_ASAP7_75t_L g9570 ( 
.A1(n_8164),
.A2(n_6731),
.B(n_7453),
.Y(n_9570)
);

AND2x4_ASAP7_75t_L g9571 ( 
.A(n_8767),
.B(n_6677),
.Y(n_9571)
);

AO21x2_ASAP7_75t_L g9572 ( 
.A1(n_8014),
.A2(n_7392),
.B(n_7352),
.Y(n_9572)
);

BUFx3_ASAP7_75t_L g9573 ( 
.A(n_8346),
.Y(n_9573)
);

BUFx2_ASAP7_75t_SL g9574 ( 
.A(n_7847),
.Y(n_9574)
);

AND2x4_ASAP7_75t_L g9575 ( 
.A(n_8767),
.B(n_6677),
.Y(n_9575)
);

INVx1_ASAP7_75t_L g9576 ( 
.A(n_8242),
.Y(n_9576)
);

INVx8_ASAP7_75t_L g9577 ( 
.A(n_8943),
.Y(n_9577)
);

INVx1_ASAP7_75t_SL g9578 ( 
.A(n_8810),
.Y(n_9578)
);

AO21x1_ASAP7_75t_L g9579 ( 
.A1(n_8121),
.A2(n_7431),
.B(n_7430),
.Y(n_9579)
);

NAND2xp5_ASAP7_75t_L g9580 ( 
.A(n_7852),
.B(n_6618),
.Y(n_9580)
);

AND2x2_ASAP7_75t_L g9581 ( 
.A(n_8824),
.B(n_7569),
.Y(n_9581)
);

BUFx3_ASAP7_75t_L g9582 ( 
.A(n_8346),
.Y(n_9582)
);

INVx4_ASAP7_75t_L g9583 ( 
.A(n_8070),
.Y(n_9583)
);

OAI21x1_ASAP7_75t_SL g9584 ( 
.A1(n_8830),
.A2(n_6832),
.B(n_6493),
.Y(n_9584)
);

NOR2x1_ASAP7_75t_R g9585 ( 
.A(n_8648),
.B(n_6677),
.Y(n_9585)
);

INVx1_ASAP7_75t_L g9586 ( 
.A(n_8242),
.Y(n_9586)
);

INVx5_ASAP7_75t_L g9587 ( 
.A(n_8581),
.Y(n_9587)
);

INVx1_ASAP7_75t_L g9588 ( 
.A(n_8242),
.Y(n_9588)
);

BUFx3_ASAP7_75t_L g9589 ( 
.A(n_8370),
.Y(n_9589)
);

AO21x2_ASAP7_75t_L g9590 ( 
.A1(n_8288),
.A2(n_8557),
.B(n_8544),
.Y(n_9590)
);

NOR2xp33_ASAP7_75t_L g9591 ( 
.A(n_8135),
.B(n_8152),
.Y(n_9591)
);

INVx4_ASAP7_75t_L g9592 ( 
.A(n_8070),
.Y(n_9592)
);

INVx2_ASAP7_75t_L g9593 ( 
.A(n_8269),
.Y(n_9593)
);

INVx1_ASAP7_75t_L g9594 ( 
.A(n_8269),
.Y(n_9594)
);

INVx1_ASAP7_75t_SL g9595 ( 
.A(n_8810),
.Y(n_9595)
);

BUFx3_ASAP7_75t_L g9596 ( 
.A(n_8370),
.Y(n_9596)
);

OR2x2_ASAP7_75t_L g9597 ( 
.A(n_8411),
.B(n_6618),
.Y(n_9597)
);

INVx2_ASAP7_75t_SL g9598 ( 
.A(n_8767),
.Y(n_9598)
);

NAND2xp5_ASAP7_75t_L g9599 ( 
.A(n_7852),
.B(n_6618),
.Y(n_9599)
);

BUFx3_ASAP7_75t_L g9600 ( 
.A(n_8370),
.Y(n_9600)
);

CKINVDCx5p33_ASAP7_75t_R g9601 ( 
.A(n_8663),
.Y(n_9601)
);

INVx1_ASAP7_75t_L g9602 ( 
.A(n_8269),
.Y(n_9602)
);

OAI21xp5_ASAP7_75t_L g9603 ( 
.A1(n_8002),
.A2(n_7315),
.B(n_7234),
.Y(n_9603)
);

INVx2_ASAP7_75t_L g9604 ( 
.A(n_8269),
.Y(n_9604)
);

INVx2_ASAP7_75t_L g9605 ( 
.A(n_8269),
.Y(n_9605)
);

BUFx3_ASAP7_75t_L g9606 ( 
.A(n_8370),
.Y(n_9606)
);

NAND2xp5_ASAP7_75t_L g9607 ( 
.A(n_7935),
.B(n_6637),
.Y(n_9607)
);

CKINVDCx6p67_ASAP7_75t_R g9608 ( 
.A(n_8608),
.Y(n_9608)
);

AOI21x1_ASAP7_75t_L g9609 ( 
.A1(n_8341),
.A2(n_7514),
.B(n_7475),
.Y(n_9609)
);

AOI22xp33_ASAP7_75t_L g9610 ( 
.A1(n_7909),
.A2(n_6969),
.B1(n_7324),
.B2(n_7233),
.Y(n_9610)
);

OAI21xp5_ASAP7_75t_L g9611 ( 
.A1(n_8002),
.A2(n_7432),
.B(n_7431),
.Y(n_9611)
);

AOI22xp33_ASAP7_75t_L g9612 ( 
.A1(n_7909),
.A2(n_6960),
.B1(n_7233),
.B2(n_7321),
.Y(n_9612)
);

INVx2_ASAP7_75t_SL g9613 ( 
.A(n_8767),
.Y(n_9613)
);

INVx4_ASAP7_75t_L g9614 ( 
.A(n_8070),
.Y(n_9614)
);

NOR2xp33_ASAP7_75t_L g9615 ( 
.A(n_8152),
.B(n_6507),
.Y(n_9615)
);

OAI21x1_ASAP7_75t_L g9616 ( 
.A1(n_8139),
.A2(n_6465),
.B(n_6574),
.Y(n_9616)
);

NAND2xp5_ASAP7_75t_L g9617 ( 
.A(n_7935),
.B(n_6637),
.Y(n_9617)
);

INVx1_ASAP7_75t_L g9618 ( 
.A(n_8269),
.Y(n_9618)
);

O2A1O1Ixp33_ASAP7_75t_L g9619 ( 
.A1(n_7951),
.A2(n_6767),
.B(n_7231),
.C(n_7194),
.Y(n_9619)
);

INVx3_ASAP7_75t_L g9620 ( 
.A(n_8581),
.Y(n_9620)
);

HB1xp67_ASAP7_75t_L g9621 ( 
.A(n_8307),
.Y(n_9621)
);

INVx1_ASAP7_75t_SL g9622 ( 
.A(n_8810),
.Y(n_9622)
);

INVx1_ASAP7_75t_L g9623 ( 
.A(n_8307),
.Y(n_9623)
);

OAI21x1_ASAP7_75t_L g9624 ( 
.A1(n_8141),
.A2(n_6574),
.B(n_6525),
.Y(n_9624)
);

NOR2xp33_ASAP7_75t_SL g9625 ( 
.A(n_8092),
.B(n_6288),
.Y(n_9625)
);

CKINVDCx20_ASAP7_75t_R g9626 ( 
.A(n_8251),
.Y(n_9626)
);

OAI21x1_ASAP7_75t_L g9627 ( 
.A1(n_8141),
.A2(n_8142),
.B(n_7939),
.Y(n_9627)
);

AOI21xp5_ASAP7_75t_L g9628 ( 
.A1(n_8166),
.A2(n_6731),
.B(n_7324),
.Y(n_9628)
);

BUFx6f_ASAP7_75t_L g9629 ( 
.A(n_8581),
.Y(n_9629)
);

OAI21xp5_ASAP7_75t_L g9630 ( 
.A1(n_7963),
.A2(n_7955),
.B(n_7937),
.Y(n_9630)
);

OAI21x1_ASAP7_75t_SL g9631 ( 
.A1(n_7941),
.A2(n_7920),
.B(n_8530),
.Y(n_9631)
);

INVx1_ASAP7_75t_L g9632 ( 
.A(n_8307),
.Y(n_9632)
);

OAI21x1_ASAP7_75t_L g9633 ( 
.A1(n_8141),
.A2(n_6574),
.B(n_6525),
.Y(n_9633)
);

INVx1_ASAP7_75t_L g9634 ( 
.A(n_8307),
.Y(n_9634)
);

INVxp33_ASAP7_75t_L g9635 ( 
.A(n_7977),
.Y(n_9635)
);

INVx5_ASAP7_75t_L g9636 ( 
.A(n_8581),
.Y(n_9636)
);

INVx2_ASAP7_75t_SL g9637 ( 
.A(n_8767),
.Y(n_9637)
);

AOI21xp5_ASAP7_75t_L g9638 ( 
.A1(n_8166),
.A2(n_6731),
.B(n_7324),
.Y(n_9638)
);

AOI21xp5_ASAP7_75t_L g9639 ( 
.A1(n_8385),
.A2(n_8397),
.B(n_8134),
.Y(n_9639)
);

NAND2xp5_ASAP7_75t_L g9640 ( 
.A(n_7942),
.B(n_6637),
.Y(n_9640)
);

AND2x2_ASAP7_75t_L g9641 ( 
.A(n_8845),
.B(n_6637),
.Y(n_9641)
);

OAI21x1_ASAP7_75t_SL g9642 ( 
.A1(n_7941),
.A2(n_6832),
.B(n_6288),
.Y(n_9642)
);

NAND2x1p5_ASAP7_75t_L g9643 ( 
.A(n_7810),
.B(n_6731),
.Y(n_9643)
);

NAND2x1p5_ASAP7_75t_L g9644 ( 
.A(n_7810),
.B(n_6731),
.Y(n_9644)
);

OAI21x1_ASAP7_75t_SL g9645 ( 
.A1(n_7941),
.A2(n_6288),
.B(n_6493),
.Y(n_9645)
);

NAND2xp5_ASAP7_75t_L g9646 ( 
.A(n_7942),
.B(n_6637),
.Y(n_9646)
);

NAND3xp33_ASAP7_75t_L g9647 ( 
.A(n_7891),
.B(n_6960),
.C(n_7324),
.Y(n_9647)
);

AND2x2_ASAP7_75t_L g9648 ( 
.A(n_8845),
.B(n_6637),
.Y(n_9648)
);

INVx2_ASAP7_75t_L g9649 ( 
.A(n_8307),
.Y(n_9649)
);

AND2x2_ASAP7_75t_L g9650 ( 
.A(n_8845),
.B(n_6637),
.Y(n_9650)
);

AND2x4_ASAP7_75t_L g9651 ( 
.A(n_8767),
.B(n_6969),
.Y(n_9651)
);

HB1xp67_ASAP7_75t_L g9652 ( 
.A(n_8307),
.Y(n_9652)
);

BUFx6f_ASAP7_75t_L g9653 ( 
.A(n_8581),
.Y(n_9653)
);

BUFx3_ASAP7_75t_L g9654 ( 
.A(n_8370),
.Y(n_9654)
);

AOI21xp5_ASAP7_75t_L g9655 ( 
.A1(n_8385),
.A2(n_6938),
.B(n_7359),
.Y(n_9655)
);

INVx1_ASAP7_75t_L g9656 ( 
.A(n_8765),
.Y(n_9656)
);

AOI22xp33_ASAP7_75t_L g9657 ( 
.A1(n_7770),
.A2(n_7321),
.B1(n_7324),
.B2(n_7233),
.Y(n_9657)
);

BUFx6f_ASAP7_75t_L g9658 ( 
.A(n_8581),
.Y(n_9658)
);

INVx3_ASAP7_75t_L g9659 ( 
.A(n_8581),
.Y(n_9659)
);

BUFx4f_ASAP7_75t_SL g9660 ( 
.A(n_8439),
.Y(n_9660)
);

INVx1_ASAP7_75t_L g9661 ( 
.A(n_8875),
.Y(n_9661)
);

OAI21x1_ASAP7_75t_SL g9662 ( 
.A1(n_7920),
.A2(n_6317),
.B(n_6493),
.Y(n_9662)
);

INVx2_ASAP7_75t_L g9663 ( 
.A(n_8810),
.Y(n_9663)
);

INVx1_ASAP7_75t_L g9664 ( 
.A(n_8875),
.Y(n_9664)
);

OAI21xp5_ASAP7_75t_L g9665 ( 
.A1(n_7963),
.A2(n_7012),
.B(n_7491),
.Y(n_9665)
);

BUFx3_ASAP7_75t_L g9666 ( 
.A(n_8370),
.Y(n_9666)
);

AND2x2_ASAP7_75t_L g9667 ( 
.A(n_8845),
.B(n_8854),
.Y(n_9667)
);

NOR2xp33_ASAP7_75t_R g9668 ( 
.A(n_7953),
.B(n_6317),
.Y(n_9668)
);

BUFx12f_ASAP7_75t_L g9669 ( 
.A(n_7693),
.Y(n_9669)
);

INVx4_ASAP7_75t_L g9670 ( 
.A(n_8070),
.Y(n_9670)
);

AND2x2_ASAP7_75t_L g9671 ( 
.A(n_8854),
.B(n_6637),
.Y(n_9671)
);

BUFx3_ASAP7_75t_L g9672 ( 
.A(n_8370),
.Y(n_9672)
);

INVx1_ASAP7_75t_L g9673 ( 
.A(n_8875),
.Y(n_9673)
);

OAI21x1_ASAP7_75t_L g9674 ( 
.A1(n_8056),
.A2(n_8060),
.B(n_8582),
.Y(n_9674)
);

AOI22x1_ASAP7_75t_L g9675 ( 
.A1(n_7902),
.A2(n_6938),
.B1(n_6776),
.B2(n_7359),
.Y(n_9675)
);

NAND2xp5_ASAP7_75t_L g9676 ( 
.A(n_8897),
.B(n_7222),
.Y(n_9676)
);

NOR2xp67_ASAP7_75t_L g9677 ( 
.A(n_7810),
.B(n_7861),
.Y(n_9677)
);

INVxp67_ASAP7_75t_SL g9678 ( 
.A(n_8575),
.Y(n_9678)
);

OA21x2_ASAP7_75t_L g9679 ( 
.A1(n_8532),
.A2(n_8552),
.B(n_8555),
.Y(n_9679)
);

NAND2xp5_ASAP7_75t_L g9680 ( 
.A(n_8897),
.B(n_7222),
.Y(n_9680)
);

AOI22xp5_ASAP7_75t_L g9681 ( 
.A1(n_7803),
.A2(n_7012),
.B1(n_7029),
.B2(n_7452),
.Y(n_9681)
);

INVxp67_ASAP7_75t_SL g9682 ( 
.A(n_8575),
.Y(n_9682)
);

INVx4_ASAP7_75t_L g9683 ( 
.A(n_8070),
.Y(n_9683)
);

OR2x2_ASAP7_75t_L g9684 ( 
.A(n_7986),
.B(n_6837),
.Y(n_9684)
);

OAI21x1_ASAP7_75t_L g9685 ( 
.A1(n_8060),
.A2(n_8582),
.B(n_8430),
.Y(n_9685)
);

BUFx3_ASAP7_75t_L g9686 ( 
.A(n_8370),
.Y(n_9686)
);

OR2x2_ASAP7_75t_L g9687 ( 
.A(n_7986),
.B(n_6837),
.Y(n_9687)
);

BUFx6f_ASAP7_75t_L g9688 ( 
.A(n_8625),
.Y(n_9688)
);

CKINVDCx16_ASAP7_75t_R g9689 ( 
.A(n_8131),
.Y(n_9689)
);

OAI21x1_ASAP7_75t_L g9690 ( 
.A1(n_8582),
.A2(n_6997),
.B(n_6955),
.Y(n_9690)
);

NAND2xp5_ASAP7_75t_L g9691 ( 
.A(n_8173),
.B(n_7222),
.Y(n_9691)
);

INVx2_ASAP7_75t_L g9692 ( 
.A(n_8810),
.Y(n_9692)
);

OAI21x1_ASAP7_75t_L g9693 ( 
.A1(n_8582),
.A2(n_6997),
.B(n_6955),
.Y(n_9693)
);

INVx1_ASAP7_75t_SL g9694 ( 
.A(n_8810),
.Y(n_9694)
);

OAI21x1_ASAP7_75t_L g9695 ( 
.A1(n_8430),
.A2(n_6997),
.B(n_6955),
.Y(n_9695)
);

OAI21x1_ASAP7_75t_L g9696 ( 
.A1(n_8430),
.A2(n_6997),
.B(n_6955),
.Y(n_9696)
);

OAI21xp5_ASAP7_75t_L g9697 ( 
.A1(n_7955),
.A2(n_7350),
.B(n_7467),
.Y(n_9697)
);

AND2x4_ASAP7_75t_L g9698 ( 
.A(n_8074),
.B(n_7453),
.Y(n_9698)
);

OAI21xp5_ASAP7_75t_L g9699 ( 
.A1(n_7937),
.A2(n_7350),
.B(n_7467),
.Y(n_9699)
);

INVxp67_ASAP7_75t_SL g9700 ( 
.A(n_8575),
.Y(n_9700)
);

NAND2xp5_ASAP7_75t_L g9701 ( 
.A(n_8173),
.B(n_7222),
.Y(n_9701)
);

NAND2xp5_ASAP7_75t_L g9702 ( 
.A(n_8334),
.B(n_7222),
.Y(n_9702)
);

OAI21x1_ASAP7_75t_L g9703 ( 
.A1(n_8430),
.A2(n_6997),
.B(n_6955),
.Y(n_9703)
);

INVx1_ASAP7_75t_SL g9704 ( 
.A(n_7757),
.Y(n_9704)
);

INVx3_ASAP7_75t_L g9705 ( 
.A(n_8625),
.Y(n_9705)
);

INVx2_ASAP7_75t_SL g9706 ( 
.A(n_8817),
.Y(n_9706)
);

AOI22xp33_ASAP7_75t_L g9707 ( 
.A1(n_7983),
.A2(n_6969),
.B1(n_7321),
.B2(n_7233),
.Y(n_9707)
);

BUFx2_ASAP7_75t_L g9708 ( 
.A(n_8524),
.Y(n_9708)
);

NAND2x1p5_ASAP7_75t_L g9709 ( 
.A(n_7861),
.B(n_6938),
.Y(n_9709)
);

INVx2_ASAP7_75t_L g9710 ( 
.A(n_8465),
.Y(n_9710)
);

AOI21xp5_ASAP7_75t_L g9711 ( 
.A1(n_8397),
.A2(n_6938),
.B(n_7324),
.Y(n_9711)
);

NAND2x1p5_ASAP7_75t_L g9712 ( 
.A(n_7861),
.B(n_7324),
.Y(n_9712)
);

AO21x2_ASAP7_75t_L g9713 ( 
.A1(n_7845),
.A2(n_6767),
.B(n_7459),
.Y(n_9713)
);

BUFx2_ASAP7_75t_L g9714 ( 
.A(n_8524),
.Y(n_9714)
);

NOR2xp67_ASAP7_75t_L g9715 ( 
.A(n_7861),
.B(n_7324),
.Y(n_9715)
);

NAND2xp5_ASAP7_75t_L g9716 ( 
.A(n_8334),
.B(n_7222),
.Y(n_9716)
);

AOI21xp33_ASAP7_75t_L g9717 ( 
.A1(n_7865),
.A2(n_6969),
.B(n_7453),
.Y(n_9717)
);

INVx2_ASAP7_75t_L g9718 ( 
.A(n_8465),
.Y(n_9718)
);

OAI21x1_ASAP7_75t_SL g9719 ( 
.A1(n_8530),
.A2(n_6317),
.B(n_7581),
.Y(n_9719)
);

NAND2xp5_ASAP7_75t_L g9720 ( 
.A(n_8336),
.B(n_7222),
.Y(n_9720)
);

NAND2xp5_ASAP7_75t_L g9721 ( 
.A(n_8336),
.B(n_7222),
.Y(n_9721)
);

INVx2_ASAP7_75t_L g9722 ( 
.A(n_8465),
.Y(n_9722)
);

OA21x2_ASAP7_75t_L g9723 ( 
.A1(n_8555),
.A2(n_8289),
.B(n_8658),
.Y(n_9723)
);

INVx4_ASAP7_75t_L g9724 ( 
.A(n_8070),
.Y(n_9724)
);

INVx1_ASAP7_75t_SL g9725 ( 
.A(n_7757),
.Y(n_9725)
);

BUFx6f_ASAP7_75t_L g9726 ( 
.A(n_8625),
.Y(n_9726)
);

INVx3_ASAP7_75t_L g9727 ( 
.A(n_8625),
.Y(n_9727)
);

AND2x2_ASAP7_75t_L g9728 ( 
.A(n_8854),
.B(n_7315),
.Y(n_9728)
);

NOR2xp33_ASAP7_75t_L g9729 ( 
.A(n_7879),
.B(n_7452),
.Y(n_9729)
);

HB1xp67_ASAP7_75t_L g9730 ( 
.A(n_8465),
.Y(n_9730)
);

AND2x4_ASAP7_75t_L g9731 ( 
.A(n_8074),
.B(n_7453),
.Y(n_9731)
);

NOR2xp33_ASAP7_75t_SL g9732 ( 
.A(n_8092),
.B(n_6317),
.Y(n_9732)
);

BUFx3_ASAP7_75t_L g9733 ( 
.A(n_8370),
.Y(n_9733)
);

OAI21xp5_ASAP7_75t_L g9734 ( 
.A1(n_7853),
.A2(n_6727),
.B(n_7452),
.Y(n_9734)
);

OAI21xp5_ASAP7_75t_L g9735 ( 
.A1(n_7853),
.A2(n_6727),
.B(n_7452),
.Y(n_9735)
);

INVx6_ASAP7_75t_L g9736 ( 
.A(n_7735),
.Y(n_9736)
);

OAI21xp5_ASAP7_75t_L g9737 ( 
.A1(n_7944),
.A2(n_6727),
.B(n_7452),
.Y(n_9737)
);

INVx3_ASAP7_75t_SL g9738 ( 
.A(n_7756),
.Y(n_9738)
);

CKINVDCx11_ASAP7_75t_R g9739 ( 
.A(n_8558),
.Y(n_9739)
);

AND2x2_ASAP7_75t_L g9740 ( 
.A(n_8854),
.B(n_6692),
.Y(n_9740)
);

OA21x2_ASAP7_75t_L g9741 ( 
.A1(n_8555),
.A2(n_8289),
.B(n_8658),
.Y(n_9741)
);

OAI21x1_ASAP7_75t_SL g9742 ( 
.A1(n_8531),
.A2(n_6317),
.B(n_7581),
.Y(n_9742)
);

OAI21xp5_ASAP7_75t_L g9743 ( 
.A1(n_7944),
.A2(n_7234),
.B(n_7432),
.Y(n_9743)
);

INVx5_ASAP7_75t_L g9744 ( 
.A(n_8625),
.Y(n_9744)
);

AOI22xp33_ASAP7_75t_L g9745 ( 
.A1(n_7983),
.A2(n_7321),
.B1(n_7233),
.B2(n_7107),
.Y(n_9745)
);

AND2x2_ASAP7_75t_L g9746 ( 
.A(n_8859),
.B(n_6692),
.Y(n_9746)
);

INVx3_ASAP7_75t_L g9747 ( 
.A(n_8625),
.Y(n_9747)
);

HB1xp67_ASAP7_75t_L g9748 ( 
.A(n_8465),
.Y(n_9748)
);

NAND2xp5_ASAP7_75t_L g9749 ( 
.A(n_8848),
.B(n_7204),
.Y(n_9749)
);

NOR2xp67_ASAP7_75t_L g9750 ( 
.A(n_7861),
.B(n_7107),
.Y(n_9750)
);

NAND2xp5_ASAP7_75t_L g9751 ( 
.A(n_8848),
.B(n_7204),
.Y(n_9751)
);

INVx3_ASAP7_75t_L g9752 ( 
.A(n_8625),
.Y(n_9752)
);

NOR2xp33_ASAP7_75t_L g9753 ( 
.A(n_7866),
.B(n_7350),
.Y(n_9753)
);

INVx1_ASAP7_75t_L g9754 ( 
.A(n_8465),
.Y(n_9754)
);

OAI21xp33_ASAP7_75t_SL g9755 ( 
.A1(n_7801),
.A2(n_7300),
.B(n_6837),
.Y(n_9755)
);

INVx8_ASAP7_75t_L g9756 ( 
.A(n_8943),
.Y(n_9756)
);

INVx1_ASAP7_75t_L g9757 ( 
.A(n_8321),
.Y(n_9757)
);

NOR2xp33_ASAP7_75t_L g9758 ( 
.A(n_7866),
.B(n_7234),
.Y(n_9758)
);

INVx2_ASAP7_75t_SL g9759 ( 
.A(n_8817),
.Y(n_9759)
);

OAI21xp5_ASAP7_75t_L g9760 ( 
.A1(n_7944),
.A2(n_7432),
.B(n_7231),
.Y(n_9760)
);

NOR2xp33_ASAP7_75t_L g9761 ( 
.A(n_7866),
.B(n_7234),
.Y(n_9761)
);

AND2x2_ASAP7_75t_L g9762 ( 
.A(n_8859),
.B(n_6691),
.Y(n_9762)
);

BUFx2_ASAP7_75t_SL g9763 ( 
.A(n_7921),
.Y(n_9763)
);

BUFx2_ASAP7_75t_L g9764 ( 
.A(n_8524),
.Y(n_9764)
);

CKINVDCx20_ASAP7_75t_R g9765 ( 
.A(n_8558),
.Y(n_9765)
);

AOI21xp33_ASAP7_75t_L g9766 ( 
.A1(n_7865),
.A2(n_6776),
.B(n_7453),
.Y(n_9766)
);

AOI22xp33_ASAP7_75t_L g9767 ( 
.A1(n_7959),
.A2(n_7359),
.B1(n_7107),
.B2(n_6938),
.Y(n_9767)
);

AND2x4_ASAP7_75t_L g9768 ( 
.A(n_8074),
.B(n_6776),
.Y(n_9768)
);

AOI21xp5_ASAP7_75t_L g9769 ( 
.A1(n_8134),
.A2(n_6828),
.B(n_7233),
.Y(n_9769)
);

NOR2x1_ASAP7_75t_R g9770 ( 
.A(n_8742),
.B(n_6776),
.Y(n_9770)
);

OR2x2_ASAP7_75t_L g9771 ( 
.A(n_7986),
.B(n_6897),
.Y(n_9771)
);

INVx1_ASAP7_75t_L g9772 ( 
.A(n_8321),
.Y(n_9772)
);

BUFx3_ASAP7_75t_L g9773 ( 
.A(n_8370),
.Y(n_9773)
);

CKINVDCx20_ASAP7_75t_R g9774 ( 
.A(n_8647),
.Y(n_9774)
);

OA21x2_ASAP7_75t_L g9775 ( 
.A1(n_8289),
.A2(n_6690),
.B(n_7315),
.Y(n_9775)
);

OR2x2_ASAP7_75t_L g9776 ( 
.A(n_7986),
.B(n_6897),
.Y(n_9776)
);

AND2x4_ASAP7_75t_L g9777 ( 
.A(n_8074),
.B(n_6776),
.Y(n_9777)
);

INVx1_ASAP7_75t_L g9778 ( 
.A(n_8321),
.Y(n_9778)
);

INVx1_ASAP7_75t_L g9779 ( 
.A(n_8321),
.Y(n_9779)
);

CKINVDCx20_ASAP7_75t_R g9780 ( 
.A(n_8647),
.Y(n_9780)
);

INVx2_ASAP7_75t_SL g9781 ( 
.A(n_8817),
.Y(n_9781)
);

BUFx12f_ASAP7_75t_L g9782 ( 
.A(n_7804),
.Y(n_9782)
);

BUFx3_ASAP7_75t_L g9783 ( 
.A(n_8370),
.Y(n_9783)
);

INVx1_ASAP7_75t_L g9784 ( 
.A(n_8321),
.Y(n_9784)
);

AND2x4_ASAP7_75t_L g9785 ( 
.A(n_8074),
.B(n_6700),
.Y(n_9785)
);

OAI21xp5_ASAP7_75t_L g9786 ( 
.A1(n_7914),
.A2(n_6690),
.B(n_7315),
.Y(n_9786)
);

INVx2_ASAP7_75t_L g9787 ( 
.A(n_8292),
.Y(n_9787)
);

OAI21xp5_ASAP7_75t_L g9788 ( 
.A1(n_7914),
.A2(n_8228),
.B(n_8217),
.Y(n_9788)
);

INVx1_ASAP7_75t_L g9789 ( 
.A(n_8321),
.Y(n_9789)
);

AOI21xp5_ASAP7_75t_L g9790 ( 
.A1(n_8373),
.A2(n_6700),
.B(n_7107),
.Y(n_9790)
);

AOI21x1_ASAP7_75t_L g9791 ( 
.A1(n_8341),
.A2(n_6688),
.B(n_7231),
.Y(n_9791)
);

AND2x4_ASAP7_75t_SL g9792 ( 
.A(n_8070),
.B(n_6317),
.Y(n_9792)
);

BUFx2_ASAP7_75t_R g9793 ( 
.A(n_7804),
.Y(n_9793)
);

CKINVDCx20_ASAP7_75t_R g9794 ( 
.A(n_8706),
.Y(n_9794)
);

CKINVDCx20_ASAP7_75t_R g9795 ( 
.A(n_8706),
.Y(n_9795)
);

INVx2_ASAP7_75t_L g9796 ( 
.A(n_8292),
.Y(n_9796)
);

INVx1_ASAP7_75t_L g9797 ( 
.A(n_8054),
.Y(n_9797)
);

BUFx12f_ASAP7_75t_L g9798 ( 
.A(n_8162),
.Y(n_9798)
);

BUFx6f_ASAP7_75t_L g9799 ( 
.A(n_8625),
.Y(n_9799)
);

AOI22xp33_ASAP7_75t_L g9800 ( 
.A1(n_7959),
.A2(n_6938),
.B1(n_7359),
.B2(n_7453),
.Y(n_9800)
);

INVxp67_ASAP7_75t_SL g9801 ( 
.A(n_8933),
.Y(n_9801)
);

OAI21x1_ASAP7_75t_SL g9802 ( 
.A1(n_8531),
.A2(n_7581),
.B(n_6440),
.Y(n_9802)
);

OAI21x1_ASAP7_75t_SL g9803 ( 
.A1(n_7750),
.A2(n_7581),
.B(n_6440),
.Y(n_9803)
);

OAI21x1_ASAP7_75t_SL g9804 ( 
.A1(n_7750),
.A2(n_6440),
.B(n_6535),
.Y(n_9804)
);

HB1xp67_ASAP7_75t_L g9805 ( 
.A(n_8567),
.Y(n_9805)
);

INVx1_ASAP7_75t_SL g9806 ( 
.A(n_7757),
.Y(n_9806)
);

OAI21x1_ASAP7_75t_SL g9807 ( 
.A1(n_7750),
.A2(n_6440),
.B(n_6535),
.Y(n_9807)
);

AOI21xp5_ASAP7_75t_L g9808 ( 
.A1(n_8373),
.A2(n_6828),
.B(n_7453),
.Y(n_9808)
);

INVx2_ASAP7_75t_L g9809 ( 
.A(n_8292),
.Y(n_9809)
);

INVx1_ASAP7_75t_L g9810 ( 
.A(n_8054),
.Y(n_9810)
);

OAI21xp33_ASAP7_75t_L g9811 ( 
.A1(n_7803),
.A2(n_6767),
.B(n_7226),
.Y(n_9811)
);

OAI21x1_ASAP7_75t_L g9812 ( 
.A1(n_7794),
.A2(n_6837),
.B(n_6295),
.Y(n_9812)
);

OAI21xp5_ASAP7_75t_L g9813 ( 
.A1(n_8217),
.A2(n_6691),
.B(n_7226),
.Y(n_9813)
);

CKINVDCx5p33_ASAP7_75t_R g9814 ( 
.A(n_8742),
.Y(n_9814)
);

INVx1_ASAP7_75t_L g9815 ( 
.A(n_8054),
.Y(n_9815)
);

OAI21xp5_ASAP7_75t_SL g9816 ( 
.A1(n_7803),
.A2(n_6828),
.B(n_7321),
.Y(n_9816)
);

OAI21x1_ASAP7_75t_L g9817 ( 
.A1(n_7794),
.A2(n_6837),
.B(n_6295),
.Y(n_9817)
);

INVx1_ASAP7_75t_L g9818 ( 
.A(n_8075),
.Y(n_9818)
);

NAND2x1p5_ASAP7_75t_L g9819 ( 
.A(n_7861),
.B(n_6828),
.Y(n_9819)
);

INVx1_ASAP7_75t_L g9820 ( 
.A(n_8075),
.Y(n_9820)
);

HB1xp67_ASAP7_75t_L g9821 ( 
.A(n_8567),
.Y(n_9821)
);

NOR2xp33_ASAP7_75t_L g9822 ( 
.A(n_7931),
.B(n_6691),
.Y(n_9822)
);

AOI21xp5_ASAP7_75t_L g9823 ( 
.A1(n_8381),
.A2(n_6828),
.B(n_7359),
.Y(n_9823)
);

INVx1_ASAP7_75t_L g9824 ( 
.A(n_8075),
.Y(n_9824)
);

INVx1_ASAP7_75t_L g9825 ( 
.A(n_8227),
.Y(n_9825)
);

NAND2xp5_ASAP7_75t_L g9826 ( 
.A(n_8852),
.B(n_7204),
.Y(n_9826)
);

AND2x4_ASAP7_75t_L g9827 ( 
.A(n_8074),
.B(n_6828),
.Y(n_9827)
);

BUFx2_ASAP7_75t_SL g9828 ( 
.A(n_7921),
.Y(n_9828)
);

AND2x4_ASAP7_75t_L g9829 ( 
.A(n_8095),
.B(n_6828),
.Y(n_9829)
);

AOI22xp33_ASAP7_75t_L g9830 ( 
.A1(n_7776),
.A2(n_7107),
.B1(n_7359),
.B2(n_7321),
.Y(n_9830)
);

BUFx3_ASAP7_75t_L g9831 ( 
.A(n_8370),
.Y(n_9831)
);

INVx1_ASAP7_75t_L g9832 ( 
.A(n_8227),
.Y(n_9832)
);

AOI21x1_ASAP7_75t_L g9833 ( 
.A1(n_8341),
.A2(n_6691),
.B(n_6652),
.Y(n_9833)
);

NAND2x1p5_ASAP7_75t_L g9834 ( 
.A(n_7861),
.B(n_7321),
.Y(n_9834)
);

AND2x6_ASAP7_75t_L g9835 ( 
.A(n_7752),
.B(n_7321),
.Y(n_9835)
);

BUFx6f_ASAP7_75t_L g9836 ( 
.A(n_8625),
.Y(n_9836)
);

NAND2x1_ASAP7_75t_L g9837 ( 
.A(n_8029),
.B(n_7437),
.Y(n_9837)
);

BUFx6f_ASAP7_75t_L g9838 ( 
.A(n_8171),
.Y(n_9838)
);

INVx1_ASAP7_75t_L g9839 ( 
.A(n_8227),
.Y(n_9839)
);

INVx1_ASAP7_75t_L g9840 ( 
.A(n_8245),
.Y(n_9840)
);

INVx6_ASAP7_75t_L g9841 ( 
.A(n_7735),
.Y(n_9841)
);

NAND2xp5_ASAP7_75t_L g9842 ( 
.A(n_8852),
.B(n_7602),
.Y(n_9842)
);

INVx2_ASAP7_75t_L g9843 ( 
.A(n_8292),
.Y(n_9843)
);

INVx1_ASAP7_75t_SL g9844 ( 
.A(n_7757),
.Y(n_9844)
);

INVx3_ASAP7_75t_L g9845 ( 
.A(n_8804),
.Y(n_9845)
);

INVx1_ASAP7_75t_L g9846 ( 
.A(n_8245),
.Y(n_9846)
);

BUFx12f_ASAP7_75t_L g9847 ( 
.A(n_8162),
.Y(n_9847)
);

AOI22x1_ASAP7_75t_L g9848 ( 
.A1(n_7902),
.A2(n_7107),
.B1(n_7359),
.B2(n_7321),
.Y(n_9848)
);

INVx3_ASAP7_75t_L g9849 ( 
.A(n_8804),
.Y(n_9849)
);

NOR2xp33_ASAP7_75t_L g9850 ( 
.A(n_7931),
.B(n_6692),
.Y(n_9850)
);

INVx2_ASAP7_75t_SL g9851 ( 
.A(n_8817),
.Y(n_9851)
);

OAI21xp5_ASAP7_75t_L g9852 ( 
.A1(n_8228),
.A2(n_6652),
.B(n_6692),
.Y(n_9852)
);

INVx1_ASAP7_75t_L g9853 ( 
.A(n_8245),
.Y(n_9853)
);

NOR2xp33_ASAP7_75t_L g9854 ( 
.A(n_8064),
.B(n_7226),
.Y(n_9854)
);

INVx4_ASAP7_75t_L g9855 ( 
.A(n_8070),
.Y(n_9855)
);

INVxp67_ASAP7_75t_L g9856 ( 
.A(n_7840),
.Y(n_9856)
);

HB1xp67_ASAP7_75t_L g9857 ( 
.A(n_8567),
.Y(n_9857)
);

AND2x4_ASAP7_75t_L g9858 ( 
.A(n_8095),
.B(n_6700),
.Y(n_9858)
);

INVx2_ASAP7_75t_L g9859 ( 
.A(n_8292),
.Y(n_9859)
);

INVx2_ASAP7_75t_SL g9860 ( 
.A(n_8817),
.Y(n_9860)
);

AOI21xp5_ASAP7_75t_L g9861 ( 
.A1(n_8381),
.A2(n_6700),
.B(n_6677),
.Y(n_9861)
);

INVx2_ASAP7_75t_L g9862 ( 
.A(n_8292),
.Y(n_9862)
);

AO21x2_ASAP7_75t_L g9863 ( 
.A1(n_8487),
.A2(n_6652),
.B(n_7226),
.Y(n_9863)
);

INVx2_ASAP7_75t_L g9864 ( 
.A(n_8292),
.Y(n_9864)
);

INVx3_ASAP7_75t_L g9865 ( 
.A(n_8804),
.Y(n_9865)
);

INVx1_ASAP7_75t_SL g9866 ( 
.A(n_7757),
.Y(n_9866)
);

HB1xp67_ASAP7_75t_L g9867 ( 
.A(n_8567),
.Y(n_9867)
);

NOR2xp33_ASAP7_75t_L g9868 ( 
.A(n_8064),
.B(n_8192),
.Y(n_9868)
);

INVx5_ASAP7_75t_L g9869 ( 
.A(n_7744),
.Y(n_9869)
);

NAND2x1_ASAP7_75t_L g9870 ( 
.A(n_8431),
.B(n_6677),
.Y(n_9870)
);

AO21x1_ASAP7_75t_L g9871 ( 
.A1(n_7919),
.A2(n_6440),
.B(n_6677),
.Y(n_9871)
);

BUFx6f_ASAP7_75t_L g9872 ( 
.A(n_8171),
.Y(n_9872)
);

INVx4_ASAP7_75t_L g9873 ( 
.A(n_8165),
.Y(n_9873)
);

INVx4_ASAP7_75t_L g9874 ( 
.A(n_8165),
.Y(n_9874)
);

HB1xp67_ASAP7_75t_L g9875 ( 
.A(n_8567),
.Y(n_9875)
);

AND2x2_ASAP7_75t_L g9876 ( 
.A(n_8859),
.B(n_6440),
.Y(n_9876)
);

INVx1_ASAP7_75t_L g9877 ( 
.A(n_8252),
.Y(n_9877)
);

INVx1_ASAP7_75t_L g9878 ( 
.A(n_8252),
.Y(n_9878)
);

NOR2xp33_ASAP7_75t_L g9879 ( 
.A(n_8064),
.B(n_6440),
.Y(n_9879)
);

AND2x2_ASAP7_75t_L g9880 ( 
.A(n_8859),
.B(n_6440),
.Y(n_9880)
);

AOI21xp5_ASAP7_75t_L g9881 ( 
.A1(n_7851),
.A2(n_6535),
.B(n_7807),
.Y(n_9881)
);

OAI21xp5_ASAP7_75t_L g9882 ( 
.A1(n_8012),
.A2(n_6535),
.B(n_8081),
.Y(n_9882)
);

AND2x4_ASAP7_75t_L g9883 ( 
.A(n_8095),
.B(n_6535),
.Y(n_9883)
);

CKINVDCx20_ASAP7_75t_R g9884 ( 
.A(n_8720),
.Y(n_9884)
);

HB1xp67_ASAP7_75t_L g9885 ( 
.A(n_8567),
.Y(n_9885)
);

OAI21x1_ASAP7_75t_L g9886 ( 
.A1(n_7822),
.A2(n_6535),
.B(n_7835),
.Y(n_9886)
);

OAI21xp5_ASAP7_75t_L g9887 ( 
.A1(n_8012),
.A2(n_6535),
.B(n_8201),
.Y(n_9887)
);

BUFx12f_ASAP7_75t_L g9888 ( 
.A(n_8162),
.Y(n_9888)
);

OR2x2_ASAP7_75t_L g9889 ( 
.A(n_7986),
.B(n_7954),
.Y(n_9889)
);

BUFx2_ASAP7_75t_L g9890 ( 
.A(n_8524),
.Y(n_9890)
);

INVx2_ASAP7_75t_SL g9891 ( 
.A(n_8817),
.Y(n_9891)
);

BUFx6f_ASAP7_75t_L g9892 ( 
.A(n_8171),
.Y(n_9892)
);

OAI21x1_ASAP7_75t_L g9893 ( 
.A1(n_7822),
.A2(n_7850),
.B(n_7835),
.Y(n_9893)
);

AND2x2_ASAP7_75t_L g9894 ( 
.A(n_8718),
.B(n_8755),
.Y(n_9894)
);

OAI21x1_ASAP7_75t_L g9895 ( 
.A1(n_7822),
.A2(n_7850),
.B(n_7835),
.Y(n_9895)
);

OAI21x1_ASAP7_75t_L g9896 ( 
.A1(n_7850),
.A2(n_7859),
.B(n_7855),
.Y(n_9896)
);

O2A1O1Ixp33_ASAP7_75t_L g9897 ( 
.A1(n_7911),
.A2(n_8107),
.B(n_7776),
.C(n_8169),
.Y(n_9897)
);

AOI21xp33_ASAP7_75t_L g9898 ( 
.A1(n_7776),
.A2(n_7985),
.B(n_7807),
.Y(n_9898)
);

OAI21x1_ASAP7_75t_L g9899 ( 
.A1(n_7850),
.A2(n_7859),
.B(n_7855),
.Y(n_9899)
);

OR2x6_ASAP7_75t_L g9900 ( 
.A(n_8021),
.B(n_8369),
.Y(n_9900)
);

AO31x2_ASAP7_75t_L g9901 ( 
.A1(n_8133),
.A2(n_8031),
.A3(n_8157),
.B(n_8659),
.Y(n_9901)
);

AO21x2_ASAP7_75t_L g9902 ( 
.A1(n_8487),
.A2(n_8065),
.B(n_8057),
.Y(n_9902)
);

INVx1_ASAP7_75t_L g9903 ( 
.A(n_8252),
.Y(n_9903)
);

OAI21xp5_ASAP7_75t_L g9904 ( 
.A1(n_8012),
.A2(n_8201),
.B(n_8126),
.Y(n_9904)
);

INVxp67_ASAP7_75t_L g9905 ( 
.A(n_7840),
.Y(n_9905)
);

NAND2xp5_ASAP7_75t_L g9906 ( 
.A(n_8866),
.B(n_8362),
.Y(n_9906)
);

OAI21x1_ASAP7_75t_L g9907 ( 
.A1(n_7868),
.A2(n_7878),
.B(n_7877),
.Y(n_9907)
);

AND2x4_ASAP7_75t_L g9908 ( 
.A(n_8095),
.B(n_8207),
.Y(n_9908)
);

OA21x2_ASAP7_75t_L g9909 ( 
.A1(n_8562),
.A2(n_8654),
.B(n_8556),
.Y(n_9909)
);

CKINVDCx12_ASAP7_75t_R g9910 ( 
.A(n_7808),
.Y(n_9910)
);

BUFx6f_ASAP7_75t_L g9911 ( 
.A(n_8171),
.Y(n_9911)
);

INVx1_ASAP7_75t_L g9912 ( 
.A(n_8280),
.Y(n_9912)
);

OAI21x1_ASAP7_75t_L g9913 ( 
.A1(n_7868),
.A2(n_7878),
.B(n_7877),
.Y(n_9913)
);

INVx2_ASAP7_75t_L g9914 ( 
.A(n_8292),
.Y(n_9914)
);

AND2x4_ASAP7_75t_L g9915 ( 
.A(n_8095),
.B(n_8207),
.Y(n_9915)
);

OA21x2_ASAP7_75t_L g9916 ( 
.A1(n_8654),
.A2(n_8556),
.B(n_8598),
.Y(n_9916)
);

INVx1_ASAP7_75t_L g9917 ( 
.A(n_8280),
.Y(n_9917)
);

BUFx3_ASAP7_75t_L g9918 ( 
.A(n_8828),
.Y(n_9918)
);

AND2x2_ASAP7_75t_L g9919 ( 
.A(n_8718),
.B(n_8755),
.Y(n_9919)
);

INVx2_ASAP7_75t_L g9920 ( 
.A(n_8292),
.Y(n_9920)
);

NAND2xp5_ASAP7_75t_L g9921 ( 
.A(n_8866),
.B(n_8362),
.Y(n_9921)
);

OAI21xp5_ASAP7_75t_L g9922 ( 
.A1(n_8126),
.A2(n_7969),
.B(n_8083),
.Y(n_9922)
);

INVxp67_ASAP7_75t_L g9923 ( 
.A(n_7840),
.Y(n_9923)
);

NAND2x1p5_ASAP7_75t_L g9924 ( 
.A(n_7861),
.B(n_7901),
.Y(n_9924)
);

OA21x2_ASAP7_75t_L g9925 ( 
.A1(n_8654),
.A2(n_8556),
.B(n_8598),
.Y(n_9925)
);

OAI21x1_ASAP7_75t_L g9926 ( 
.A1(n_7877),
.A2(n_7888),
.B(n_7878),
.Y(n_9926)
);

AO21x2_ASAP7_75t_L g9927 ( 
.A1(n_8057),
.A2(n_8065),
.B(n_8705),
.Y(n_9927)
);

OAI21x1_ASAP7_75t_L g9928 ( 
.A1(n_7877),
.A2(n_7888),
.B(n_7878),
.Y(n_9928)
);

OAI21x1_ASAP7_75t_L g9929 ( 
.A1(n_7888),
.A2(n_7896),
.B(n_7890),
.Y(n_9929)
);

OAI21x1_ASAP7_75t_L g9930 ( 
.A1(n_7888),
.A2(n_7896),
.B(n_7890),
.Y(n_9930)
);

HB1xp67_ASAP7_75t_L g9931 ( 
.A(n_8567),
.Y(n_9931)
);

NAND2xp5_ASAP7_75t_L g9932 ( 
.A(n_8366),
.B(n_8383),
.Y(n_9932)
);

CKINVDCx5p33_ASAP7_75t_R g9933 ( 
.A(n_8742),
.Y(n_9933)
);

AND2x4_ASAP7_75t_L g9934 ( 
.A(n_8095),
.B(n_8207),
.Y(n_9934)
);

INVx1_ASAP7_75t_L g9935 ( 
.A(n_8280),
.Y(n_9935)
);

AO21x2_ASAP7_75t_L g9936 ( 
.A1(n_8705),
.A2(n_8753),
.B(n_7851),
.Y(n_9936)
);

AO21x2_ASAP7_75t_L g9937 ( 
.A1(n_8753),
.A2(n_8283),
.B(n_7988),
.Y(n_9937)
);

HB1xp67_ASAP7_75t_L g9938 ( 
.A(n_8567),
.Y(n_9938)
);

INVx1_ASAP7_75t_L g9939 ( 
.A(n_7984),
.Y(n_9939)
);

HB1xp67_ASAP7_75t_L g9940 ( 
.A(n_8567),
.Y(n_9940)
);

BUFx6f_ASAP7_75t_L g9941 ( 
.A(n_8171),
.Y(n_9941)
);

OAI21xp5_ASAP7_75t_L g9942 ( 
.A1(n_8126),
.A2(n_7969),
.B(n_8083),
.Y(n_9942)
);

INVx1_ASAP7_75t_L g9943 ( 
.A(n_7984),
.Y(n_9943)
);

AO21x2_ASAP7_75t_L g9944 ( 
.A1(n_8283),
.A2(n_7988),
.B(n_8316),
.Y(n_9944)
);

HB1xp67_ASAP7_75t_L g9945 ( 
.A(n_8585),
.Y(n_9945)
);

BUFx3_ASAP7_75t_L g9946 ( 
.A(n_8828),
.Y(n_9946)
);

INVx3_ASAP7_75t_L g9947 ( 
.A(n_8804),
.Y(n_9947)
);

OAI21xp5_ASAP7_75t_L g9948 ( 
.A1(n_7985),
.A2(n_8107),
.B(n_8234),
.Y(n_9948)
);

INVx1_ASAP7_75t_L g9949 ( 
.A(n_7984),
.Y(n_9949)
);

NAND3xp33_ASAP7_75t_L g9950 ( 
.A(n_7998),
.B(n_7956),
.C(n_8048),
.Y(n_9950)
);

OAI21x1_ASAP7_75t_L g9951 ( 
.A1(n_7890),
.A2(n_7900),
.B(n_7896),
.Y(n_9951)
);

OAI21x1_ASAP7_75t_SL g9952 ( 
.A1(n_7867),
.A2(n_8041),
.B(n_8018),
.Y(n_9952)
);

AO21x2_ASAP7_75t_L g9953 ( 
.A1(n_8316),
.A2(n_7875),
.B(n_8235),
.Y(n_9953)
);

BUFx6f_ASAP7_75t_L g9954 ( 
.A(n_8171),
.Y(n_9954)
);

INVx1_ASAP7_75t_L g9955 ( 
.A(n_8444),
.Y(n_9955)
);

INVx2_ASAP7_75t_SL g9956 ( 
.A(n_8817),
.Y(n_9956)
);

AO21x2_ASAP7_75t_L g9957 ( 
.A1(n_7875),
.A2(n_8235),
.B(n_8801),
.Y(n_9957)
);

OAI21x1_ASAP7_75t_L g9958 ( 
.A1(n_7890),
.A2(n_7900),
.B(n_7896),
.Y(n_9958)
);

AND2x2_ASAP7_75t_SL g9959 ( 
.A(n_7883),
.B(n_8035),
.Y(n_9959)
);

NOR2xp33_ASAP7_75t_SL g9960 ( 
.A(n_7741),
.B(n_8031),
.Y(n_9960)
);

OAI21x1_ASAP7_75t_L g9961 ( 
.A1(n_7900),
.A2(n_7790),
.B(n_7788),
.Y(n_9961)
);

NOR2xp33_ASAP7_75t_L g9962 ( 
.A(n_8192),
.B(n_8016),
.Y(n_9962)
);

INVx1_ASAP7_75t_L g9963 ( 
.A(n_8444),
.Y(n_9963)
);

OAI21x1_ASAP7_75t_L g9964 ( 
.A1(n_7900),
.A2(n_7790),
.B(n_7788),
.Y(n_9964)
);

BUFx5_ASAP7_75t_L g9965 ( 
.A(n_8768),
.Y(n_9965)
);

OAI21xp33_ASAP7_75t_L g9966 ( 
.A1(n_7956),
.A2(n_8619),
.B(n_7839),
.Y(n_9966)
);

BUFx6f_ASAP7_75t_L g9967 ( 
.A(n_8171),
.Y(n_9967)
);

BUFx12f_ASAP7_75t_L g9968 ( 
.A(n_8162),
.Y(n_9968)
);

OAI21xp5_ASAP7_75t_L g9969 ( 
.A1(n_8234),
.A2(n_7919),
.B(n_7998),
.Y(n_9969)
);

NOR2xp33_ASAP7_75t_L g9970 ( 
.A(n_8016),
.B(n_8619),
.Y(n_9970)
);

OA21x2_ASAP7_75t_L g9971 ( 
.A1(n_8556),
.A2(n_8604),
.B(n_8602),
.Y(n_9971)
);

OR2x2_ASAP7_75t_L g9972 ( 
.A(n_7986),
.B(n_7954),
.Y(n_9972)
);

OAI21x1_ASAP7_75t_L g9973 ( 
.A1(n_8195),
.A2(n_8578),
.B(n_8572),
.Y(n_9973)
);

AND2x4_ASAP7_75t_L g9974 ( 
.A(n_8207),
.B(n_7921),
.Y(n_9974)
);

INVx6_ASAP7_75t_SL g9975 ( 
.A(n_8021),
.Y(n_9975)
);

OAI21x1_ASAP7_75t_SL g9976 ( 
.A1(n_7867),
.A2(n_8041),
.B(n_8018),
.Y(n_9976)
);

INVx1_ASAP7_75t_L g9977 ( 
.A(n_8444),
.Y(n_9977)
);

AO21x2_ASAP7_75t_L g9978 ( 
.A1(n_7875),
.A2(n_8801),
.B(n_7925),
.Y(n_9978)
);

INVx1_ASAP7_75t_L g9979 ( 
.A(n_8451),
.Y(n_9979)
);

INVx1_ASAP7_75t_L g9980 ( 
.A(n_8451),
.Y(n_9980)
);

OA21x2_ASAP7_75t_L g9981 ( 
.A1(n_8602),
.A2(n_8604),
.B(n_8578),
.Y(n_9981)
);

BUFx3_ASAP7_75t_L g9982 ( 
.A(n_8828),
.Y(n_9982)
);

INVx2_ASAP7_75t_L g9983 ( 
.A(n_8399),
.Y(n_9983)
);

BUFx12f_ASAP7_75t_L g9984 ( 
.A(n_8282),
.Y(n_9984)
);

OAI21x1_ASAP7_75t_L g9985 ( 
.A1(n_8195),
.A2(n_8578),
.B(n_8572),
.Y(n_9985)
);

AO21x2_ASAP7_75t_L g9986 ( 
.A1(n_7875),
.A2(n_8801),
.B(n_7925),
.Y(n_9986)
);

NAND2xp5_ASAP7_75t_L g9987 ( 
.A(n_8366),
.B(n_8383),
.Y(n_9987)
);

INVx1_ASAP7_75t_L g9988 ( 
.A(n_8451),
.Y(n_9988)
);

INVx4_ASAP7_75t_L g9989 ( 
.A(n_8165),
.Y(n_9989)
);

BUFx3_ASAP7_75t_L g9990 ( 
.A(n_8837),
.Y(n_9990)
);

OAI21x1_ASAP7_75t_L g9991 ( 
.A1(n_8572),
.A2(n_8578),
.B(n_8847),
.Y(n_9991)
);

INVx1_ASAP7_75t_L g9992 ( 
.A(n_8451),
.Y(n_9992)
);

INVx2_ASAP7_75t_SL g9993 ( 
.A(n_8103),
.Y(n_9993)
);

NAND2x1p5_ASAP7_75t_L g9994 ( 
.A(n_7861),
.B(n_7901),
.Y(n_9994)
);

AOI21xp5_ASAP7_75t_L g9995 ( 
.A1(n_8326),
.A2(n_8155),
.B(n_8175),
.Y(n_9995)
);

AND2x2_ASAP7_75t_L g9996 ( 
.A(n_8718),
.B(n_8755),
.Y(n_9996)
);

INVx6_ASAP7_75t_L g9997 ( 
.A(n_7735),
.Y(n_9997)
);

OAI21xp33_ASAP7_75t_L g9998 ( 
.A1(n_7956),
.A2(n_7839),
.B(n_7791),
.Y(n_9998)
);

INVx2_ASAP7_75t_L g9999 ( 
.A(n_8399),
.Y(n_9999)
);

OAI21x1_ASAP7_75t_L g10000 ( 
.A1(n_8856),
.A2(n_8863),
.B(n_8883),
.Y(n_10000)
);

OAI21x1_ASAP7_75t_L g10001 ( 
.A1(n_8863),
.A2(n_8896),
.B(n_8883),
.Y(n_10001)
);

OR2x6_ASAP7_75t_L g10002 ( 
.A(n_8021),
.B(n_8369),
.Y(n_10002)
);

HB1xp67_ASAP7_75t_L g10003 ( 
.A(n_8585),
.Y(n_10003)
);

BUFx3_ASAP7_75t_L g10004 ( 
.A(n_8837),
.Y(n_10004)
);

AOI22xp33_ASAP7_75t_L g10005 ( 
.A1(n_8708),
.A2(n_7801),
.B1(n_8076),
.B2(n_7965),
.Y(n_10005)
);

BUFx2_ASAP7_75t_SL g10006 ( 
.A(n_7960),
.Y(n_10006)
);

OA21x2_ASAP7_75t_L g10007 ( 
.A1(n_8787),
.A2(n_8809),
.B(n_8807),
.Y(n_10007)
);

INVx1_ASAP7_75t_L g10008 ( 
.A(n_8451),
.Y(n_10008)
);

OAI21x1_ASAP7_75t_SL g10009 ( 
.A1(n_7867),
.A2(n_8041),
.B(n_8018),
.Y(n_10009)
);

AO21x2_ASAP7_75t_L g10010 ( 
.A1(n_7875),
.A2(n_8290),
.B(n_8079),
.Y(n_10010)
);

NAND2x1p5_ASAP7_75t_L g10011 ( 
.A(n_7901),
.B(n_8103),
.Y(n_10011)
);

INVx4_ASAP7_75t_L g10012 ( 
.A(n_8165),
.Y(n_10012)
);

AO21x2_ASAP7_75t_L g10013 ( 
.A1(n_7875),
.A2(n_8290),
.B(n_8079),
.Y(n_10013)
);

OAI21x1_ASAP7_75t_L g10014 ( 
.A1(n_8883),
.A2(n_8898),
.B(n_8896),
.Y(n_10014)
);

OAI21x1_ASAP7_75t_L g10015 ( 
.A1(n_8883),
.A2(n_8898),
.B(n_8896),
.Y(n_10015)
);

OAI21x1_ASAP7_75t_L g10016 ( 
.A1(n_8896),
.A2(n_8901),
.B(n_8898),
.Y(n_10016)
);

CKINVDCx20_ASAP7_75t_R g10017 ( 
.A(n_8720),
.Y(n_10017)
);

AO21x2_ASAP7_75t_L g10018 ( 
.A1(n_8419),
.A2(n_8375),
.B(n_8086),
.Y(n_10018)
);

INVx1_ASAP7_75t_SL g10019 ( 
.A(n_7757),
.Y(n_10019)
);

OAI21xp5_ASAP7_75t_L g10020 ( 
.A1(n_8234),
.A2(n_8169),
.B(n_8048),
.Y(n_10020)
);

NAND2xp5_ASAP7_75t_L g10021 ( 
.A(n_8733),
.B(n_8743),
.Y(n_10021)
);

INVx2_ASAP7_75t_L g10022 ( 
.A(n_8399),
.Y(n_10022)
);

INVx2_ASAP7_75t_SL g10023 ( 
.A(n_8103),
.Y(n_10023)
);

BUFx6f_ASAP7_75t_L g10024 ( 
.A(n_8171),
.Y(n_10024)
);

AOI22xp33_ASAP7_75t_L g10025 ( 
.A1(n_8708),
.A2(n_7801),
.B1(n_8076),
.B2(n_7965),
.Y(n_10025)
);

OA21x2_ASAP7_75t_L g10026 ( 
.A1(n_8787),
.A2(n_8809),
.B(n_8807),
.Y(n_10026)
);

INVx8_ASAP7_75t_L g10027 ( 
.A(n_8943),
.Y(n_10027)
);

INVx1_ASAP7_75t_L g10028 ( 
.A(n_8451),
.Y(n_10028)
);

INVx2_ASAP7_75t_L g10029 ( 
.A(n_8399),
.Y(n_10029)
);

INVx1_ASAP7_75t_L g10030 ( 
.A(n_8451),
.Y(n_10030)
);

OR2x2_ASAP7_75t_L g10031 ( 
.A(n_7986),
.B(n_7954),
.Y(n_10031)
);

INVx5_ASAP7_75t_L g10032 ( 
.A(n_7744),
.Y(n_10032)
);

BUFx6f_ASAP7_75t_L g10033 ( 
.A(n_8171),
.Y(n_10033)
);

AND2x4_ASAP7_75t_L g10034 ( 
.A(n_8207),
.B(n_7960),
.Y(n_10034)
);

INVx1_ASAP7_75t_L g10035 ( 
.A(n_8451),
.Y(n_10035)
);

BUFx6f_ASAP7_75t_L g10036 ( 
.A(n_8689),
.Y(n_10036)
);

NAND2xp5_ASAP7_75t_L g10037 ( 
.A(n_8733),
.B(n_8743),
.Y(n_10037)
);

NAND2x1p5_ASAP7_75t_L g10038 ( 
.A(n_7901),
.B(n_8103),
.Y(n_10038)
);

OA21x2_ASAP7_75t_L g10039 ( 
.A1(n_8844),
.A2(n_8890),
.B(n_8889),
.Y(n_10039)
);

INVx2_ASAP7_75t_L g10040 ( 
.A(n_8399),
.Y(n_10040)
);

BUFx2_ASAP7_75t_R g10041 ( 
.A(n_8222),
.Y(n_10041)
);

AOI21xp5_ASAP7_75t_L g10042 ( 
.A1(n_8326),
.A2(n_8155),
.B(n_8175),
.Y(n_10042)
);

NOR2x1_ASAP7_75t_SL g10043 ( 
.A(n_8165),
.B(n_8208),
.Y(n_10043)
);

AOI21xp5_ASAP7_75t_L g10044 ( 
.A1(n_8310),
.A2(n_8320),
.B(n_8324),
.Y(n_10044)
);

NOR2xp33_ASAP7_75t_L g10045 ( 
.A(n_7858),
.B(n_7801),
.Y(n_10045)
);

INVx1_ASAP7_75t_L g10046 ( 
.A(n_8451),
.Y(n_10046)
);

NAND2x1p5_ASAP7_75t_L g10047 ( 
.A(n_7901),
.B(n_8103),
.Y(n_10047)
);

BUFx6f_ASAP7_75t_L g10048 ( 
.A(n_8689),
.Y(n_10048)
);

INVx4_ASAP7_75t_L g10049 ( 
.A(n_8165),
.Y(n_10049)
);

INVx1_ASAP7_75t_L g10050 ( 
.A(n_8483),
.Y(n_10050)
);

INVx5_ASAP7_75t_L g10051 ( 
.A(n_7744),
.Y(n_10051)
);

AND2x2_ASAP7_75t_L g10052 ( 
.A(n_8718),
.B(n_8755),
.Y(n_10052)
);

INVx5_ASAP7_75t_SL g10053 ( 
.A(n_7744),
.Y(n_10053)
);

OAI21x1_ASAP7_75t_SL g10054 ( 
.A1(n_8431),
.A2(n_7710),
.B(n_8032),
.Y(n_10054)
);

OA21x2_ASAP7_75t_L g10055 ( 
.A1(n_8844),
.A2(n_8890),
.B(n_8889),
.Y(n_10055)
);

BUFx3_ASAP7_75t_L g10056 ( 
.A(n_8837),
.Y(n_10056)
);

INVx1_ASAP7_75t_L g10057 ( 
.A(n_8483),
.Y(n_10057)
);

AOI22x1_ASAP7_75t_L g10058 ( 
.A1(n_8042),
.A2(n_8408),
.B1(n_8071),
.B2(n_8404),
.Y(n_10058)
);

AND2x4_ASAP7_75t_L g10059 ( 
.A(n_8207),
.B(n_7960),
.Y(n_10059)
);

OAI21xp5_ASAP7_75t_L g10060 ( 
.A1(n_8266),
.A2(n_8256),
.B(n_7764),
.Y(n_10060)
);

INVx2_ASAP7_75t_L g10061 ( 
.A(n_8399),
.Y(n_10061)
);

OAI21x1_ASAP7_75t_L g10062 ( 
.A1(n_7940),
.A2(n_7946),
.B(n_7945),
.Y(n_10062)
);

BUFx3_ASAP7_75t_L g10063 ( 
.A(n_8103),
.Y(n_10063)
);

INVx1_ASAP7_75t_L g10064 ( 
.A(n_8483),
.Y(n_10064)
);

BUFx2_ASAP7_75t_L g10065 ( 
.A(n_8689),
.Y(n_10065)
);

NAND2xp5_ASAP7_75t_L g10066 ( 
.A(n_8747),
.B(n_8386),
.Y(n_10066)
);

INVx2_ASAP7_75t_L g10067 ( 
.A(n_8399),
.Y(n_10067)
);

NOR2xp33_ASAP7_75t_L g10068 ( 
.A(n_7858),
.B(n_7801),
.Y(n_10068)
);

INVx1_ASAP7_75t_L g10069 ( 
.A(n_8483),
.Y(n_10069)
);

AO21x2_ASAP7_75t_L g10070 ( 
.A1(n_8419),
.A2(n_8375),
.B(n_8086),
.Y(n_10070)
);

AOI22xp5_ASAP7_75t_L g10071 ( 
.A1(n_7791),
.A2(n_8084),
.B1(n_8167),
.B2(n_8140),
.Y(n_10071)
);

AOI21xp5_ASAP7_75t_L g10072 ( 
.A1(n_8310),
.A2(n_8320),
.B(n_8324),
.Y(n_10072)
);

OR2x2_ASAP7_75t_L g10073 ( 
.A(n_7986),
.B(n_7954),
.Y(n_10073)
);

NAND2xp5_ASAP7_75t_L g10074 ( 
.A(n_8747),
.B(n_8386),
.Y(n_10074)
);

INVx1_ASAP7_75t_L g10075 ( 
.A(n_8483),
.Y(n_10075)
);

INVx1_ASAP7_75t_SL g10076 ( 
.A(n_8862),
.Y(n_10076)
);

INVx1_ASAP7_75t_SL g10077 ( 
.A(n_8862),
.Y(n_10077)
);

OA21x2_ASAP7_75t_L g10078 ( 
.A1(n_8909),
.A2(n_8910),
.B(n_8785),
.Y(n_10078)
);

BUFx4f_ASAP7_75t_L g10079 ( 
.A(n_8165),
.Y(n_10079)
);

INVx2_ASAP7_75t_L g10080 ( 
.A(n_8399),
.Y(n_10080)
);

INVx2_ASAP7_75t_SL g10081 ( 
.A(n_8103),
.Y(n_10081)
);

NOR2xp33_ASAP7_75t_L g10082 ( 
.A(n_7858),
.B(n_7823),
.Y(n_10082)
);

AND2x2_ASAP7_75t_L g10083 ( 
.A(n_8756),
.B(n_7894),
.Y(n_10083)
);

AND2x4_ASAP7_75t_L g10084 ( 
.A(n_8027),
.B(n_8860),
.Y(n_10084)
);

INVx1_ASAP7_75t_L g10085 ( 
.A(n_8483),
.Y(n_10085)
);

BUFx12f_ASAP7_75t_L g10086 ( 
.A(n_8282),
.Y(n_10086)
);

OAI21x1_ASAP7_75t_L g10087 ( 
.A1(n_7979),
.A2(n_8882),
.B(n_8873),
.Y(n_10087)
);

BUFx2_ASAP7_75t_R g10088 ( 
.A(n_8222),
.Y(n_10088)
);

O2A1O1Ixp33_ASAP7_75t_L g10089 ( 
.A1(n_7911),
.A2(n_8024),
.B(n_8042),
.C(n_8167),
.Y(n_10089)
);

CKINVDCx5p33_ASAP7_75t_R g10090 ( 
.A(n_8742),
.Y(n_10090)
);

INVx6_ASAP7_75t_L g10091 ( 
.A(n_7735),
.Y(n_10091)
);

OAI22xp5_ASAP7_75t_L g10092 ( 
.A1(n_7827),
.A2(n_8040),
.B1(n_7893),
.B2(n_8140),
.Y(n_10092)
);

OAI21x1_ASAP7_75t_SL g10093 ( 
.A1(n_8431),
.A2(n_7710),
.B(n_8032),
.Y(n_10093)
);

OA21x2_ASAP7_75t_L g10094 ( 
.A1(n_8909),
.A2(n_8910),
.B(n_8785),
.Y(n_10094)
);

INVx1_ASAP7_75t_L g10095 ( 
.A(n_8483),
.Y(n_10095)
);

INVxp67_ASAP7_75t_L g10096 ( 
.A(n_8170),
.Y(n_10096)
);

AO21x2_ASAP7_75t_L g10097 ( 
.A1(n_8686),
.A2(n_8693),
.B(n_8193),
.Y(n_10097)
);

OAI21x1_ASAP7_75t_L g10098 ( 
.A1(n_8873),
.A2(n_8905),
.B(n_8882),
.Y(n_10098)
);

OAI21xp5_ASAP7_75t_L g10099 ( 
.A1(n_8266),
.A2(n_8256),
.B(n_7764),
.Y(n_10099)
);

INVx6_ASAP7_75t_L g10100 ( 
.A(n_7735),
.Y(n_10100)
);

OAI21xp5_ASAP7_75t_L g10101 ( 
.A1(n_8395),
.A2(n_8193),
.B(n_8013),
.Y(n_10101)
);

AND2x4_ASAP7_75t_L g10102 ( 
.A(n_8027),
.B(n_8860),
.Y(n_10102)
);

OR2x6_ASAP7_75t_L g10103 ( 
.A(n_8021),
.B(n_8369),
.Y(n_10103)
);

NAND2x1p5_ASAP7_75t_L g10104 ( 
.A(n_7901),
.B(n_8103),
.Y(n_10104)
);

AOI22x1_ASAP7_75t_L g10105 ( 
.A1(n_8408),
.A2(n_8071),
.B1(n_8404),
.B2(n_8180),
.Y(n_10105)
);

INVx4_ASAP7_75t_L g10106 ( 
.A(n_8165),
.Y(n_10106)
);

INVx1_ASAP7_75t_L g10107 ( 
.A(n_8483),
.Y(n_10107)
);

OAI21x1_ASAP7_75t_L g10108 ( 
.A1(n_8882),
.A2(n_8918),
.B(n_8905),
.Y(n_10108)
);

AOI22xp5_ASAP7_75t_L g10109 ( 
.A1(n_8084),
.A2(n_8295),
.B1(n_8111),
.B2(n_7943),
.Y(n_10109)
);

BUFx6f_ASAP7_75t_L g10110 ( 
.A(n_8689),
.Y(n_10110)
);

AO21x2_ASAP7_75t_L g10111 ( 
.A1(n_8686),
.A2(n_8693),
.B(n_8432),
.Y(n_10111)
);

INVx2_ASAP7_75t_SL g10112 ( 
.A(n_8103),
.Y(n_10112)
);

NAND2xp5_ASAP7_75t_L g10113 ( 
.A(n_8390),
.B(n_8118),
.Y(n_10113)
);

AOI21xp5_ASAP7_75t_L g10114 ( 
.A1(n_8577),
.A2(n_8541),
.B(n_8024),
.Y(n_10114)
);

AO31x2_ASAP7_75t_L g10115 ( 
.A1(n_8157),
.A2(n_8659),
.A3(n_8669),
.B(n_8040),
.Y(n_10115)
);

BUFx4f_ASAP7_75t_SL g10116 ( 
.A(n_8078),
.Y(n_10116)
);

AO21x2_ASAP7_75t_L g10117 ( 
.A1(n_8432),
.A2(n_8668),
.B(n_8635),
.Y(n_10117)
);

OA21x2_ASAP7_75t_L g10118 ( 
.A1(n_8784),
.A2(n_8731),
.B(n_8668),
.Y(n_10118)
);

OAI21x1_ASAP7_75t_L g10119 ( 
.A1(n_8882),
.A2(n_8918),
.B(n_8905),
.Y(n_10119)
);

OAI21x1_ASAP7_75t_L g10120 ( 
.A1(n_8905),
.A2(n_8918),
.B(n_8426),
.Y(n_10120)
);

OR2x6_ASAP7_75t_L g10121 ( 
.A(n_8369),
.B(n_7744),
.Y(n_10121)
);

OAI21x1_ASAP7_75t_L g10122 ( 
.A1(n_8918),
.A2(n_8426),
.B(n_8631),
.Y(n_10122)
);

INVx1_ASAP7_75t_L g10123 ( 
.A(n_8483),
.Y(n_10123)
);

AO21x2_ASAP7_75t_L g10124 ( 
.A1(n_8635),
.A2(n_8680),
.B(n_8673),
.Y(n_10124)
);

NAND2xp5_ASAP7_75t_L g10125 ( 
.A(n_8390),
.B(n_8118),
.Y(n_10125)
);

OAI21x1_ASAP7_75t_L g10126 ( 
.A1(n_8426),
.A2(n_8637),
.B(n_8631),
.Y(n_10126)
);

INVx2_ASAP7_75t_L g10127 ( 
.A(n_8399),
.Y(n_10127)
);

INVx1_ASAP7_75t_L g10128 ( 
.A(n_8591),
.Y(n_10128)
);

OAI21x1_ASAP7_75t_L g10129 ( 
.A1(n_8426),
.A2(n_8637),
.B(n_8631),
.Y(n_10129)
);

HB1xp67_ASAP7_75t_L g10130 ( 
.A(n_8585),
.Y(n_10130)
);

NAND2x1p5_ASAP7_75t_L g10131 ( 
.A(n_7901),
.B(n_8103),
.Y(n_10131)
);

INVx3_ASAP7_75t_L g10132 ( 
.A(n_8899),
.Y(n_10132)
);

INVx1_ASAP7_75t_L g10133 ( 
.A(n_8591),
.Y(n_10133)
);

NAND2xp5_ASAP7_75t_L g10134 ( 
.A(n_8119),
.B(n_8900),
.Y(n_10134)
);

CKINVDCx6p67_ASAP7_75t_R g10135 ( 
.A(n_8608),
.Y(n_10135)
);

OAI21x1_ASAP7_75t_L g10136 ( 
.A1(n_8631),
.A2(n_8651),
.B(n_8637),
.Y(n_10136)
);

INVx6_ASAP7_75t_L g10137 ( 
.A(n_8300),
.Y(n_10137)
);

OAI21xp5_ASAP7_75t_L g10138 ( 
.A1(n_8395),
.A2(n_8013),
.B(n_8143),
.Y(n_10138)
);

OA21x2_ASAP7_75t_L g10139 ( 
.A1(n_8784),
.A2(n_8731),
.B(n_8680),
.Y(n_10139)
);

OA21x2_ASAP7_75t_L g10140 ( 
.A1(n_8293),
.A2(n_8163),
.B(n_8727),
.Y(n_10140)
);

O2A1O1Ixp33_ASAP7_75t_L g10141 ( 
.A1(n_8470),
.A2(n_8052),
.B(n_7741),
.C(n_8028),
.Y(n_10141)
);

INVx1_ASAP7_75t_L g10142 ( 
.A(n_8591),
.Y(n_10142)
);

INVx1_ASAP7_75t_SL g10143 ( 
.A(n_8862),
.Y(n_10143)
);

OAI21x1_ASAP7_75t_L g10144 ( 
.A1(n_8637),
.A2(n_8651),
.B(n_8205),
.Y(n_10144)
);

OAI21x1_ASAP7_75t_L g10145 ( 
.A1(n_8651),
.A2(n_8205),
.B(n_8204),
.Y(n_10145)
);

NOR2x1_ASAP7_75t_R g10146 ( 
.A(n_8608),
.B(n_8282),
.Y(n_10146)
);

OAI21x1_ASAP7_75t_L g10147 ( 
.A1(n_8651),
.A2(n_8205),
.B(n_8204),
.Y(n_10147)
);

CKINVDCx16_ASAP7_75t_R g10148 ( 
.A(n_8737),
.Y(n_10148)
);

AOI22xp33_ASAP7_75t_L g10149 ( 
.A1(n_7982),
.A2(n_8295),
.B1(n_7827),
.B2(n_8047),
.Y(n_10149)
);

INVx1_ASAP7_75t_L g10150 ( 
.A(n_8593),
.Y(n_10150)
);

AOI321xp33_ASAP7_75t_L g10151 ( 
.A1(n_8143),
.A2(n_8571),
.A3(n_7982),
.B1(n_8111),
.B2(n_8047),
.C(n_7697),
.Y(n_10151)
);

CKINVDCx5p33_ASAP7_75t_R g10152 ( 
.A(n_8078),
.Y(n_10152)
);

AOI22xp33_ASAP7_75t_L g10153 ( 
.A1(n_7827),
.A2(n_8194),
.B1(n_8028),
.B2(n_8052),
.Y(n_10153)
);

INVx3_ASAP7_75t_L g10154 ( 
.A(n_8899),
.Y(n_10154)
);

INVx3_ASAP7_75t_L g10155 ( 
.A(n_8899),
.Y(n_10155)
);

OR2x2_ASAP7_75t_L g10156 ( 
.A(n_7954),
.B(n_7957),
.Y(n_10156)
);

AOI21xp5_ASAP7_75t_L g10157 ( 
.A1(n_8577),
.A2(n_8541),
.B(n_8428),
.Y(n_10157)
);

NOR2xp33_ASAP7_75t_L g10158 ( 
.A(n_7823),
.B(n_7826),
.Y(n_10158)
);

INVx6_ASAP7_75t_L g10159 ( 
.A(n_8300),
.Y(n_10159)
);

NOR2xp67_ASAP7_75t_L g10160 ( 
.A(n_7901),
.B(n_8300),
.Y(n_10160)
);

BUFx2_ASAP7_75t_L g10161 ( 
.A(n_8689),
.Y(n_10161)
);

OA21x2_ASAP7_75t_L g10162 ( 
.A1(n_8293),
.A2(n_8163),
.B(n_8727),
.Y(n_10162)
);

OAI21xp5_ASAP7_75t_L g10163 ( 
.A1(n_8395),
.A2(n_8013),
.B(n_8085),
.Y(n_10163)
);

INVx1_ASAP7_75t_L g10164 ( 
.A(n_8593),
.Y(n_10164)
);

NAND2xp5_ASAP7_75t_L g10165 ( 
.A(n_8119),
.B(n_8900),
.Y(n_10165)
);

OAI21x1_ASAP7_75t_L g10166 ( 
.A1(n_8211),
.A2(n_8232),
.B(n_8226),
.Y(n_10166)
);

AO21x1_ASAP7_75t_L g10167 ( 
.A1(n_8446),
.A2(n_8462),
.B(n_8170),
.Y(n_10167)
);

OAI21xp5_ASAP7_75t_L g10168 ( 
.A1(n_8013),
.A2(n_8085),
.B(n_8259),
.Y(n_10168)
);

INVx3_ASAP7_75t_L g10169 ( 
.A(n_8899),
.Y(n_10169)
);

INVx1_ASAP7_75t_L g10170 ( 
.A(n_8593),
.Y(n_10170)
);

OAI21x1_ASAP7_75t_L g10171 ( 
.A1(n_8211),
.A2(n_8232),
.B(n_8226),
.Y(n_10171)
);

BUFx2_ASAP7_75t_L g10172 ( 
.A(n_8689),
.Y(n_10172)
);

BUFx2_ASAP7_75t_L g10173 ( 
.A(n_8689),
.Y(n_10173)
);

NAND2xp5_ASAP7_75t_L g10174 ( 
.A(n_8900),
.B(n_8838),
.Y(n_10174)
);

NOR2xp33_ASAP7_75t_SL g10175 ( 
.A(n_8061),
.B(n_7792),
.Y(n_10175)
);

OAI21x1_ASAP7_75t_L g10176 ( 
.A1(n_8232),
.A2(n_8237),
.B(n_8236),
.Y(n_10176)
);

INVx1_ASAP7_75t_L g10177 ( 
.A(n_8595),
.Y(n_10177)
);

OAI21x1_ASAP7_75t_SL g10178 ( 
.A1(n_8032),
.A2(n_8285),
.B(n_7705),
.Y(n_10178)
);

INVx2_ASAP7_75t_L g10179 ( 
.A(n_8644),
.Y(n_10179)
);

OA21x2_ASAP7_75t_L g10180 ( 
.A1(n_8727),
.A2(n_8732),
.B(n_8922),
.Y(n_10180)
);

BUFx6f_ASAP7_75t_L g10181 ( 
.A(n_8689),
.Y(n_10181)
);

INVx1_ASAP7_75t_L g10182 ( 
.A(n_8595),
.Y(n_10182)
);

OAI21x1_ASAP7_75t_L g10183 ( 
.A1(n_8236),
.A2(n_8238),
.B(n_8237),
.Y(n_10183)
);

OA21x2_ASAP7_75t_L g10184 ( 
.A1(n_8732),
.A2(n_8923),
.B(n_8922),
.Y(n_10184)
);

OAI21x1_ASAP7_75t_L g10185 ( 
.A1(n_8236),
.A2(n_8238),
.B(n_8237),
.Y(n_10185)
);

OAI21xp5_ASAP7_75t_SL g10186 ( 
.A1(n_7697),
.A2(n_8361),
.B(n_8391),
.Y(n_10186)
);

AND2x2_ASAP7_75t_L g10187 ( 
.A(n_8756),
.B(n_7894),
.Y(n_10187)
);

NOR2xp67_ASAP7_75t_SL g10188 ( 
.A(n_7717),
.B(n_8337),
.Y(n_10188)
);

NOR2x1_ASAP7_75t_SL g10189 ( 
.A(n_8165),
.B(n_8208),
.Y(n_10189)
);

BUFx2_ASAP7_75t_L g10190 ( 
.A(n_8689),
.Y(n_10190)
);

OAI21x1_ASAP7_75t_SL g10191 ( 
.A1(n_8285),
.A2(n_7705),
.B(n_8528),
.Y(n_10191)
);

INVx1_ASAP7_75t_L g10192 ( 
.A(n_8595),
.Y(n_10192)
);

NOR2x1_ASAP7_75t_SL g10193 ( 
.A(n_8208),
.B(n_8943),
.Y(n_10193)
);

OAI21x1_ASAP7_75t_SL g10194 ( 
.A1(n_9003),
.A2(n_7705),
.B(n_8425),
.Y(n_10194)
);

INVx2_ASAP7_75t_L g10195 ( 
.A(n_9435),
.Y(n_10195)
);

INVx1_ASAP7_75t_L g10196 ( 
.A(n_10128),
.Y(n_10196)
);

INVx1_ASAP7_75t_L g10197 ( 
.A(n_10128),
.Y(n_10197)
);

INVx2_ASAP7_75t_L g10198 ( 
.A(n_9435),
.Y(n_10198)
);

AND2x4_ASAP7_75t_L g10199 ( 
.A(n_9589),
.B(n_7930),
.Y(n_10199)
);

NAND2xp5_ASAP7_75t_L g10200 ( 
.A(n_10096),
.B(n_8332),
.Y(n_10200)
);

NOR2xp67_ASAP7_75t_L g10201 ( 
.A(n_9467),
.B(n_7930),
.Y(n_10201)
);

OA21x2_ASAP7_75t_L g10202 ( 
.A1(n_9486),
.A2(n_8238),
.B(n_8237),
.Y(n_10202)
);

INVx2_ASAP7_75t_SL g10203 ( 
.A(n_9441),
.Y(n_10203)
);

OAI21x1_ASAP7_75t_L g10204 ( 
.A1(n_9135),
.A2(n_8584),
.B(n_8583),
.Y(n_10204)
);

OAI21x1_ASAP7_75t_L g10205 ( 
.A1(n_9135),
.A2(n_8584),
.B(n_8583),
.Y(n_10205)
);

OA21x2_ASAP7_75t_L g10206 ( 
.A1(n_9486),
.A2(n_8249),
.B(n_8238),
.Y(n_10206)
);

INVx1_ASAP7_75t_L g10207 ( 
.A(n_10128),
.Y(n_10207)
);

NAND2xp5_ASAP7_75t_L g10208 ( 
.A(n_10096),
.B(n_8332),
.Y(n_10208)
);

AOI21xp5_ASAP7_75t_L g10209 ( 
.A1(n_9473),
.A2(n_8470),
.B(n_8519),
.Y(n_10209)
);

OAI21x1_ASAP7_75t_L g10210 ( 
.A1(n_9135),
.A2(n_8590),
.B(n_8588),
.Y(n_10210)
);

AO31x2_ASAP7_75t_L g10211 ( 
.A1(n_9003),
.A2(n_8255),
.A3(n_8570),
.B(n_8669),
.Y(n_10211)
);

INVx2_ASAP7_75t_SL g10212 ( 
.A(n_9441),
.Y(n_10212)
);

INVx1_ASAP7_75t_L g10213 ( 
.A(n_10128),
.Y(n_10213)
);

AO21x1_ASAP7_75t_L g10214 ( 
.A1(n_9137),
.A2(n_8462),
.B(n_8446),
.Y(n_10214)
);

NAND2xp5_ASAP7_75t_L g10215 ( 
.A(n_10096),
.B(n_7989),
.Y(n_10215)
);

INVx1_ASAP7_75t_SL g10216 ( 
.A(n_9087),
.Y(n_10216)
);

AO31x2_ASAP7_75t_L g10217 ( 
.A1(n_9003),
.A2(n_8255),
.A3(n_8570),
.B(n_8573),
.Y(n_10217)
);

INVx2_ASAP7_75t_SL g10218 ( 
.A(n_9441),
.Y(n_10218)
);

INVx6_ASAP7_75t_L g10219 ( 
.A(n_9073),
.Y(n_10219)
);

OAI21x1_ASAP7_75t_L g10220 ( 
.A1(n_9135),
.A2(n_8590),
.B(n_8588),
.Y(n_10220)
);

INVx2_ASAP7_75t_L g10221 ( 
.A(n_9435),
.Y(n_10221)
);

INVx1_ASAP7_75t_L g10222 ( 
.A(n_10133),
.Y(n_10222)
);

AND2x4_ASAP7_75t_L g10223 ( 
.A(n_9589),
.B(n_7930),
.Y(n_10223)
);

OAI21x1_ASAP7_75t_L g10224 ( 
.A1(n_9135),
.A2(n_8603),
.B(n_8596),
.Y(n_10224)
);

OA21x2_ASAP7_75t_L g10225 ( 
.A1(n_9486),
.A2(n_8268),
.B(n_8249),
.Y(n_10225)
);

AO31x2_ASAP7_75t_L g10226 ( 
.A1(n_9003),
.A2(n_9319),
.A3(n_10167),
.B(n_9012),
.Y(n_10226)
);

AO31x2_ASAP7_75t_L g10227 ( 
.A1(n_9003),
.A2(n_8255),
.A3(n_8573),
.B(n_8313),
.Y(n_10227)
);

INVx1_ASAP7_75t_L g10228 ( 
.A(n_10133),
.Y(n_10228)
);

AOI22xp33_ASAP7_75t_L g10229 ( 
.A1(n_8975),
.A2(n_7827),
.B1(n_8194),
.B2(n_8071),
.Y(n_10229)
);

OA21x2_ASAP7_75t_L g10230 ( 
.A1(n_9539),
.A2(n_8268),
.B(n_8249),
.Y(n_10230)
);

BUFx2_ASAP7_75t_L g10231 ( 
.A(n_9975),
.Y(n_10231)
);

AND2x4_ASAP7_75t_L g10232 ( 
.A(n_9589),
.B(n_7930),
.Y(n_10232)
);

CKINVDCx6p67_ASAP7_75t_R g10233 ( 
.A(n_9143),
.Y(n_10233)
);

BUFx3_ASAP7_75t_L g10234 ( 
.A(n_9073),
.Y(n_10234)
);

INVx1_ASAP7_75t_L g10235 ( 
.A(n_10133),
.Y(n_10235)
);

AOI22x1_ASAP7_75t_L g10236 ( 
.A1(n_9630),
.A2(n_8071),
.B1(n_8305),
.B2(n_8282),
.Y(n_10236)
);

NOR2xp33_ASAP7_75t_SL g10237 ( 
.A(n_9208),
.B(n_7808),
.Y(n_10237)
);

AO31x2_ASAP7_75t_L g10238 ( 
.A1(n_9319),
.A2(n_8573),
.A3(n_8313),
.B(n_8673),
.Y(n_10238)
);

BUFx3_ASAP7_75t_L g10239 ( 
.A(n_9073),
.Y(n_10239)
);

AOI22xp33_ASAP7_75t_L g10240 ( 
.A1(n_8975),
.A2(n_7827),
.B1(n_8194),
.B2(n_8071),
.Y(n_10240)
);

INVx1_ASAP7_75t_L g10241 ( 
.A(n_10133),
.Y(n_10241)
);

NOR2xp67_ASAP7_75t_L g10242 ( 
.A(n_9467),
.B(n_8007),
.Y(n_10242)
);

AOI21x1_ASAP7_75t_L g10243 ( 
.A1(n_9088),
.A2(n_8053),
.B(n_8045),
.Y(n_10243)
);

AND2x2_ASAP7_75t_L g10244 ( 
.A(n_9876),
.B(n_8007),
.Y(n_10244)
);

NAND2x1_ASAP7_75t_L g10245 ( 
.A(n_9952),
.B(n_9976),
.Y(n_10245)
);

INVx4_ASAP7_75t_SL g10246 ( 
.A(n_9388),
.Y(n_10246)
);

INVx5_ASAP7_75t_L g10247 ( 
.A(n_10148),
.Y(n_10247)
);

OA21x2_ASAP7_75t_L g10248 ( 
.A1(n_9539),
.A2(n_8268),
.B(n_8249),
.Y(n_10248)
);

OAI21x1_ASAP7_75t_L g10249 ( 
.A1(n_9136),
.A2(n_8603),
.B(n_8596),
.Y(n_10249)
);

INVx1_ASAP7_75t_L g10250 ( 
.A(n_10142),
.Y(n_10250)
);

INVx1_ASAP7_75t_SL g10251 ( 
.A(n_9087),
.Y(n_10251)
);

INVxp67_ASAP7_75t_SL g10252 ( 
.A(n_9012),
.Y(n_10252)
);

NAND2xp5_ASAP7_75t_L g10253 ( 
.A(n_9932),
.B(n_7989),
.Y(n_10253)
);

AOI21x1_ASAP7_75t_L g10254 ( 
.A1(n_9088),
.A2(n_8053),
.B(n_8045),
.Y(n_10254)
);

AO31x2_ASAP7_75t_L g10255 ( 
.A1(n_9319),
.A2(n_8633),
.A3(n_8766),
.B(n_8761),
.Y(n_10255)
);

OAI21x1_ASAP7_75t_L g10256 ( 
.A1(n_9136),
.A2(n_8600),
.B(n_8621),
.Y(n_10256)
);

INVx1_ASAP7_75t_L g10257 ( 
.A(n_10142),
.Y(n_10257)
);

INVx1_ASAP7_75t_L g10258 ( 
.A(n_10142),
.Y(n_10258)
);

OAI21x1_ASAP7_75t_SL g10259 ( 
.A1(n_9473),
.A2(n_8425),
.B(n_8361),
.Y(n_10259)
);

INVx2_ASAP7_75t_L g10260 ( 
.A(n_9323),
.Y(n_10260)
);

INVx1_ASAP7_75t_L g10261 ( 
.A(n_10142),
.Y(n_10261)
);

INVx1_ASAP7_75t_L g10262 ( 
.A(n_10150),
.Y(n_10262)
);

OR3x4_ASAP7_75t_SL g10263 ( 
.A(n_9143),
.B(n_9014),
.C(n_10041),
.Y(n_10263)
);

INVx2_ASAP7_75t_L g10264 ( 
.A(n_9323),
.Y(n_10264)
);

NAND2xp5_ASAP7_75t_L g10265 ( 
.A(n_9932),
.B(n_9987),
.Y(n_10265)
);

AOI21x1_ASAP7_75t_L g10266 ( 
.A1(n_9088),
.A2(n_8053),
.B(n_8045),
.Y(n_10266)
);

OA21x2_ASAP7_75t_L g10267 ( 
.A1(n_9539),
.A2(n_8272),
.B(n_8268),
.Y(n_10267)
);

NAND2x1p5_ASAP7_75t_L g10268 ( 
.A(n_9110),
.B(n_8208),
.Y(n_10268)
);

AOI21xp33_ASAP7_75t_L g10269 ( 
.A1(n_9206),
.A2(n_8319),
.B(n_8629),
.Y(n_10269)
);

INVx1_ASAP7_75t_L g10270 ( 
.A(n_10150),
.Y(n_10270)
);

BUFx8_ASAP7_75t_L g10271 ( 
.A(n_9148),
.Y(n_10271)
);

CKINVDCx5p33_ASAP7_75t_R g10272 ( 
.A(n_9422),
.Y(n_10272)
);

INVx2_ASAP7_75t_L g10273 ( 
.A(n_9323),
.Y(n_10273)
);

INVx1_ASAP7_75t_L g10274 ( 
.A(n_10150),
.Y(n_10274)
);

OAI21x1_ASAP7_75t_SL g10275 ( 
.A1(n_9473),
.A2(n_8391),
.B(n_8427),
.Y(n_10275)
);

OAI21x1_ASAP7_75t_L g10276 ( 
.A1(n_9136),
.A2(n_8600),
.B(n_8621),
.Y(n_10276)
);

NAND2xp5_ASAP7_75t_L g10277 ( 
.A(n_9932),
.B(n_7990),
.Y(n_10277)
);

HB1xp67_ASAP7_75t_L g10278 ( 
.A(n_9205),
.Y(n_10278)
);

OAI21x1_ASAP7_75t_L g10279 ( 
.A1(n_9136),
.A2(n_8600),
.B(n_8624),
.Y(n_10279)
);

OAI21x1_ASAP7_75t_L g10280 ( 
.A1(n_9136),
.A2(n_8624),
.B(n_8412),
.Y(n_10280)
);

OAI21x1_ASAP7_75t_L g10281 ( 
.A1(n_8991),
.A2(n_8412),
.B(n_8417),
.Y(n_10281)
);

INVx2_ASAP7_75t_L g10282 ( 
.A(n_9323),
.Y(n_10282)
);

BUFx2_ASAP7_75t_L g10283 ( 
.A(n_9975),
.Y(n_10283)
);

NAND2xp5_ASAP7_75t_L g10284 ( 
.A(n_9987),
.B(n_7990),
.Y(n_10284)
);

NOR2xp67_ASAP7_75t_SL g10285 ( 
.A(n_9208),
.B(n_8608),
.Y(n_10285)
);

BUFx2_ASAP7_75t_L g10286 ( 
.A(n_9975),
.Y(n_10286)
);

OAI21x1_ASAP7_75t_L g10287 ( 
.A1(n_8991),
.A2(n_8417),
.B(n_8489),
.Y(n_10287)
);

OA21x2_ASAP7_75t_L g10288 ( 
.A1(n_9656),
.A2(n_8275),
.B(n_8272),
.Y(n_10288)
);

OAI21xp33_ASAP7_75t_L g10289 ( 
.A1(n_9591),
.A2(n_8571),
.B(n_8330),
.Y(n_10289)
);

OAI21x1_ASAP7_75t_L g10290 ( 
.A1(n_8991),
.A2(n_8489),
.B(n_8664),
.Y(n_10290)
);

OAI21xp5_ASAP7_75t_L g10291 ( 
.A1(n_9630),
.A2(n_8493),
.B(n_8330),
.Y(n_10291)
);

NAND2xp5_ASAP7_75t_L g10292 ( 
.A(n_9987),
.B(n_7893),
.Y(n_10292)
);

INVx2_ASAP7_75t_L g10293 ( 
.A(n_9323),
.Y(n_10293)
);

INVx2_ASAP7_75t_L g10294 ( 
.A(n_9323),
.Y(n_10294)
);

BUFx2_ASAP7_75t_L g10295 ( 
.A(n_9975),
.Y(n_10295)
);

OA21x2_ASAP7_75t_L g10296 ( 
.A1(n_9656),
.A2(n_8275),
.B(n_8272),
.Y(n_10296)
);

OAI21x1_ASAP7_75t_L g10297 ( 
.A1(n_8991),
.A2(n_8489),
.B(n_8664),
.Y(n_10297)
);

AO21x2_ASAP7_75t_L g10298 ( 
.A1(n_10163),
.A2(n_8428),
.B(n_8247),
.Y(n_10298)
);

BUFx3_ASAP7_75t_L g10299 ( 
.A(n_9073),
.Y(n_10299)
);

OAI21x1_ASAP7_75t_L g10300 ( 
.A1(n_8991),
.A2(n_8489),
.B(n_8664),
.Y(n_10300)
);

INVx1_ASAP7_75t_L g10301 ( 
.A(n_10150),
.Y(n_10301)
);

OA21x2_ASAP7_75t_L g10302 ( 
.A1(n_9656),
.A2(n_8275),
.B(n_8272),
.Y(n_10302)
);

OA21x2_ASAP7_75t_L g10303 ( 
.A1(n_9656),
.A2(n_8275),
.B(n_8922),
.Y(n_10303)
);

OR2x2_ASAP7_75t_L g10304 ( 
.A(n_10156),
.B(n_8384),
.Y(n_10304)
);

INVx1_ASAP7_75t_L g10305 ( 
.A(n_10164),
.Y(n_10305)
);

AO21x2_ASAP7_75t_L g10306 ( 
.A1(n_10163),
.A2(n_8247),
.B(n_8246),
.Y(n_10306)
);

OR2x2_ASAP7_75t_L g10307 ( 
.A(n_10156),
.B(n_8384),
.Y(n_10307)
);

AO31x2_ASAP7_75t_L g10308 ( 
.A1(n_9319),
.A2(n_10167),
.A3(n_9012),
.B(n_8980),
.Y(n_10308)
);

NAND2xp5_ASAP7_75t_L g10309 ( 
.A(n_10082),
.B(n_8564),
.Y(n_10309)
);

BUFx2_ASAP7_75t_L g10310 ( 
.A(n_9975),
.Y(n_10310)
);

AOI21x1_ASAP7_75t_L g10311 ( 
.A1(n_9088),
.A2(n_8367),
.B(n_8732),
.Y(n_10311)
);

INVx1_ASAP7_75t_L g10312 ( 
.A(n_10164),
.Y(n_10312)
);

NAND2xp5_ASAP7_75t_L g10313 ( 
.A(n_10082),
.B(n_8564),
.Y(n_10313)
);

AOI21x1_ASAP7_75t_L g10314 ( 
.A1(n_10188),
.A2(n_8367),
.B(n_8941),
.Y(n_10314)
);

OA21x2_ASAP7_75t_L g10315 ( 
.A1(n_9661),
.A2(n_9673),
.B(n_9664),
.Y(n_10315)
);

OAI21x1_ASAP7_75t_L g10316 ( 
.A1(n_9188),
.A2(n_8672),
.B(n_8664),
.Y(n_10316)
);

INVx1_ASAP7_75t_L g10317 ( 
.A(n_10164),
.Y(n_10317)
);

INVx3_ASAP7_75t_L g10318 ( 
.A(n_9589),
.Y(n_10318)
);

NAND2x1p5_ASAP7_75t_L g10319 ( 
.A(n_9110),
.B(n_8208),
.Y(n_10319)
);

OAI21x1_ASAP7_75t_L g10320 ( 
.A1(n_9188),
.A2(n_8678),
.B(n_8672),
.Y(n_10320)
);

INVx1_ASAP7_75t_L g10321 ( 
.A(n_10164),
.Y(n_10321)
);

OAI21x1_ASAP7_75t_L g10322 ( 
.A1(n_9188),
.A2(n_8678),
.B(n_8672),
.Y(n_10322)
);

INVx3_ASAP7_75t_L g10323 ( 
.A(n_9589),
.Y(n_10323)
);

NAND2xp5_ASAP7_75t_L g10324 ( 
.A(n_10082),
.B(n_7829),
.Y(n_10324)
);

AOI22xp5_ASAP7_75t_L g10325 ( 
.A1(n_9591),
.A2(n_7943),
.B1(n_8129),
.B2(n_7953),
.Y(n_10325)
);

OAI21x1_ASAP7_75t_L g10326 ( 
.A1(n_9188),
.A2(n_8678),
.B(n_8672),
.Y(n_10326)
);

BUFx2_ASAP7_75t_L g10327 ( 
.A(n_9975),
.Y(n_10327)
);

AO31x2_ASAP7_75t_L g10328 ( 
.A1(n_9319),
.A2(n_10167),
.A3(n_9012),
.B(n_8980),
.Y(n_10328)
);

A2O1A1Ixp33_ASAP7_75t_L g10329 ( 
.A1(n_10089),
.A2(n_8561),
.B(n_8576),
.C(n_8452),
.Y(n_10329)
);

INVx1_ASAP7_75t_L g10330 ( 
.A(n_10170),
.Y(n_10330)
);

NOR2xp33_ASAP7_75t_R g10331 ( 
.A(n_9014),
.B(n_8481),
.Y(n_10331)
);

AO21x2_ASAP7_75t_L g10332 ( 
.A1(n_10163),
.A2(n_8246),
.B(n_8516),
.Y(n_10332)
);

INVx3_ASAP7_75t_L g10333 ( 
.A(n_9589),
.Y(n_10333)
);

OAI21x1_ASAP7_75t_L g10334 ( 
.A1(n_9188),
.A2(n_8690),
.B(n_8678),
.Y(n_10334)
);

OR2x2_ASAP7_75t_L g10335 ( 
.A(n_10156),
.B(n_8384),
.Y(n_10335)
);

OAI21x1_ASAP7_75t_L g10336 ( 
.A1(n_8978),
.A2(n_8696),
.B(n_8690),
.Y(n_10336)
);

INVx3_ASAP7_75t_L g10337 ( 
.A(n_9596),
.Y(n_10337)
);

NAND2xp5_ASAP7_75t_L g10338 ( 
.A(n_9022),
.B(n_7829),
.Y(n_10338)
);

OA21x2_ASAP7_75t_L g10339 ( 
.A1(n_9661),
.A2(n_8923),
.B(n_8922),
.Y(n_10339)
);

OR2x2_ASAP7_75t_L g10340 ( 
.A(n_10156),
.B(n_9889),
.Y(n_10340)
);

OAI21x1_ASAP7_75t_L g10341 ( 
.A1(n_8978),
.A2(n_8696),
.B(n_8690),
.Y(n_10341)
);

NAND2xp5_ASAP7_75t_L g10342 ( 
.A(n_9022),
.B(n_7922),
.Y(n_10342)
);

OAI21x1_ASAP7_75t_L g10343 ( 
.A1(n_8978),
.A2(n_9522),
.B(n_9609),
.Y(n_10343)
);

AO21x2_ASAP7_75t_L g10344 ( 
.A1(n_9639),
.A2(n_8516),
.B(n_8319),
.Y(n_10344)
);

OR2x6_ASAP7_75t_L g10345 ( 
.A(n_10114),
.B(n_9441),
.Y(n_10345)
);

NOR3xp33_ASAP7_75t_SL g10346 ( 
.A(n_9630),
.B(n_8466),
.C(n_8481),
.Y(n_10346)
);

INVx2_ASAP7_75t_L g10347 ( 
.A(n_9435),
.Y(n_10347)
);

OR2x2_ASAP7_75t_L g10348 ( 
.A(n_10156),
.B(n_8384),
.Y(n_10348)
);

NAND2xp5_ASAP7_75t_L g10349 ( 
.A(n_9022),
.B(n_10113),
.Y(n_10349)
);

INVx2_ASAP7_75t_L g10350 ( 
.A(n_9435),
.Y(n_10350)
);

OAI21x1_ASAP7_75t_L g10351 ( 
.A1(n_8978),
.A2(n_8696),
.B(n_8690),
.Y(n_10351)
);

INVx1_ASAP7_75t_L g10352 ( 
.A(n_10170),
.Y(n_10352)
);

INVx2_ASAP7_75t_L g10353 ( 
.A(n_9435),
.Y(n_10353)
);

INVx1_ASAP7_75t_L g10354 ( 
.A(n_10170),
.Y(n_10354)
);

HB1xp67_ASAP7_75t_L g10355 ( 
.A(n_9205),
.Y(n_10355)
);

INVx1_ASAP7_75t_L g10356 ( 
.A(n_10170),
.Y(n_10356)
);

INVx1_ASAP7_75t_L g10357 ( 
.A(n_10177),
.Y(n_10357)
);

NAND2x1p5_ASAP7_75t_L g10358 ( 
.A(n_9110),
.B(n_9370),
.Y(n_10358)
);

INVx2_ASAP7_75t_L g10359 ( 
.A(n_9435),
.Y(n_10359)
);

NAND2xp5_ASAP7_75t_L g10360 ( 
.A(n_10113),
.B(n_10125),
.Y(n_10360)
);

AO21x1_ASAP7_75t_L g10361 ( 
.A1(n_9137),
.A2(n_8479),
.B(n_8482),
.Y(n_10361)
);

AO31x2_ASAP7_75t_L g10362 ( 
.A1(n_10167),
.A2(n_8633),
.A3(n_8766),
.B(n_8761),
.Y(n_10362)
);

AO21x1_ASAP7_75t_L g10363 ( 
.A1(n_9137),
.A2(n_8479),
.B(n_8482),
.Y(n_10363)
);

HB1xp67_ASAP7_75t_L g10364 ( 
.A(n_9205),
.Y(n_10364)
);

AND2x4_ASAP7_75t_L g10365 ( 
.A(n_9596),
.B(n_9600),
.Y(n_10365)
);

AOI22x1_ASAP7_75t_L g10366 ( 
.A1(n_9560),
.A2(n_8071),
.B1(n_8305),
.B2(n_8180),
.Y(n_10366)
);

INVxp67_ASAP7_75t_SL g10367 ( 
.A(n_9012),
.Y(n_10367)
);

NAND2xp5_ASAP7_75t_L g10368 ( 
.A(n_10113),
.B(n_7922),
.Y(n_10368)
);

CKINVDCx11_ASAP7_75t_R g10369 ( 
.A(n_9014),
.Y(n_10369)
);

AND2x4_ASAP7_75t_L g10370 ( 
.A(n_9596),
.B(n_8007),
.Y(n_10370)
);

INVx1_ASAP7_75t_L g10371 ( 
.A(n_10177),
.Y(n_10371)
);

INVx2_ASAP7_75t_L g10372 ( 
.A(n_9435),
.Y(n_10372)
);

INVx3_ASAP7_75t_L g10373 ( 
.A(n_9596),
.Y(n_10373)
);

INVx2_ASAP7_75t_L g10374 ( 
.A(n_9323),
.Y(n_10374)
);

INVx2_ASAP7_75t_L g10375 ( 
.A(n_9323),
.Y(n_10375)
);

OAI21x1_ASAP7_75t_L g10376 ( 
.A1(n_8978),
.A2(n_9522),
.B(n_9609),
.Y(n_10376)
);

CKINVDCx20_ASAP7_75t_R g10377 ( 
.A(n_9149),
.Y(n_10377)
);

BUFx6f_ASAP7_75t_L g10378 ( 
.A(n_9110),
.Y(n_10378)
);

CKINVDCx11_ASAP7_75t_R g10379 ( 
.A(n_9143),
.Y(n_10379)
);

INVx2_ASAP7_75t_L g10380 ( 
.A(n_9323),
.Y(n_10380)
);

AOI21x1_ASAP7_75t_L g10381 ( 
.A1(n_10188),
.A2(n_8367),
.B(n_8941),
.Y(n_10381)
);

INVxp67_ASAP7_75t_L g10382 ( 
.A(n_9868),
.Y(n_10382)
);

AO21x2_ASAP7_75t_L g10383 ( 
.A1(n_9639),
.A2(n_8116),
.B(n_8574),
.Y(n_10383)
);

OAI21x1_ASAP7_75t_L g10384 ( 
.A1(n_9522),
.A2(n_8707),
.B(n_8696),
.Y(n_10384)
);

INVx1_ASAP7_75t_L g10385 ( 
.A(n_10177),
.Y(n_10385)
);

NAND2xp5_ASAP7_75t_L g10386 ( 
.A(n_10125),
.B(n_7826),
.Y(n_10386)
);

INVx3_ASAP7_75t_L g10387 ( 
.A(n_9596),
.Y(n_10387)
);

AO21x2_ASAP7_75t_L g10388 ( 
.A1(n_9639),
.A2(n_8116),
.B(n_8574),
.Y(n_10388)
);

INVx2_ASAP7_75t_L g10389 ( 
.A(n_9435),
.Y(n_10389)
);

OAI21x1_ASAP7_75t_L g10390 ( 
.A1(n_9522),
.A2(n_8719),
.B(n_8707),
.Y(n_10390)
);

OAI21x1_ASAP7_75t_L g10391 ( 
.A1(n_9522),
.A2(n_8719),
.B(n_8707),
.Y(n_10391)
);

AO21x1_ASAP7_75t_L g10392 ( 
.A1(n_9868),
.A2(n_9206),
.B(n_9898),
.Y(n_10392)
);

BUFx3_ASAP7_75t_L g10393 ( 
.A(n_9073),
.Y(n_10393)
);

INVx1_ASAP7_75t_L g10394 ( 
.A(n_10177),
.Y(n_10394)
);

INVx1_ASAP7_75t_L g10395 ( 
.A(n_10182),
.Y(n_10395)
);

A2O1A1Ixp33_ASAP7_75t_L g10396 ( 
.A1(n_10089),
.A2(n_8561),
.B(n_8576),
.C(n_8452),
.Y(n_10396)
);

OAI21x1_ASAP7_75t_L g10397 ( 
.A1(n_9609),
.A2(n_8719),
.B(n_8707),
.Y(n_10397)
);

OAI21x1_ASAP7_75t_L g10398 ( 
.A1(n_9609),
.A2(n_8721),
.B(n_8719),
.Y(n_10398)
);

INVx2_ASAP7_75t_L g10399 ( 
.A(n_9336),
.Y(n_10399)
);

AOI21xp5_ASAP7_75t_L g10400 ( 
.A1(n_10044),
.A2(n_8526),
.B(n_8519),
.Y(n_10400)
);

INVx1_ASAP7_75t_L g10401 ( 
.A(n_10182),
.Y(n_10401)
);

NAND3xp33_ASAP7_75t_L g10402 ( 
.A(n_9560),
.B(n_8153),
.C(n_8746),
.Y(n_10402)
);

OA21x2_ASAP7_75t_L g10403 ( 
.A1(n_9661),
.A2(n_8938),
.B(n_8923),
.Y(n_10403)
);

AO31x2_ASAP7_75t_L g10404 ( 
.A1(n_10167),
.A2(n_8594),
.A3(n_8347),
.B(n_8871),
.Y(n_10404)
);

OAI21x1_ASAP7_75t_L g10405 ( 
.A1(n_9203),
.A2(n_8721),
.B(n_8923),
.Y(n_10405)
);

INVx1_ASAP7_75t_L g10406 ( 
.A(n_10182),
.Y(n_10406)
);

OAI21x1_ASAP7_75t_L g10407 ( 
.A1(n_9203),
.A2(n_8721),
.B(n_8938),
.Y(n_10407)
);

AND2x2_ASAP7_75t_L g10408 ( 
.A(n_9876),
.B(n_8007),
.Y(n_10408)
);

OAI21xp5_ASAP7_75t_L g10409 ( 
.A1(n_9560),
.A2(n_8493),
.B(n_8129),
.Y(n_10409)
);

INVx1_ASAP7_75t_SL g10410 ( 
.A(n_9087),
.Y(n_10410)
);

OAI21x1_ASAP7_75t_L g10411 ( 
.A1(n_9203),
.A2(n_8721),
.B(n_8938),
.Y(n_10411)
);

OAI21x1_ASAP7_75t_L g10412 ( 
.A1(n_9203),
.A2(n_8945),
.B(n_8938),
.Y(n_10412)
);

NOR2xp33_ASAP7_75t_L g10413 ( 
.A(n_8975),
.B(n_7836),
.Y(n_10413)
);

INVx1_ASAP7_75t_L g10414 ( 
.A(n_10182),
.Y(n_10414)
);

INVx1_ASAP7_75t_L g10415 ( 
.A(n_10192),
.Y(n_10415)
);

NAND2xp5_ASAP7_75t_L g10416 ( 
.A(n_10125),
.B(n_7818),
.Y(n_10416)
);

AOI21x1_ASAP7_75t_L g10417 ( 
.A1(n_10188),
.A2(n_8941),
.B(n_8670),
.Y(n_10417)
);

INVx1_ASAP7_75t_L g10418 ( 
.A(n_10192),
.Y(n_10418)
);

AOI21x1_ASAP7_75t_L g10419 ( 
.A1(n_10188),
.A2(n_8670),
.B(n_8665),
.Y(n_10419)
);

NOR2x1_ASAP7_75t_SL g10420 ( 
.A(n_9272),
.B(n_8044),
.Y(n_10420)
);

OAI21x1_ASAP7_75t_L g10421 ( 
.A1(n_9203),
.A2(n_8947),
.B(n_8945),
.Y(n_10421)
);

INVx1_ASAP7_75t_SL g10422 ( 
.A(n_9134),
.Y(n_10422)
);

BUFx10_ASAP7_75t_L g10423 ( 
.A(n_9056),
.Y(n_10423)
);

AO21x2_ASAP7_75t_L g10424 ( 
.A1(n_10157),
.A2(n_8574),
.B(n_8223),
.Y(n_10424)
);

OAI21x1_ASAP7_75t_L g10425 ( 
.A1(n_9213),
.A2(n_8947),
.B(n_8945),
.Y(n_10425)
);

OAI21x1_ASAP7_75t_L g10426 ( 
.A1(n_9213),
.A2(n_8947),
.B(n_8945),
.Y(n_10426)
);

AND2x2_ASAP7_75t_L g10427 ( 
.A(n_9876),
.B(n_8019),
.Y(n_10427)
);

OAI21x1_ASAP7_75t_L g10428 ( 
.A1(n_9213),
.A2(n_8950),
.B(n_8947),
.Y(n_10428)
);

INVx1_ASAP7_75t_L g10429 ( 
.A(n_10192),
.Y(n_10429)
);

NAND2xp5_ASAP7_75t_L g10430 ( 
.A(n_9906),
.B(n_7818),
.Y(n_10430)
);

BUFx2_ASAP7_75t_L g10431 ( 
.A(n_9975),
.Y(n_10431)
);

OA21x2_ASAP7_75t_L g10432 ( 
.A1(n_9661),
.A2(n_8954),
.B(n_8950),
.Y(n_10432)
);

OAI21x1_ASAP7_75t_L g10433 ( 
.A1(n_9213),
.A2(n_8954),
.B(n_8950),
.Y(n_10433)
);

CKINVDCx5p33_ASAP7_75t_R g10434 ( 
.A(n_9422),
.Y(n_10434)
);

BUFx8_ASAP7_75t_L g10435 ( 
.A(n_9148),
.Y(n_10435)
);

INVx1_ASAP7_75t_L g10436 ( 
.A(n_10192),
.Y(n_10436)
);

AND2x2_ASAP7_75t_L g10437 ( 
.A(n_9876),
.B(n_8019),
.Y(n_10437)
);

AO21x2_ASAP7_75t_L g10438 ( 
.A1(n_10157),
.A2(n_8223),
.B(n_8172),
.Y(n_10438)
);

INVx1_ASAP7_75t_L g10439 ( 
.A(n_9801),
.Y(n_10439)
);

OA21x2_ASAP7_75t_L g10440 ( 
.A1(n_9664),
.A2(n_8954),
.B(n_8950),
.Y(n_10440)
);

HB1xp67_ASAP7_75t_L g10441 ( 
.A(n_9205),
.Y(n_10441)
);

INVx3_ASAP7_75t_L g10442 ( 
.A(n_9596),
.Y(n_10442)
);

AND2x4_ASAP7_75t_L g10443 ( 
.A(n_9600),
.B(n_8027),
.Y(n_10443)
);

OR2x2_ASAP7_75t_L g10444 ( 
.A(n_9889),
.B(n_8384),
.Y(n_10444)
);

CKINVDCx20_ASAP7_75t_R g10445 ( 
.A(n_9149),
.Y(n_10445)
);

BUFx2_ASAP7_75t_L g10446 ( 
.A(n_9975),
.Y(n_10446)
);

CKINVDCx5p33_ASAP7_75t_R g10447 ( 
.A(n_9422),
.Y(n_10447)
);

NOR2x1_ASAP7_75t_L g10448 ( 
.A(n_9868),
.B(n_8435),
.Y(n_10448)
);

INVx2_ASAP7_75t_L g10449 ( 
.A(n_9336),
.Y(n_10449)
);

NAND2xp5_ASAP7_75t_L g10450 ( 
.A(n_9906),
.B(n_8087),
.Y(n_10450)
);

AO21x2_ASAP7_75t_L g10451 ( 
.A1(n_10157),
.A2(n_8223),
.B(n_8172),
.Y(n_10451)
);

HB1xp67_ASAP7_75t_L g10452 ( 
.A(n_9205),
.Y(n_10452)
);

NAND2xp5_ASAP7_75t_SL g10453 ( 
.A(n_9898),
.B(n_8746),
.Y(n_10453)
);

CKINVDCx11_ASAP7_75t_R g10454 ( 
.A(n_9739),
.Y(n_10454)
);

INVx1_ASAP7_75t_L g10455 ( 
.A(n_9801),
.Y(n_10455)
);

INVx1_ASAP7_75t_L g10456 ( 
.A(n_9801),
.Y(n_10456)
);

AO31x2_ASAP7_75t_L g10457 ( 
.A1(n_8980),
.A2(n_8594),
.A3(n_8347),
.B(n_8871),
.Y(n_10457)
);

BUFx6f_ASAP7_75t_L g10458 ( 
.A(n_9110),
.Y(n_10458)
);

OAI21x1_ASAP7_75t_L g10459 ( 
.A1(n_9213),
.A2(n_9551),
.B(n_10114),
.Y(n_10459)
);

INVx6_ASAP7_75t_L g10460 ( 
.A(n_9073),
.Y(n_10460)
);

OR2x6_ASAP7_75t_L g10461 ( 
.A(n_10114),
.B(n_8876),
.Y(n_10461)
);

OAI21x1_ASAP7_75t_L g10462 ( 
.A1(n_9551),
.A2(n_8956),
.B(n_8954),
.Y(n_10462)
);

OAI21xp5_ASAP7_75t_L g10463 ( 
.A1(n_9897),
.A2(n_10089),
.B(n_9591),
.Y(n_10463)
);

AO21x2_ASAP7_75t_L g10464 ( 
.A1(n_9678),
.A2(n_8223),
.B(n_8172),
.Y(n_10464)
);

INVx3_ASAP7_75t_SL g10465 ( 
.A(n_9056),
.Y(n_10465)
);

AO21x2_ASAP7_75t_L g10466 ( 
.A1(n_9678),
.A2(n_8223),
.B(n_8172),
.Y(n_10466)
);

OAI21xp5_ASAP7_75t_L g10467 ( 
.A1(n_9897),
.A2(n_8493),
.B(n_8418),
.Y(n_10467)
);

INVx2_ASAP7_75t_L g10468 ( 
.A(n_9336),
.Y(n_10468)
);

OAI21x1_ASAP7_75t_L g10469 ( 
.A1(n_9551),
.A2(n_8964),
.B(n_8956),
.Y(n_10469)
);

INVx1_ASAP7_75t_L g10470 ( 
.A(n_9664),
.Y(n_10470)
);

NAND2xp5_ASAP7_75t_L g10471 ( 
.A(n_9906),
.B(n_8087),
.Y(n_10471)
);

AO21x2_ASAP7_75t_L g10472 ( 
.A1(n_9678),
.A2(n_8223),
.B(n_8172),
.Y(n_10472)
);

AO31x2_ASAP7_75t_L g10473 ( 
.A1(n_8980),
.A2(n_8944),
.A3(n_8968),
.B(n_8599),
.Y(n_10473)
);

HB1xp67_ASAP7_75t_L g10474 ( 
.A(n_9205),
.Y(n_10474)
);

HB1xp67_ASAP7_75t_L g10475 ( 
.A(n_9205),
.Y(n_10475)
);

INVx1_ASAP7_75t_L g10476 ( 
.A(n_9664),
.Y(n_10476)
);

NOR2xp33_ASAP7_75t_SL g10477 ( 
.A(n_9208),
.B(n_7808),
.Y(n_10477)
);

AND2x4_ASAP7_75t_L g10478 ( 
.A(n_9600),
.B(n_8250),
.Y(n_10478)
);

OAI21x1_ASAP7_75t_L g10479 ( 
.A1(n_9551),
.A2(n_8964),
.B(n_8956),
.Y(n_10479)
);

AND2x4_ASAP7_75t_L g10480 ( 
.A(n_9600),
.B(n_8250),
.Y(n_10480)
);

HB1xp67_ASAP7_75t_L g10481 ( 
.A(n_9205),
.Y(n_10481)
);

INVx3_ASAP7_75t_L g10482 ( 
.A(n_9600),
.Y(n_10482)
);

OAI21x1_ASAP7_75t_L g10483 ( 
.A1(n_9002),
.A2(n_8964),
.B(n_8956),
.Y(n_10483)
);

INVx1_ASAP7_75t_L g10484 ( 
.A(n_9673),
.Y(n_10484)
);

OAI21x1_ASAP7_75t_L g10485 ( 
.A1(n_9002),
.A2(n_8965),
.B(n_8964),
.Y(n_10485)
);

INVx2_ASAP7_75t_L g10486 ( 
.A(n_9439),
.Y(n_10486)
);

INVx1_ASAP7_75t_L g10487 ( 
.A(n_9673),
.Y(n_10487)
);

AOI221xp5_ASAP7_75t_L g10488 ( 
.A1(n_9206),
.A2(n_8746),
.B1(n_8751),
.B2(n_8153),
.C(n_8629),
.Y(n_10488)
);

AOI21xp33_ASAP7_75t_SL g10489 ( 
.A1(n_9897),
.A2(n_8427),
.B(n_8416),
.Y(n_10489)
);

OAI22xp5_ASAP7_75t_L g10490 ( 
.A1(n_10149),
.A2(n_8061),
.B1(n_7883),
.B2(n_8035),
.Y(n_10490)
);

OAI21xp5_ASAP7_75t_L g10491 ( 
.A1(n_9528),
.A2(n_8418),
.B(n_8259),
.Y(n_10491)
);

AND2x2_ASAP7_75t_L g10492 ( 
.A(n_9876),
.B(n_8019),
.Y(n_10492)
);

INVx1_ASAP7_75t_L g10493 ( 
.A(n_9673),
.Y(n_10493)
);

OAI21x1_ASAP7_75t_L g10494 ( 
.A1(n_9002),
.A2(n_8970),
.B(n_8965),
.Y(n_10494)
);

OAI21x1_ASAP7_75t_L g10495 ( 
.A1(n_9002),
.A2(n_8970),
.B(n_8965),
.Y(n_10495)
);

OAI21x1_ASAP7_75t_L g10496 ( 
.A1(n_9002),
.A2(n_8970),
.B(n_8965),
.Y(n_10496)
);

OA21x2_ASAP7_75t_L g10497 ( 
.A1(n_10101),
.A2(n_8970),
.B(n_8392),
.Y(n_10497)
);

AOI21xp5_ASAP7_75t_L g10498 ( 
.A1(n_10044),
.A2(n_8526),
.B(n_8433),
.Y(n_10498)
);

NAND2x1p5_ASAP7_75t_L g10499 ( 
.A(n_9110),
.B(n_8208),
.Y(n_10499)
);

INVx3_ASAP7_75t_L g10500 ( 
.A(n_9600),
.Y(n_10500)
);

INVx1_ASAP7_75t_L g10501 ( 
.A(n_9797),
.Y(n_10501)
);

AOI21xp5_ASAP7_75t_L g10502 ( 
.A1(n_10044),
.A2(n_8433),
.B(n_7756),
.Y(n_10502)
);

NAND2xp5_ASAP7_75t_L g10503 ( 
.A(n_9921),
.B(n_8094),
.Y(n_10503)
);

OAI21x1_ASAP7_75t_SL g10504 ( 
.A1(n_9032),
.A2(n_8436),
.B(n_8551),
.Y(n_10504)
);

NAND2xp5_ASAP7_75t_L g10505 ( 
.A(n_9921),
.B(n_10158),
.Y(n_10505)
);

INVx2_ASAP7_75t_L g10506 ( 
.A(n_9439),
.Y(n_10506)
);

OAI21x1_ASAP7_75t_L g10507 ( 
.A1(n_9273),
.A2(n_7692),
.B(n_8422),
.Y(n_10507)
);

INVx1_ASAP7_75t_L g10508 ( 
.A(n_9797),
.Y(n_10508)
);

OAI21x1_ASAP7_75t_L g10509 ( 
.A1(n_9273),
.A2(n_7692),
.B(n_8422),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_9797),
.Y(n_10510)
);

INVx2_ASAP7_75t_L g10511 ( 
.A(n_9439),
.Y(n_10511)
);

CKINVDCx5p33_ASAP7_75t_R g10512 ( 
.A(n_9739),
.Y(n_10512)
);

OA21x2_ASAP7_75t_L g10513 ( 
.A1(n_10101),
.A2(n_8392),
.B(n_8380),
.Y(n_10513)
);

CKINVDCx6p67_ASAP7_75t_R g10514 ( 
.A(n_9388),
.Y(n_10514)
);

INVx1_ASAP7_75t_L g10515 ( 
.A(n_9797),
.Y(n_10515)
);

INVx3_ASAP7_75t_L g10516 ( 
.A(n_9606),
.Y(n_10516)
);

AOI21xp5_ASAP7_75t_L g10517 ( 
.A1(n_10072),
.A2(n_7756),
.B(n_7763),
.Y(n_10517)
);

OAI21x1_ASAP7_75t_L g10518 ( 
.A1(n_9273),
.A2(n_7692),
.B(n_8422),
.Y(n_10518)
);

OAI21x1_ASAP7_75t_L g10519 ( 
.A1(n_9273),
.A2(n_7692),
.B(n_8422),
.Y(n_10519)
);

INVx1_ASAP7_75t_L g10520 ( 
.A(n_9810),
.Y(n_10520)
);

INVx1_ASAP7_75t_L g10521 ( 
.A(n_9810),
.Y(n_10521)
);

INVx2_ASAP7_75t_L g10522 ( 
.A(n_9439),
.Y(n_10522)
);

INVx1_ASAP7_75t_L g10523 ( 
.A(n_9810),
.Y(n_10523)
);

INVx1_ASAP7_75t_L g10524 ( 
.A(n_9810),
.Y(n_10524)
);

AND2x4_ASAP7_75t_L g10525 ( 
.A(n_9606),
.B(n_8250),
.Y(n_10525)
);

INVx1_ASAP7_75t_L g10526 ( 
.A(n_9815),
.Y(n_10526)
);

NAND2x1p5_ASAP7_75t_L g10527 ( 
.A(n_9110),
.B(n_8208),
.Y(n_10527)
);

NAND2xp5_ASAP7_75t_L g10528 ( 
.A(n_9921),
.B(n_8094),
.Y(n_10528)
);

OAI21xp5_ASAP7_75t_L g10529 ( 
.A1(n_9528),
.A2(n_8418),
.B(n_8464),
.Y(n_10529)
);

AOI22xp33_ASAP7_75t_L g10530 ( 
.A1(n_9544),
.A2(n_8194),
.B1(n_8071),
.B2(n_8180),
.Y(n_10530)
);

AO31x2_ASAP7_75t_L g10531 ( 
.A1(n_8980),
.A2(n_8944),
.A3(n_8968),
.B(n_8599),
.Y(n_10531)
);

OAI21x1_ASAP7_75t_L g10532 ( 
.A1(n_9791),
.A2(n_8424),
.B(n_8438),
.Y(n_10532)
);

OAI21x1_ASAP7_75t_L g10533 ( 
.A1(n_9791),
.A2(n_8424),
.B(n_8438),
.Y(n_10533)
);

OAI21x1_ASAP7_75t_L g10534 ( 
.A1(n_9791),
.A2(n_8424),
.B(n_8438),
.Y(n_10534)
);

OA21x2_ASAP7_75t_L g10535 ( 
.A1(n_10101),
.A2(n_10168),
.B(n_9700),
.Y(n_10535)
);

CKINVDCx5p33_ASAP7_75t_R g10536 ( 
.A(n_9739),
.Y(n_10536)
);

INVx1_ASAP7_75t_L g10537 ( 
.A(n_9815),
.Y(n_10537)
);

AOI21xp5_ASAP7_75t_L g10538 ( 
.A1(n_10072),
.A2(n_7756),
.B(n_7763),
.Y(n_10538)
);

OR2x6_ASAP7_75t_L g10539 ( 
.A(n_9441),
.B(n_8876),
.Y(n_10539)
);

AOI21x1_ASAP7_75t_L g10540 ( 
.A1(n_9815),
.A2(n_8697),
.B(n_8665),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_9815),
.Y(n_10541)
);

INVx2_ASAP7_75t_L g10542 ( 
.A(n_9439),
.Y(n_10542)
);

INVx1_ASAP7_75t_L g10543 ( 
.A(n_9818),
.Y(n_10543)
);

AOI21xp5_ASAP7_75t_L g10544 ( 
.A1(n_10072),
.A2(n_7756),
.B(n_8260),
.Y(n_10544)
);

NAND2x1p5_ASAP7_75t_L g10545 ( 
.A(n_9110),
.B(n_8208),
.Y(n_10545)
);

AO31x2_ASAP7_75t_L g10546 ( 
.A1(n_9871),
.A2(n_8968),
.A3(n_8777),
.B(n_8782),
.Y(n_10546)
);

AND2x2_ASAP7_75t_L g10547 ( 
.A(n_9880),
.B(n_9346),
.Y(n_10547)
);

OAI21x1_ASAP7_75t_L g10548 ( 
.A1(n_9791),
.A2(n_8424),
.B(n_8508),
.Y(n_10548)
);

INVx2_ASAP7_75t_L g10549 ( 
.A(n_9439),
.Y(n_10549)
);

NAND2x1p5_ASAP7_75t_L g10550 ( 
.A(n_9110),
.B(n_8208),
.Y(n_10550)
);

OAI21x1_ASAP7_75t_L g10551 ( 
.A1(n_9833),
.A2(n_8508),
.B(n_8392),
.Y(n_10551)
);

OAI21xp33_ASAP7_75t_L g10552 ( 
.A1(n_9544),
.A2(n_8122),
.B(n_8112),
.Y(n_10552)
);

AND2x2_ASAP7_75t_L g10553 ( 
.A(n_9880),
.B(n_8019),
.Y(n_10553)
);

NAND2xp5_ASAP7_75t_L g10554 ( 
.A(n_10158),
.B(n_8775),
.Y(n_10554)
);

AND2x2_ASAP7_75t_L g10555 ( 
.A(n_9880),
.B(n_8093),
.Y(n_10555)
);

AOI21xp5_ASAP7_75t_L g10556 ( 
.A1(n_9898),
.A2(n_9032),
.B(n_9995),
.Y(n_10556)
);

AO31x2_ASAP7_75t_L g10557 ( 
.A1(n_9871),
.A2(n_8968),
.A3(n_8777),
.B(n_8782),
.Y(n_10557)
);

NOR2xp33_ASAP7_75t_L g10558 ( 
.A(n_9277),
.B(n_7836),
.Y(n_10558)
);

OAI21xp5_ASAP7_75t_L g10559 ( 
.A1(n_9528),
.A2(n_8418),
.B(n_8464),
.Y(n_10559)
);

OAI21x1_ASAP7_75t_L g10560 ( 
.A1(n_9833),
.A2(n_8508),
.B(n_8392),
.Y(n_10560)
);

OAI21xp5_ASAP7_75t_L g10561 ( 
.A1(n_9528),
.A2(n_8464),
.B(n_8640),
.Y(n_10561)
);

OAI21x1_ASAP7_75t_L g10562 ( 
.A1(n_9833),
.A2(n_8380),
.B(n_8476),
.Y(n_10562)
);

INVx2_ASAP7_75t_L g10563 ( 
.A(n_9439),
.Y(n_10563)
);

A2O1A1Ixp33_ASAP7_75t_L g10564 ( 
.A1(n_9966),
.A2(n_8402),
.B(n_7765),
.C(n_7977),
.Y(n_10564)
);

INVx1_ASAP7_75t_L g10565 ( 
.A(n_9818),
.Y(n_10565)
);

OAI21xp5_ASAP7_75t_L g10566 ( 
.A1(n_9119),
.A2(n_8464),
.B(n_8640),
.Y(n_10566)
);

NOR2xp33_ASAP7_75t_L g10567 ( 
.A(n_9277),
.B(n_8423),
.Y(n_10567)
);

NAND2x1p5_ASAP7_75t_L g10568 ( 
.A(n_9370),
.B(n_8067),
.Y(n_10568)
);

OA21x2_ASAP7_75t_L g10569 ( 
.A1(n_10168),
.A2(n_8380),
.B(n_8476),
.Y(n_10569)
);

OR2x2_ASAP7_75t_L g10570 ( 
.A(n_9889),
.B(n_8384),
.Y(n_10570)
);

AO31x2_ASAP7_75t_L g10571 ( 
.A1(n_9871),
.A2(n_8769),
.A3(n_8827),
.B(n_8388),
.Y(n_10571)
);

OR2x2_ASAP7_75t_L g10572 ( 
.A(n_9889),
.B(n_8384),
.Y(n_10572)
);

NAND2xp5_ASAP7_75t_L g10573 ( 
.A(n_10158),
.B(n_8775),
.Y(n_10573)
);

BUFx2_ASAP7_75t_L g10574 ( 
.A(n_9975),
.Y(n_10574)
);

INVx2_ASAP7_75t_L g10575 ( 
.A(n_9439),
.Y(n_10575)
);

AND2x4_ASAP7_75t_L g10576 ( 
.A(n_9606),
.B(n_8250),
.Y(n_10576)
);

AO21x2_ASAP7_75t_L g10577 ( 
.A1(n_9682),
.A2(n_9700),
.B(n_10168),
.Y(n_10577)
);

INVx2_ASAP7_75t_L g10578 ( 
.A(n_9439),
.Y(n_10578)
);

OAI21x1_ASAP7_75t_L g10579 ( 
.A1(n_9833),
.A2(n_8380),
.B(n_8476),
.Y(n_10579)
);

OAI21x1_ASAP7_75t_L g10580 ( 
.A1(n_9069),
.A2(n_8476),
.B(n_8741),
.Y(n_10580)
);

BUFx2_ASAP7_75t_R g10581 ( 
.A(n_9056),
.Y(n_10581)
);

NOR2xp33_ASAP7_75t_SL g10582 ( 
.A(n_9208),
.B(n_8298),
.Y(n_10582)
);

NAND2x1p5_ASAP7_75t_L g10583 ( 
.A(n_9370),
.B(n_9229),
.Y(n_10583)
);

INVx1_ASAP7_75t_L g10584 ( 
.A(n_9818),
.Y(n_10584)
);

INVx1_ASAP7_75t_SL g10585 ( 
.A(n_9134),
.Y(n_10585)
);

CKINVDCx11_ASAP7_75t_R g10586 ( 
.A(n_9388),
.Y(n_10586)
);

NAND2xp5_ASAP7_75t_L g10587 ( 
.A(n_10066),
.B(n_8793),
.Y(n_10587)
);

NAND2xp5_ASAP7_75t_SL g10588 ( 
.A(n_9208),
.B(n_9255),
.Y(n_10588)
);

INVx2_ASAP7_75t_L g10589 ( 
.A(n_9447),
.Y(n_10589)
);

INVx2_ASAP7_75t_L g10590 ( 
.A(n_9447),
.Y(n_10590)
);

AOI21x1_ASAP7_75t_L g10591 ( 
.A1(n_9818),
.A2(n_8697),
.B(n_7707),
.Y(n_10591)
);

AND2x2_ASAP7_75t_L g10592 ( 
.A(n_9880),
.B(n_8093),
.Y(n_10592)
);

OR2x2_ASAP7_75t_L g10593 ( 
.A(n_9889),
.B(n_8384),
.Y(n_10593)
);

INVx1_ASAP7_75t_L g10594 ( 
.A(n_9820),
.Y(n_10594)
);

INVx1_ASAP7_75t_L g10595 ( 
.A(n_9820),
.Y(n_10595)
);

INVx2_ASAP7_75t_L g10596 ( 
.A(n_9447),
.Y(n_10596)
);

BUFx3_ASAP7_75t_L g10597 ( 
.A(n_9073),
.Y(n_10597)
);

OR2x6_ASAP7_75t_L g10598 ( 
.A(n_9441),
.B(n_8876),
.Y(n_10598)
);

INVx2_ASAP7_75t_L g10599 ( 
.A(n_9447),
.Y(n_10599)
);

CKINVDCx12_ASAP7_75t_R g10600 ( 
.A(n_10146),
.Y(n_10600)
);

INVx1_ASAP7_75t_L g10601 ( 
.A(n_9820),
.Y(n_10601)
);

BUFx3_ASAP7_75t_L g10602 ( 
.A(n_9073),
.Y(n_10602)
);

OAI21x1_ASAP7_75t_L g10603 ( 
.A1(n_9069),
.A2(n_8741),
.B(n_8748),
.Y(n_10603)
);

BUFx3_ASAP7_75t_L g10604 ( 
.A(n_9073),
.Y(n_10604)
);

NOR2x1_ASAP7_75t_SL g10605 ( 
.A(n_9272),
.B(n_8044),
.Y(n_10605)
);

INVx2_ASAP7_75t_L g10606 ( 
.A(n_9447),
.Y(n_10606)
);

INVx2_ASAP7_75t_SL g10607 ( 
.A(n_9441),
.Y(n_10607)
);

INVx1_ASAP7_75t_L g10608 ( 
.A(n_9820),
.Y(n_10608)
);

INVx1_ASAP7_75t_L g10609 ( 
.A(n_9824),
.Y(n_10609)
);

AO21x2_ASAP7_75t_L g10610 ( 
.A1(n_9682),
.A2(n_8172),
.B(n_8130),
.Y(n_10610)
);

OAI21xp5_ASAP7_75t_L g10611 ( 
.A1(n_9119),
.A2(n_8122),
.B(n_8112),
.Y(n_10611)
);

HB1xp67_ASAP7_75t_L g10612 ( 
.A(n_9205),
.Y(n_10612)
);

AND2x4_ASAP7_75t_L g10613 ( 
.A(n_9606),
.B(n_8250),
.Y(n_10613)
);

AO21x2_ASAP7_75t_L g10614 ( 
.A1(n_9682),
.A2(n_8130),
.B(n_8622),
.Y(n_10614)
);

INVx1_ASAP7_75t_L g10615 ( 
.A(n_9824),
.Y(n_10615)
);

OA21x2_ASAP7_75t_L g10616 ( 
.A1(n_9700),
.A2(n_8622),
.B(n_8616),
.Y(n_10616)
);

A2O1A1Ixp33_ASAP7_75t_L g10617 ( 
.A1(n_9966),
.A2(n_8402),
.B(n_7765),
.C(n_7977),
.Y(n_10617)
);

AOI21xp33_ASAP7_75t_L g10618 ( 
.A1(n_9544),
.A2(n_8379),
.B(n_8180),
.Y(n_10618)
);

BUFx6f_ASAP7_75t_L g10619 ( 
.A(n_9060),
.Y(n_10619)
);

NOR2xp33_ASAP7_75t_L g10620 ( 
.A(n_9277),
.B(n_8423),
.Y(n_10620)
);

OAI21x1_ASAP7_75t_L g10621 ( 
.A1(n_9069),
.A2(n_8741),
.B(n_8748),
.Y(n_10621)
);

INVx1_ASAP7_75t_L g10622 ( 
.A(n_9824),
.Y(n_10622)
);

AND2x2_ASAP7_75t_L g10623 ( 
.A(n_9880),
.B(n_8093),
.Y(n_10623)
);

OAI21x1_ASAP7_75t_L g10624 ( 
.A1(n_9069),
.A2(n_8748),
.B(n_8692),
.Y(n_10624)
);

BUFx8_ASAP7_75t_L g10625 ( 
.A(n_9148),
.Y(n_10625)
);

OR2x6_ASAP7_75t_L g10626 ( 
.A(n_9441),
.B(n_8281),
.Y(n_10626)
);

NAND3xp33_ASAP7_75t_L g10627 ( 
.A(n_9969),
.B(n_8153),
.C(n_8751),
.Y(n_10627)
);

AND2x4_ASAP7_75t_L g10628 ( 
.A(n_9606),
.B(n_9654),
.Y(n_10628)
);

OAI21x1_ASAP7_75t_L g10629 ( 
.A1(n_9069),
.A2(n_8748),
.B(n_8692),
.Y(n_10629)
);

OAI21x1_ASAP7_75t_L g10630 ( 
.A1(n_9318),
.A2(n_9080),
.B(n_9557),
.Y(n_10630)
);

HB1xp67_ASAP7_75t_L g10631 ( 
.A(n_9205),
.Y(n_10631)
);

OR2x6_ASAP7_75t_L g10632 ( 
.A(n_9441),
.B(n_8369),
.Y(n_10632)
);

AOI21xp5_ASAP7_75t_L g10633 ( 
.A1(n_9032),
.A2(n_10042),
.B(n_9995),
.Y(n_10633)
);

INVx2_ASAP7_75t_L g10634 ( 
.A(n_9336),
.Y(n_10634)
);

INVxp67_ASAP7_75t_L g10635 ( 
.A(n_9962),
.Y(n_10635)
);

INVx2_ASAP7_75t_L g10636 ( 
.A(n_9336),
.Y(n_10636)
);

NOR2xp67_ASAP7_75t_L g10637 ( 
.A(n_9467),
.B(n_8044),
.Y(n_10637)
);

BUFx4f_ASAP7_75t_SL g10638 ( 
.A(n_9388),
.Y(n_10638)
);

OAI21x1_ASAP7_75t_L g10639 ( 
.A1(n_9318),
.A2(n_8692),
.B(n_8691),
.Y(n_10639)
);

INVx1_ASAP7_75t_L g10640 ( 
.A(n_9824),
.Y(n_10640)
);

HB1xp67_ASAP7_75t_L g10641 ( 
.A(n_9205),
.Y(n_10641)
);

AND2x2_ASAP7_75t_L g10642 ( 
.A(n_9346),
.B(n_8093),
.Y(n_10642)
);

AND2x2_ASAP7_75t_L g10643 ( 
.A(n_9346),
.B(n_7894),
.Y(n_10643)
);

INVx3_ASAP7_75t_SL g10644 ( 
.A(n_9025),
.Y(n_10644)
);

OAI21x1_ASAP7_75t_L g10645 ( 
.A1(n_9318),
.A2(n_9080),
.B(n_9557),
.Y(n_10645)
);

INVx2_ASAP7_75t_L g10646 ( 
.A(n_9336),
.Y(n_10646)
);

AOI22xp5_ASAP7_75t_L g10647 ( 
.A1(n_9277),
.A2(n_8194),
.B1(n_8377),
.B2(n_7772),
.Y(n_10647)
);

A2O1A1Ixp33_ASAP7_75t_L g10648 ( 
.A1(n_9966),
.A2(n_8459),
.B(n_7687),
.C(n_8264),
.Y(n_10648)
);

INVx1_ASAP7_75t_L g10649 ( 
.A(n_9825),
.Y(n_10649)
);

INVx2_ASAP7_75t_L g10650 ( 
.A(n_9336),
.Y(n_10650)
);

NAND2x1p5_ASAP7_75t_L g10651 ( 
.A(n_9370),
.B(n_8067),
.Y(n_10651)
);

AOI21xp5_ASAP7_75t_L g10652 ( 
.A1(n_9995),
.A2(n_8260),
.B(n_8271),
.Y(n_10652)
);

OAI21x1_ASAP7_75t_L g10653 ( 
.A1(n_9318),
.A2(n_9080),
.B(n_9557),
.Y(n_10653)
);

AO31x2_ASAP7_75t_L g10654 ( 
.A1(n_9871),
.A2(n_8769),
.A3(n_8827),
.B(n_8388),
.Y(n_10654)
);

AND2x2_ASAP7_75t_L g10655 ( 
.A(n_9346),
.B(n_7894),
.Y(n_10655)
);

INVx1_ASAP7_75t_L g10656 ( 
.A(n_9825),
.Y(n_10656)
);

AO21x2_ASAP7_75t_L g10657 ( 
.A1(n_8982),
.A2(n_8447),
.B(n_8445),
.Y(n_10657)
);

OAI22xp5_ASAP7_75t_L g10658 ( 
.A1(n_10149),
.A2(n_8035),
.B1(n_7883),
.B2(n_8174),
.Y(n_10658)
);

OAI21x1_ASAP7_75t_L g10659 ( 
.A1(n_9318),
.A2(n_8739),
.B(n_8691),
.Y(n_10659)
);

INVx2_ASAP7_75t_L g10660 ( 
.A(n_9336),
.Y(n_10660)
);

HB1xp67_ASAP7_75t_L g10661 ( 
.A(n_9205),
.Y(n_10661)
);

INVx1_ASAP7_75t_L g10662 ( 
.A(n_9825),
.Y(n_10662)
);

OAI21x1_ASAP7_75t_L g10663 ( 
.A1(n_9080),
.A2(n_8739),
.B(n_8691),
.Y(n_10663)
);

OAI22xp33_ASAP7_75t_L g10664 ( 
.A1(n_10071),
.A2(n_7772),
.B1(n_8174),
.B2(n_8224),
.Y(n_10664)
);

BUFx3_ASAP7_75t_L g10665 ( 
.A(n_9131),
.Y(n_10665)
);

NOR2xp67_ASAP7_75t_L g10666 ( 
.A(n_9467),
.B(n_8044),
.Y(n_10666)
);

INVx1_ASAP7_75t_SL g10667 ( 
.A(n_9134),
.Y(n_10667)
);

OAI21x1_ASAP7_75t_L g10668 ( 
.A1(n_9080),
.A2(n_8739),
.B(n_8265),
.Y(n_10668)
);

OR2x6_ASAP7_75t_L g10669 ( 
.A(n_9441),
.B(n_8369),
.Y(n_10669)
);

OAI21x1_ASAP7_75t_L g10670 ( 
.A1(n_9557),
.A2(n_8265),
.B(n_8262),
.Y(n_10670)
);

NAND2xp5_ASAP7_75t_L g10671 ( 
.A(n_10066),
.B(n_8793),
.Y(n_10671)
);

OAI21x1_ASAP7_75t_L g10672 ( 
.A1(n_9557),
.A2(n_10136),
.B(n_10129),
.Y(n_10672)
);

INVx1_ASAP7_75t_L g10673 ( 
.A(n_9825),
.Y(n_10673)
);

INVx1_ASAP7_75t_L g10674 ( 
.A(n_9832),
.Y(n_10674)
);

INVx2_ASAP7_75t_L g10675 ( 
.A(n_9447),
.Y(n_10675)
);

NOR2xp67_ASAP7_75t_L g10676 ( 
.A(n_8995),
.B(n_8168),
.Y(n_10676)
);

OAI21x1_ASAP7_75t_L g10677 ( 
.A1(n_10136),
.A2(n_10129),
.B(n_10126),
.Y(n_10677)
);

BUFx2_ASAP7_75t_L g10678 ( 
.A(n_9606),
.Y(n_10678)
);

OAI21x1_ASAP7_75t_L g10679 ( 
.A1(n_10136),
.A2(n_8262),
.B(n_8864),
.Y(n_10679)
);

OAI21x1_ASAP7_75t_L g10680 ( 
.A1(n_10136),
.A2(n_8865),
.B(n_8864),
.Y(n_10680)
);

NOR2xp67_ASAP7_75t_L g10681 ( 
.A(n_8995),
.B(n_8168),
.Y(n_10681)
);

INVx1_ASAP7_75t_L g10682 ( 
.A(n_9832),
.Y(n_10682)
);

NOR2xp33_ASAP7_75t_L g10683 ( 
.A(n_9970),
.B(n_7897),
.Y(n_10683)
);

NOR2x1_ASAP7_75t_R g10684 ( 
.A(n_9388),
.B(n_8338),
.Y(n_10684)
);

INVxp67_ASAP7_75t_SL g10685 ( 
.A(n_9414),
.Y(n_10685)
);

CKINVDCx5p33_ASAP7_75t_R g10686 ( 
.A(n_10152),
.Y(n_10686)
);

OAI21x1_ASAP7_75t_L g10687 ( 
.A1(n_10136),
.A2(n_8865),
.B(n_8864),
.Y(n_10687)
);

NAND2x1p5_ASAP7_75t_L g10688 ( 
.A(n_9370),
.B(n_8067),
.Y(n_10688)
);

INVx3_ASAP7_75t_L g10689 ( 
.A(n_9654),
.Y(n_10689)
);

AOI21xp5_ASAP7_75t_L g10690 ( 
.A1(n_10042),
.A2(n_8271),
.B(n_8264),
.Y(n_10690)
);

OAI21x1_ASAP7_75t_L g10691 ( 
.A1(n_10126),
.A2(n_8865),
.B(n_8864),
.Y(n_10691)
);

OAI21xp5_ASAP7_75t_L g10692 ( 
.A1(n_9119),
.A2(n_8379),
.B(n_8109),
.Y(n_10692)
);

NAND2xp5_ASAP7_75t_L g10693 ( 
.A(n_10066),
.B(n_8795),
.Y(n_10693)
);

NAND4xp25_ASAP7_75t_L g10694 ( 
.A(n_9969),
.B(n_10020),
.C(n_10151),
.D(n_9950),
.Y(n_10694)
);

INVx1_ASAP7_75t_L g10695 ( 
.A(n_9832),
.Y(n_10695)
);

CKINVDCx6p67_ASAP7_75t_R g10696 ( 
.A(n_9388),
.Y(n_10696)
);

OAI221xp5_ASAP7_75t_SL g10697 ( 
.A1(n_10149),
.A2(n_8224),
.B1(n_8377),
.B2(n_8109),
.C(n_8174),
.Y(n_10697)
);

NAND2x1p5_ASAP7_75t_L g10698 ( 
.A(n_9370),
.B(n_8435),
.Y(n_10698)
);

OAI21x1_ASAP7_75t_L g10699 ( 
.A1(n_10126),
.A2(n_8865),
.B(n_8447),
.Y(n_10699)
);

OAI21x1_ASAP7_75t_L g10700 ( 
.A1(n_10126),
.A2(n_8456),
.B(n_8445),
.Y(n_10700)
);

INVx1_ASAP7_75t_L g10701 ( 
.A(n_9832),
.Y(n_10701)
);

AOI21xp5_ASAP7_75t_L g10702 ( 
.A1(n_10042),
.A2(n_8553),
.B(n_8543),
.Y(n_10702)
);

NAND2xp5_ASAP7_75t_L g10703 ( 
.A(n_10074),
.B(n_8795),
.Y(n_10703)
);

AO31x2_ASAP7_75t_L g10704 ( 
.A1(n_9871),
.A2(n_8156),
.A3(n_8840),
.B(n_8834),
.Y(n_10704)
);

A2O1A1Ixp33_ASAP7_75t_L g10705 ( 
.A1(n_9966),
.A2(n_10068),
.B(n_10045),
.C(n_9942),
.Y(n_10705)
);

INVx1_ASAP7_75t_L g10706 ( 
.A(n_9839),
.Y(n_10706)
);

AO21x2_ASAP7_75t_L g10707 ( 
.A1(n_8982),
.A2(n_8469),
.B(n_8456),
.Y(n_10707)
);

CKINVDCx16_ASAP7_75t_R g10708 ( 
.A(n_9201),
.Y(n_10708)
);

OA21x2_ASAP7_75t_L g10709 ( 
.A1(n_9881),
.A2(n_8616),
.B(n_8186),
.Y(n_10709)
);

AO21x2_ASAP7_75t_L g10710 ( 
.A1(n_8982),
.A2(n_8474),
.B(n_8469),
.Y(n_10710)
);

BUFx6f_ASAP7_75t_L g10711 ( 
.A(n_9060),
.Y(n_10711)
);

OAI21x1_ASAP7_75t_L g10712 ( 
.A1(n_10126),
.A2(n_8477),
.B(n_8474),
.Y(n_10712)
);

NAND2xp5_ASAP7_75t_L g10713 ( 
.A(n_10074),
.B(n_10174),
.Y(n_10713)
);

NAND2xp5_ASAP7_75t_L g10714 ( 
.A(n_10074),
.B(n_7993),
.Y(n_10714)
);

NAND2x1p5_ASAP7_75t_L g10715 ( 
.A(n_9370),
.B(n_8435),
.Y(n_10715)
);

A2O1A1Ixp33_ASAP7_75t_L g10716 ( 
.A1(n_10045),
.A2(n_8459),
.B(n_7687),
.C(n_8224),
.Y(n_10716)
);

INVx2_ASAP7_75t_L g10717 ( 
.A(n_9336),
.Y(n_10717)
);

OA21x2_ASAP7_75t_L g10718 ( 
.A1(n_9881),
.A2(n_8616),
.B(n_8186),
.Y(n_10718)
);

INVx1_ASAP7_75t_L g10719 ( 
.A(n_9839),
.Y(n_10719)
);

OAI21xp33_ASAP7_75t_SL g10720 ( 
.A1(n_9922),
.A2(n_8035),
.B(n_7883),
.Y(n_10720)
);

AOI22x1_ASAP7_75t_L g10721 ( 
.A1(n_9922),
.A2(n_8180),
.B1(n_8523),
.B2(n_8416),
.Y(n_10721)
);

INVx2_ASAP7_75t_L g10722 ( 
.A(n_9337),
.Y(n_10722)
);

OAI21x1_ASAP7_75t_L g10723 ( 
.A1(n_10129),
.A2(n_8488),
.B(n_8477),
.Y(n_10723)
);

NOR2xp67_ASAP7_75t_L g10724 ( 
.A(n_8995),
.B(n_8168),
.Y(n_10724)
);

INVx3_ASAP7_75t_L g10725 ( 
.A(n_9654),
.Y(n_10725)
);

AOI22xp33_ASAP7_75t_L g10726 ( 
.A1(n_10020),
.A2(n_9950),
.B1(n_9904),
.B2(n_9998),
.Y(n_10726)
);

NAND2xp5_ASAP7_75t_L g10727 ( 
.A(n_10174),
.B(n_7993),
.Y(n_10727)
);

CKINVDCx12_ASAP7_75t_R g10728 ( 
.A(n_10146),
.Y(n_10728)
);

CKINVDCx11_ASAP7_75t_R g10729 ( 
.A(n_9489),
.Y(n_10729)
);

NAND2xp5_ASAP7_75t_L g10730 ( 
.A(n_10174),
.B(n_7994),
.Y(n_10730)
);

OAI21x1_ASAP7_75t_L g10731 ( 
.A1(n_10129),
.A2(n_8494),
.B(n_8488),
.Y(n_10731)
);

AOI211xp5_ASAP7_75t_L g10732 ( 
.A1(n_9948),
.A2(n_8327),
.B(n_8216),
.C(n_8770),
.Y(n_10732)
);

OAI21x1_ASAP7_75t_L g10733 ( 
.A1(n_10129),
.A2(n_8502),
.B(n_8494),
.Y(n_10733)
);

INVx4_ASAP7_75t_L g10734 ( 
.A(n_9148),
.Y(n_10734)
);

INVx1_ASAP7_75t_L g10735 ( 
.A(n_9839),
.Y(n_10735)
);

BUFx12f_ASAP7_75t_L g10736 ( 
.A(n_9489),
.Y(n_10736)
);

AND2x2_ASAP7_75t_L g10737 ( 
.A(n_9403),
.B(n_7948),
.Y(n_10737)
);

INVx1_ASAP7_75t_L g10738 ( 
.A(n_9839),
.Y(n_10738)
);

O2A1O1Ixp33_ASAP7_75t_L g10739 ( 
.A1(n_10020),
.A2(n_8216),
.B(n_8463),
.C(n_8327),
.Y(n_10739)
);

OA21x2_ASAP7_75t_L g10740 ( 
.A1(n_9881),
.A2(n_8616),
.B(n_8185),
.Y(n_10740)
);

AOI21x1_ASAP7_75t_L g10741 ( 
.A1(n_9840),
.A2(n_7707),
.B(n_8082),
.Y(n_10741)
);

AND2x2_ASAP7_75t_L g10742 ( 
.A(n_9403),
.B(n_9451),
.Y(n_10742)
);

INVx2_ASAP7_75t_L g10743 ( 
.A(n_9447),
.Y(n_10743)
);

INVx1_ASAP7_75t_L g10744 ( 
.A(n_9840),
.Y(n_10744)
);

INVx2_ASAP7_75t_L g10745 ( 
.A(n_9447),
.Y(n_10745)
);

AO21x2_ASAP7_75t_L g10746 ( 
.A1(n_9011),
.A2(n_8502),
.B(n_8507),
.Y(n_10746)
);

INVx1_ASAP7_75t_L g10747 ( 
.A(n_9840),
.Y(n_10747)
);

OA21x2_ASAP7_75t_L g10748 ( 
.A1(n_9972),
.A2(n_10073),
.B(n_10031),
.Y(n_10748)
);

AO21x2_ASAP7_75t_L g10749 ( 
.A1(n_9011),
.A2(n_8507),
.B(n_8554),
.Y(n_10749)
);

AO31x2_ASAP7_75t_L g10750 ( 
.A1(n_9037),
.A2(n_8156),
.A3(n_8840),
.B(n_8834),
.Y(n_10750)
);

OAI21x1_ASAP7_75t_L g10751 ( 
.A1(n_10144),
.A2(n_8724),
.B(n_8723),
.Y(n_10751)
);

NOR3xp33_ASAP7_75t_L g10752 ( 
.A(n_9948),
.B(n_9942),
.C(n_9922),
.Y(n_10752)
);

BUFx6f_ASAP7_75t_L g10753 ( 
.A(n_9060),
.Y(n_10753)
);

AO31x2_ASAP7_75t_L g10754 ( 
.A1(n_9037),
.A2(n_8527),
.A3(n_8874),
.B(n_8364),
.Y(n_10754)
);

OAI21x1_ASAP7_75t_L g10755 ( 
.A1(n_10144),
.A2(n_8724),
.B(n_8723),
.Y(n_10755)
);

OAI21x1_ASAP7_75t_L g10756 ( 
.A1(n_10144),
.A2(n_8724),
.B(n_8723),
.Y(n_10756)
);

OAI21x1_ASAP7_75t_L g10757 ( 
.A1(n_10144),
.A2(n_8724),
.B(n_8723),
.Y(n_10757)
);

OR2x2_ASAP7_75t_L g10758 ( 
.A(n_9972),
.B(n_8384),
.Y(n_10758)
);

BUFx8_ASAP7_75t_L g10759 ( 
.A(n_9148),
.Y(n_10759)
);

AO21x2_ASAP7_75t_L g10760 ( 
.A1(n_9011),
.A2(n_8554),
.B(n_8559),
.Y(n_10760)
);

OAI21x1_ASAP7_75t_L g10761 ( 
.A1(n_10144),
.A2(n_8869),
.B(n_8868),
.Y(n_10761)
);

AO21x2_ASAP7_75t_L g10762 ( 
.A1(n_9424),
.A2(n_8559),
.B(n_8605),
.Y(n_10762)
);

AOI21xp5_ASAP7_75t_L g10763 ( 
.A1(n_9942),
.A2(n_8553),
.B(n_8543),
.Y(n_10763)
);

OAI21x1_ASAP7_75t_SL g10764 ( 
.A1(n_9904),
.A2(n_8436),
.B(n_8551),
.Y(n_10764)
);

OAI22xp5_ASAP7_75t_L g10765 ( 
.A1(n_10071),
.A2(n_8377),
.B1(n_8339),
.B2(n_8180),
.Y(n_10765)
);

OA21x2_ASAP7_75t_L g10766 ( 
.A1(n_9972),
.A2(n_8185),
.B(n_8496),
.Y(n_10766)
);

OAI21x1_ASAP7_75t_L g10767 ( 
.A1(n_9226),
.A2(n_8869),
.B(n_8868),
.Y(n_10767)
);

AOI21xp5_ASAP7_75t_L g10768 ( 
.A1(n_10138),
.A2(n_8400),
.B(n_8180),
.Y(n_10768)
);

NAND2x1p5_ASAP7_75t_L g10769 ( 
.A(n_9370),
.B(n_8300),
.Y(n_10769)
);

BUFx4f_ASAP7_75t_SL g10770 ( 
.A(n_9489),
.Y(n_10770)
);

OAI21x1_ASAP7_75t_L g10771 ( 
.A1(n_9226),
.A2(n_8879),
.B(n_8877),
.Y(n_10771)
);

CKINVDCx5p33_ASAP7_75t_R g10772 ( 
.A(n_10152),
.Y(n_10772)
);

AO21x2_ASAP7_75t_L g10773 ( 
.A1(n_9424),
.A2(n_8605),
.B(n_8188),
.Y(n_10773)
);

OAI21x1_ASAP7_75t_L g10774 ( 
.A1(n_9226),
.A2(n_8879),
.B(n_8877),
.Y(n_10774)
);

INVx2_ASAP7_75t_L g10775 ( 
.A(n_9447),
.Y(n_10775)
);

INVx1_ASAP7_75t_L g10776 ( 
.A(n_9840),
.Y(n_10776)
);

AND2x4_ASAP7_75t_L g10777 ( 
.A(n_9654),
.B(n_8250),
.Y(n_10777)
);

OAI21x1_ASAP7_75t_SL g10778 ( 
.A1(n_9904),
.A2(n_8168),
.B(n_8285),
.Y(n_10778)
);

INVx3_ASAP7_75t_L g10779 ( 
.A(n_9654),
.Y(n_10779)
);

AO21x1_ASAP7_75t_L g10780 ( 
.A1(n_10045),
.A2(n_8511),
.B(n_8911),
.Y(n_10780)
);

OAI21x1_ASAP7_75t_L g10781 ( 
.A1(n_9226),
.A2(n_8886),
.B(n_8851),
.Y(n_10781)
);

AO31x2_ASAP7_75t_L g10782 ( 
.A1(n_9037),
.A2(n_8527),
.A3(n_8874),
.B(n_8364),
.Y(n_10782)
);

NAND2xp5_ASAP7_75t_L g10783 ( 
.A(n_10134),
.B(n_7994),
.Y(n_10783)
);

HB1xp67_ASAP7_75t_L g10784 ( 
.A(n_9205),
.Y(n_10784)
);

INVx2_ASAP7_75t_L g10785 ( 
.A(n_9462),
.Y(n_10785)
);

INVx1_ASAP7_75t_L g10786 ( 
.A(n_9846),
.Y(n_10786)
);

AO31x2_ASAP7_75t_L g10787 ( 
.A1(n_9414),
.A2(n_8527),
.A3(n_8874),
.B(n_8364),
.Y(n_10787)
);

BUFx2_ASAP7_75t_R g10788 ( 
.A(n_9219),
.Y(n_10788)
);

INVx1_ASAP7_75t_L g10789 ( 
.A(n_9846),
.Y(n_10789)
);

INVx2_ASAP7_75t_SL g10790 ( 
.A(n_9441),
.Y(n_10790)
);

OA21x2_ASAP7_75t_L g10791 ( 
.A1(n_9972),
.A2(n_8496),
.B(n_8851),
.Y(n_10791)
);

AND2x2_ASAP7_75t_L g10792 ( 
.A(n_9403),
.B(n_7948),
.Y(n_10792)
);

CKINVDCx11_ASAP7_75t_R g10793 ( 
.A(n_9489),
.Y(n_10793)
);

AND2x4_ASAP7_75t_L g10794 ( 
.A(n_9654),
.B(n_8279),
.Y(n_10794)
);

AOI21x1_ASAP7_75t_L g10795 ( 
.A1(n_9846),
.A2(n_7707),
.B(n_8082),
.Y(n_10795)
);

HB1xp67_ASAP7_75t_L g10796 ( 
.A(n_9200),
.Y(n_10796)
);

NAND2xp5_ASAP7_75t_L g10797 ( 
.A(n_10134),
.B(n_8001),
.Y(n_10797)
);

INVx2_ASAP7_75t_L g10798 ( 
.A(n_9462),
.Y(n_10798)
);

NAND2x1p5_ASAP7_75t_L g10799 ( 
.A(n_9370),
.B(n_8300),
.Y(n_10799)
);

OAI21xp5_ASAP7_75t_L g10800 ( 
.A1(n_9948),
.A2(n_8463),
.B(n_8389),
.Y(n_10800)
);

INVx2_ASAP7_75t_SL g10801 ( 
.A(n_9577),
.Y(n_10801)
);

OAI21x1_ASAP7_75t_L g10802 ( 
.A1(n_9226),
.A2(n_8886),
.B(n_8580),
.Y(n_10802)
);

OA21x2_ASAP7_75t_L g10803 ( 
.A1(n_9972),
.A2(n_8188),
.B(n_8187),
.Y(n_10803)
);

OA21x2_ASAP7_75t_L g10804 ( 
.A1(n_10031),
.A2(n_8187),
.B(n_8627),
.Y(n_10804)
);

OA21x2_ASAP7_75t_L g10805 ( 
.A1(n_10031),
.A2(n_8628),
.B(n_8627),
.Y(n_10805)
);

NOR2xp33_ASAP7_75t_L g10806 ( 
.A(n_9970),
.B(n_7897),
.Y(n_10806)
);

OA21x2_ASAP7_75t_L g10807 ( 
.A1(n_10031),
.A2(n_8630),
.B(n_8628),
.Y(n_10807)
);

AO21x2_ASAP7_75t_L g10808 ( 
.A1(n_9424),
.A2(n_8609),
.B(n_8387),
.Y(n_10808)
);

NAND2xp5_ASAP7_75t_L g10809 ( 
.A(n_10134),
.B(n_10165),
.Y(n_10809)
);

BUFx12f_ASAP7_75t_SL g10810 ( 
.A(n_8988),
.Y(n_10810)
);

AOI21xp5_ASAP7_75t_L g10811 ( 
.A1(n_10138),
.A2(n_8400),
.B(n_7737),
.Y(n_10811)
);

CKINVDCx20_ASAP7_75t_R g10812 ( 
.A(n_9149),
.Y(n_10812)
);

OA21x2_ASAP7_75t_L g10813 ( 
.A1(n_10031),
.A2(n_8656),
.B(n_8630),
.Y(n_10813)
);

OR2x2_ASAP7_75t_L g10814 ( 
.A(n_10073),
.B(n_8396),
.Y(n_10814)
);

AOI21x1_ASAP7_75t_L g10815 ( 
.A1(n_9846),
.A2(n_8200),
.B(n_8082),
.Y(n_10815)
);

NOR2xp33_ASAP7_75t_L g10816 ( 
.A(n_9970),
.B(n_7837),
.Y(n_10816)
);

CKINVDCx5p33_ASAP7_75t_R g10817 ( 
.A(n_9794),
.Y(n_10817)
);

INVx1_ASAP7_75t_L g10818 ( 
.A(n_9853),
.Y(n_10818)
);

INVx1_ASAP7_75t_L g10819 ( 
.A(n_9853),
.Y(n_10819)
);

AOI21x1_ASAP7_75t_L g10820 ( 
.A1(n_9853),
.A2(n_8200),
.B(n_8884),
.Y(n_10820)
);

BUFx6f_ASAP7_75t_L g10821 ( 
.A(n_9060),
.Y(n_10821)
);

OAI21x1_ASAP7_75t_L g10822 ( 
.A1(n_10145),
.A2(n_8580),
.B(n_7746),
.Y(n_10822)
);

OAI21x1_ASAP7_75t_L g10823 ( 
.A1(n_10145),
.A2(n_7746),
.B(n_7721),
.Y(n_10823)
);

OAI21x1_ASAP7_75t_L g10824 ( 
.A1(n_10145),
.A2(n_7746),
.B(n_7721),
.Y(n_10824)
);

HB1xp67_ASAP7_75t_L g10825 ( 
.A(n_9200),
.Y(n_10825)
);

AOI21x1_ASAP7_75t_L g10826 ( 
.A1(n_9853),
.A2(n_8200),
.B(n_8884),
.Y(n_10826)
);

AOI22xp5_ASAP7_75t_L g10827 ( 
.A1(n_10071),
.A2(n_8339),
.B1(n_8413),
.B2(n_8403),
.Y(n_10827)
);

AOI22xp33_ASAP7_75t_SL g10828 ( 
.A1(n_10068),
.A2(n_8407),
.B1(n_8501),
.B2(n_7685),
.Y(n_10828)
);

AND2x4_ASAP7_75t_L g10829 ( 
.A(n_9666),
.B(n_8279),
.Y(n_10829)
);

OAI21x1_ASAP7_75t_L g10830 ( 
.A1(n_10145),
.A2(n_7746),
.B(n_7721),
.Y(n_10830)
);

NAND2x1p5_ASAP7_75t_L g10831 ( 
.A(n_9229),
.B(n_8300),
.Y(n_10831)
);

NOR2x1_ASAP7_75t_SL g10832 ( 
.A(n_9272),
.B(n_7749),
.Y(n_10832)
);

AND2x4_ASAP7_75t_L g10833 ( 
.A(n_9666),
.B(n_8279),
.Y(n_10833)
);

BUFx6f_ASAP7_75t_L g10834 ( 
.A(n_9060),
.Y(n_10834)
);

AO21x2_ASAP7_75t_L g10835 ( 
.A1(n_9978),
.A2(n_8609),
.B(n_8387),
.Y(n_10835)
);

INVx1_ASAP7_75t_L g10836 ( 
.A(n_9877),
.Y(n_10836)
);

INVx1_ASAP7_75t_L g10837 ( 
.A(n_9877),
.Y(n_10837)
);

AND2x4_ASAP7_75t_L g10838 ( 
.A(n_9666),
.B(n_8279),
.Y(n_10838)
);

OAI21x1_ASAP7_75t_L g10839 ( 
.A1(n_10145),
.A2(n_7721),
.B(n_8656),
.Y(n_10839)
);

INVx1_ASAP7_75t_L g10840 ( 
.A(n_9877),
.Y(n_10840)
);

NAND2xp5_ASAP7_75t_L g10841 ( 
.A(n_10165),
.B(n_8001),
.Y(n_10841)
);

OAI21x1_ASAP7_75t_L g10842 ( 
.A1(n_10147),
.A2(n_8958),
.B(n_8797),
.Y(n_10842)
);

INVx2_ASAP7_75t_L g10843 ( 
.A(n_9337),
.Y(n_10843)
);

AOI21xp5_ASAP7_75t_L g10844 ( 
.A1(n_10138),
.A2(n_7737),
.B(n_7730),
.Y(n_10844)
);

NAND2xp5_ASAP7_75t_L g10845 ( 
.A(n_10165),
.B(n_8184),
.Y(n_10845)
);

NAND2x1p5_ASAP7_75t_L g10846 ( 
.A(n_9229),
.B(n_8300),
.Y(n_10846)
);

BUFx3_ASAP7_75t_L g10847 ( 
.A(n_9131),
.Y(n_10847)
);

INVx2_ASAP7_75t_L g10848 ( 
.A(n_9337),
.Y(n_10848)
);

INVx1_ASAP7_75t_L g10849 ( 
.A(n_9877),
.Y(n_10849)
);

AOI21xp5_ASAP7_75t_L g10850 ( 
.A1(n_9960),
.A2(n_7730),
.B(n_8160),
.Y(n_10850)
);

NAND2xp5_ASAP7_75t_L g10851 ( 
.A(n_9432),
.B(n_8184),
.Y(n_10851)
);

OAI21x1_ASAP7_75t_L g10852 ( 
.A1(n_10147),
.A2(n_8958),
.B(n_8797),
.Y(n_10852)
);

INVx1_ASAP7_75t_L g10853 ( 
.A(n_9878),
.Y(n_10853)
);

BUFx3_ASAP7_75t_L g10854 ( 
.A(n_9131),
.Y(n_10854)
);

INVx1_ASAP7_75t_L g10855 ( 
.A(n_9878),
.Y(n_10855)
);

OAI21x1_ASAP7_75t_L g10856 ( 
.A1(n_10147),
.A2(n_8958),
.B(n_8797),
.Y(n_10856)
);

OA21x2_ASAP7_75t_L g10857 ( 
.A1(n_10073),
.A2(n_8698),
.B(n_8569),
.Y(n_10857)
);

OR2x2_ASAP7_75t_L g10858 ( 
.A(n_10073),
.B(n_8396),
.Y(n_10858)
);

INVx1_ASAP7_75t_L g10859 ( 
.A(n_9878),
.Y(n_10859)
);

INVx1_ASAP7_75t_L g10860 ( 
.A(n_9878),
.Y(n_10860)
);

INVx2_ASAP7_75t_L g10861 ( 
.A(n_9337),
.Y(n_10861)
);

INVx6_ASAP7_75t_L g10862 ( 
.A(n_9131),
.Y(n_10862)
);

OAI21x1_ASAP7_75t_L g10863 ( 
.A1(n_10147),
.A2(n_8958),
.B(n_8832),
.Y(n_10863)
);

HB1xp67_ASAP7_75t_L g10864 ( 
.A(n_9200),
.Y(n_10864)
);

OA21x2_ASAP7_75t_L g10865 ( 
.A1(n_10073),
.A2(n_8698),
.B(n_8569),
.Y(n_10865)
);

NAND2xp5_ASAP7_75t_SL g10866 ( 
.A(n_9255),
.B(n_8751),
.Y(n_10866)
);

INVx4_ASAP7_75t_L g10867 ( 
.A(n_9148),
.Y(n_10867)
);

OAI21x1_ASAP7_75t_L g10868 ( 
.A1(n_10147),
.A2(n_8832),
.B(n_8267),
.Y(n_10868)
);

NAND3xp33_ASAP7_75t_SL g10869 ( 
.A(n_9969),
.B(n_7699),
.C(n_8560),
.Y(n_10869)
);

AND2x4_ASAP7_75t_L g10870 ( 
.A(n_9666),
.B(n_8279),
.Y(n_10870)
);

OAI21x1_ASAP7_75t_L g10871 ( 
.A1(n_9685),
.A2(n_8832),
.B(n_8267),
.Y(n_10871)
);

OAI21x1_ASAP7_75t_L g10872 ( 
.A1(n_9685),
.A2(n_8267),
.B(n_7766),
.Y(n_10872)
);

OAI21x1_ASAP7_75t_L g10873 ( 
.A1(n_9685),
.A2(n_8267),
.B(n_7766),
.Y(n_10873)
);

OA21x2_ASAP7_75t_L g10874 ( 
.A1(n_9685),
.A2(n_8278),
.B(n_8276),
.Y(n_10874)
);

OAI21x1_ASAP7_75t_L g10875 ( 
.A1(n_9685),
.A2(n_7766),
.B(n_7760),
.Y(n_10875)
);

AOI21x1_ASAP7_75t_L g10876 ( 
.A1(n_9903),
.A2(n_8891),
.B(n_8884),
.Y(n_10876)
);

BUFx12f_ASAP7_75t_L g10877 ( 
.A(n_9489),
.Y(n_10877)
);

HB1xp67_ASAP7_75t_L g10878 ( 
.A(n_9330),
.Y(n_10878)
);

AO21x2_ASAP7_75t_L g10879 ( 
.A1(n_9978),
.A2(n_9986),
.B(n_9943),
.Y(n_10879)
);

INVx1_ASAP7_75t_L g10880 ( 
.A(n_9903),
.Y(n_10880)
);

INVx2_ASAP7_75t_L g10881 ( 
.A(n_9337),
.Y(n_10881)
);

OAI21x1_ASAP7_75t_L g10882 ( 
.A1(n_10122),
.A2(n_7766),
.B(n_7760),
.Y(n_10882)
);

INVx2_ASAP7_75t_L g10883 ( 
.A(n_9337),
.Y(n_10883)
);

CKINVDCx5p33_ASAP7_75t_R g10884 ( 
.A(n_9794),
.Y(n_10884)
);

NAND2xp5_ASAP7_75t_L g10885 ( 
.A(n_9432),
.B(n_8190),
.Y(n_10885)
);

NOR2xp33_ASAP7_75t_L g10886 ( 
.A(n_9950),
.B(n_9962),
.Y(n_10886)
);

OAI21xp5_ASAP7_75t_L g10887 ( 
.A1(n_9950),
.A2(n_8389),
.B(n_8522),
.Y(n_10887)
);

HB1xp67_ASAP7_75t_L g10888 ( 
.A(n_9330),
.Y(n_10888)
);

INVx1_ASAP7_75t_L g10889 ( 
.A(n_9903),
.Y(n_10889)
);

OAI21x1_ASAP7_75t_SL g10890 ( 
.A1(n_10141),
.A2(n_8528),
.B(n_8712),
.Y(n_10890)
);

OAI21x1_ASAP7_75t_SL g10891 ( 
.A1(n_10141),
.A2(n_8528),
.B(n_8712),
.Y(n_10891)
);

NAND2x1p5_ASAP7_75t_L g10892 ( 
.A(n_9229),
.B(n_8300),
.Y(n_10892)
);

NAND2x1p5_ASAP7_75t_L g10893 ( 
.A(n_9229),
.B(n_8300),
.Y(n_10893)
);

OAI21xp5_ASAP7_75t_L g10894 ( 
.A1(n_10071),
.A2(n_10109),
.B(n_9788),
.Y(n_10894)
);

INVx1_ASAP7_75t_L g10895 ( 
.A(n_9903),
.Y(n_10895)
);

OA21x2_ASAP7_75t_L g10896 ( 
.A1(n_9627),
.A2(n_8278),
.B(n_8276),
.Y(n_10896)
);

AO21x2_ASAP7_75t_L g10897 ( 
.A1(n_9978),
.A2(n_8387),
.B(n_8340),
.Y(n_10897)
);

OR2x6_ASAP7_75t_L g10898 ( 
.A(n_9577),
.B(n_8369),
.Y(n_10898)
);

INVx3_ASAP7_75t_L g10899 ( 
.A(n_9666),
.Y(n_10899)
);

OAI21x1_ASAP7_75t_L g10900 ( 
.A1(n_10122),
.A2(n_7760),
.B(n_7759),
.Y(n_10900)
);

NAND3xp33_ASAP7_75t_L g10901 ( 
.A(n_9788),
.B(n_8560),
.C(n_8506),
.Y(n_10901)
);

NOR2xp67_ASAP7_75t_L g10902 ( 
.A(n_8995),
.B(n_7749),
.Y(n_10902)
);

INVx1_ASAP7_75t_L g10903 ( 
.A(n_9912),
.Y(n_10903)
);

AND2x2_ASAP7_75t_L g10904 ( 
.A(n_9403),
.B(n_7948),
.Y(n_10904)
);

INVx1_ASAP7_75t_L g10905 ( 
.A(n_9912),
.Y(n_10905)
);

AO21x2_ASAP7_75t_L g10906 ( 
.A1(n_9978),
.A2(n_8340),
.B(n_8722),
.Y(n_10906)
);

BUFx8_ASAP7_75t_L g10907 ( 
.A(n_9161),
.Y(n_10907)
);

INVx3_ASAP7_75t_L g10908 ( 
.A(n_9666),
.Y(n_10908)
);

AOI21xp5_ASAP7_75t_L g10909 ( 
.A1(n_9960),
.A2(n_9788),
.B(n_10141),
.Y(n_10909)
);

INVx2_ASAP7_75t_L g10910 ( 
.A(n_9462),
.Y(n_10910)
);

BUFx2_ASAP7_75t_L g10911 ( 
.A(n_9672),
.Y(n_10911)
);

OAI21x1_ASAP7_75t_L g10912 ( 
.A1(n_10122),
.A2(n_7760),
.B(n_7759),
.Y(n_10912)
);

INVx1_ASAP7_75t_L g10913 ( 
.A(n_9912),
.Y(n_10913)
);

HB1xp67_ASAP7_75t_L g10914 ( 
.A(n_9330),
.Y(n_10914)
);

OAI21x1_ASAP7_75t_L g10915 ( 
.A1(n_10122),
.A2(n_7759),
.B(n_8114),
.Y(n_10915)
);

HB1xp67_ASAP7_75t_L g10916 ( 
.A(n_9556),
.Y(n_10916)
);

OA21x2_ASAP7_75t_L g10917 ( 
.A1(n_9627),
.A2(n_8715),
.B(n_8579),
.Y(n_10917)
);

AOI22xp5_ASAP7_75t_L g10918 ( 
.A1(n_9998),
.A2(n_10109),
.B1(n_10092),
.B2(n_10186),
.Y(n_10918)
);

BUFx2_ASAP7_75t_R g10919 ( 
.A(n_9219),
.Y(n_10919)
);

NAND2xp5_ASAP7_75t_L g10920 ( 
.A(n_9432),
.B(n_8190),
.Y(n_10920)
);

NAND2xp5_ASAP7_75t_L g10921 ( 
.A(n_9389),
.B(n_8199),
.Y(n_10921)
);

OAI21x1_ASAP7_75t_L g10922 ( 
.A1(n_10122),
.A2(n_7759),
.B(n_8114),
.Y(n_10922)
);

INVx2_ASAP7_75t_SL g10923 ( 
.A(n_9577),
.Y(n_10923)
);

OAI21x1_ASAP7_75t_L g10924 ( 
.A1(n_9398),
.A2(n_9434),
.B(n_9417),
.Y(n_10924)
);

OAI21xp5_ASAP7_75t_L g10925 ( 
.A1(n_10109),
.A2(n_8389),
.B(n_8522),
.Y(n_10925)
);

AND2x2_ASAP7_75t_L g10926 ( 
.A(n_9451),
.B(n_7948),
.Y(n_10926)
);

OA21x2_ASAP7_75t_L g10927 ( 
.A1(n_9627),
.A2(n_8715),
.B(n_8579),
.Y(n_10927)
);

AND2x2_ASAP7_75t_L g10928 ( 
.A(n_9451),
.B(n_7949),
.Y(n_10928)
);

AND2x2_ASAP7_75t_L g10929 ( 
.A(n_9451),
.B(n_7949),
.Y(n_10929)
);

INVx1_ASAP7_75t_L g10930 ( 
.A(n_9912),
.Y(n_10930)
);

AOI21x1_ASAP7_75t_L g10931 ( 
.A1(n_9917),
.A2(n_8932),
.B(n_8891),
.Y(n_10931)
);

INVx1_ASAP7_75t_L g10932 ( 
.A(n_9917),
.Y(n_10932)
);

OAI21x1_ASAP7_75t_L g10933 ( 
.A1(n_9398),
.A2(n_8114),
.B(n_8389),
.Y(n_10933)
);

INVx1_ASAP7_75t_SL g10934 ( 
.A(n_9428),
.Y(n_10934)
);

INVx1_ASAP7_75t_L g10935 ( 
.A(n_9917),
.Y(n_10935)
);

INVx2_ASAP7_75t_L g10936 ( 
.A(n_9462),
.Y(n_10936)
);

INVx1_ASAP7_75t_L g10937 ( 
.A(n_9917),
.Y(n_10937)
);

INVx1_ASAP7_75t_L g10938 ( 
.A(n_9935),
.Y(n_10938)
);

NOR2xp67_ASAP7_75t_L g10939 ( 
.A(n_9816),
.B(n_9254),
.Y(n_10939)
);

OAI21xp5_ASAP7_75t_L g10940 ( 
.A1(n_10109),
.A2(n_8339),
.B(n_8506),
.Y(n_10940)
);

INVx1_ASAP7_75t_L g10941 ( 
.A(n_9935),
.Y(n_10941)
);

AO21x2_ASAP7_75t_L g10942 ( 
.A1(n_9978),
.A2(n_8340),
.B(n_8722),
.Y(n_10942)
);

NAND2xp5_ASAP7_75t_L g10943 ( 
.A(n_9389),
.B(n_8199),
.Y(n_10943)
);

OAI21x1_ASAP7_75t_L g10944 ( 
.A1(n_9398),
.A2(n_8114),
.B(n_8398),
.Y(n_10944)
);

AOI21xp5_ASAP7_75t_L g10945 ( 
.A1(n_9960),
.A2(n_8160),
.B(n_8538),
.Y(n_10945)
);

OAI21x1_ASAP7_75t_L g10946 ( 
.A1(n_9398),
.A2(n_8410),
.B(n_8398),
.Y(n_10946)
);

INVx2_ASAP7_75t_L g10947 ( 
.A(n_9462),
.Y(n_10947)
);

CKINVDCx20_ASAP7_75t_R g10948 ( 
.A(n_9225),
.Y(n_10948)
);

NAND2xp5_ASAP7_75t_L g10949 ( 
.A(n_9389),
.B(n_8308),
.Y(n_10949)
);

NAND2xp5_ASAP7_75t_L g10950 ( 
.A(n_9395),
.B(n_8308),
.Y(n_10950)
);

OAI21x1_ASAP7_75t_L g10951 ( 
.A1(n_9398),
.A2(n_8410),
.B(n_8398),
.Y(n_10951)
);

NOR2xp33_ASAP7_75t_L g10952 ( 
.A(n_9962),
.B(n_10186),
.Y(n_10952)
);

OAI21x1_ASAP7_75t_L g10953 ( 
.A1(n_9417),
.A2(n_9434),
.B(n_9973),
.Y(n_10953)
);

OAI21x1_ASAP7_75t_SL g10954 ( 
.A1(n_9407),
.A2(n_7904),
.B(n_7792),
.Y(n_10954)
);

INVx2_ASAP7_75t_L g10955 ( 
.A(n_9337),
.Y(n_10955)
);

INVx1_ASAP7_75t_L g10956 ( 
.A(n_9935),
.Y(n_10956)
);

OAI21x1_ASAP7_75t_L g10957 ( 
.A1(n_9417),
.A2(n_9434),
.B(n_9973),
.Y(n_10957)
);

INVx1_ASAP7_75t_L g10958 ( 
.A(n_9935),
.Y(n_10958)
);

A2O1A1Ixp33_ASAP7_75t_L g10959 ( 
.A1(n_10068),
.A2(n_8538),
.B(n_7701),
.C(n_8329),
.Y(n_10959)
);

INVx3_ASAP7_75t_L g10960 ( 
.A(n_9672),
.Y(n_10960)
);

INVx2_ASAP7_75t_L g10961 ( 
.A(n_9337),
.Y(n_10961)
);

OAI21xp5_ASAP7_75t_L g10962 ( 
.A1(n_10060),
.A2(n_8770),
.B(n_8309),
.Y(n_10962)
);

OA21x2_ASAP7_75t_L g10963 ( 
.A1(n_9627),
.A2(n_8547),
.B(n_8786),
.Y(n_10963)
);

OAI21x1_ASAP7_75t_L g10964 ( 
.A1(n_9417),
.A2(n_8410),
.B(n_8398),
.Y(n_10964)
);

INVx1_ASAP7_75t_L g10965 ( 
.A(n_9508),
.Y(n_10965)
);

OA21x2_ASAP7_75t_L g10966 ( 
.A1(n_9627),
.A2(n_8547),
.B(n_8786),
.Y(n_10966)
);

OAI21x1_ASAP7_75t_L g10967 ( 
.A1(n_9417),
.A2(n_8410),
.B(n_8398),
.Y(n_10967)
);

OAI21x1_ASAP7_75t_L g10968 ( 
.A1(n_9434),
.A2(n_8410),
.B(n_8398),
.Y(n_10968)
);

OAI21x1_ASAP7_75t_L g10969 ( 
.A1(n_9434),
.A2(n_8415),
.B(n_8410),
.Y(n_10969)
);

INVx4_ASAP7_75t_L g10970 ( 
.A(n_9161),
.Y(n_10970)
);

INVx2_ASAP7_75t_SL g10971 ( 
.A(n_9577),
.Y(n_10971)
);

NAND2x1p5_ASAP7_75t_L g10972 ( 
.A(n_9229),
.B(n_8300),
.Y(n_10972)
);

OAI21x1_ASAP7_75t_L g10973 ( 
.A1(n_9973),
.A2(n_9985),
.B(n_9373),
.Y(n_10973)
);

INVx1_ASAP7_75t_L g10974 ( 
.A(n_9508),
.Y(n_10974)
);

INVx1_ASAP7_75t_L g10975 ( 
.A(n_9508),
.Y(n_10975)
);

INVx2_ASAP7_75t_L g10976 ( 
.A(n_9337),
.Y(n_10976)
);

NAND2xp5_ASAP7_75t_L g10977 ( 
.A(n_9395),
.B(n_8317),
.Y(n_10977)
);

NAND2xp5_ASAP7_75t_L g10978 ( 
.A(n_9395),
.B(n_8317),
.Y(n_10978)
);

OA21x2_ASAP7_75t_L g10979 ( 
.A1(n_9695),
.A2(n_8907),
.B(n_8906),
.Y(n_10979)
);

AO31x2_ASAP7_75t_L g10980 ( 
.A1(n_9552),
.A2(n_9579),
.A3(n_9414),
.B(n_9879),
.Y(n_10980)
);

NAND3xp33_ASAP7_75t_L g10981 ( 
.A(n_10151),
.B(n_10058),
.C(n_10060),
.Y(n_10981)
);

INVx2_ASAP7_75t_L g10982 ( 
.A(n_9462),
.Y(n_10982)
);

AOI22xp5_ASAP7_75t_L g10983 ( 
.A1(n_9998),
.A2(n_10092),
.B1(n_10186),
.B2(n_10005),
.Y(n_10983)
);

OAI21x1_ASAP7_75t_L g10984 ( 
.A1(n_9973),
.A2(n_8461),
.B(n_8415),
.Y(n_10984)
);

AO31x2_ASAP7_75t_L g10985 ( 
.A1(n_9552),
.A2(n_8527),
.A3(n_8364),
.B(n_8240),
.Y(n_10985)
);

BUFx8_ASAP7_75t_L g10986 ( 
.A(n_9161),
.Y(n_10986)
);

INVx1_ASAP7_75t_L g10987 ( 
.A(n_9508),
.Y(n_10987)
);

INVx1_ASAP7_75t_L g10988 ( 
.A(n_9508),
.Y(n_10988)
);

OA21x2_ASAP7_75t_L g10989 ( 
.A1(n_9695),
.A2(n_8907),
.B(n_8906),
.Y(n_10989)
);

OAI21x1_ASAP7_75t_L g10990 ( 
.A1(n_9973),
.A2(n_8461),
.B(n_8415),
.Y(n_10990)
);

OA21x2_ASAP7_75t_L g10991 ( 
.A1(n_9695),
.A2(n_9703),
.B(n_9696),
.Y(n_10991)
);

BUFx3_ASAP7_75t_L g10992 ( 
.A(n_9131),
.Y(n_10992)
);

INVx2_ASAP7_75t_L g10993 ( 
.A(n_9462),
.Y(n_10993)
);

NAND2xp5_ASAP7_75t_L g10994 ( 
.A(n_9408),
.B(n_9111),
.Y(n_10994)
);

INVx2_ASAP7_75t_L g10995 ( 
.A(n_9462),
.Y(n_10995)
);

OAI21xp5_ASAP7_75t_L g10996 ( 
.A1(n_10060),
.A2(n_8309),
.B(n_8294),
.Y(n_10996)
);

INVx1_ASAP7_75t_L g10997 ( 
.A(n_9667),
.Y(n_10997)
);

OA21x2_ASAP7_75t_L g10998 ( 
.A1(n_9695),
.A2(n_8917),
.B(n_8908),
.Y(n_10998)
);

OAI21x1_ASAP7_75t_SL g10999 ( 
.A1(n_9407),
.A2(n_7904),
.B(n_7792),
.Y(n_10999)
);

NAND2xp5_ASAP7_75t_SL g11000 ( 
.A(n_9255),
.B(n_8475),
.Y(n_11000)
);

NAND2xp5_ASAP7_75t_L g11001 ( 
.A(n_9408),
.B(n_8872),
.Y(n_11001)
);

BUFx6f_ASAP7_75t_L g11002 ( 
.A(n_9060),
.Y(n_11002)
);

OAI21x1_ASAP7_75t_L g11003 ( 
.A1(n_9985),
.A2(n_9373),
.B(n_9886),
.Y(n_11003)
);

AOI22xp5_ASAP7_75t_L g11004 ( 
.A1(n_9998),
.A2(n_8403),
.B1(n_8413),
.B2(n_8437),
.Y(n_11004)
);

AO21x2_ASAP7_75t_L g11005 ( 
.A1(n_9978),
.A2(n_8413),
.B(n_8403),
.Y(n_11005)
);

OAI21x1_ASAP7_75t_SL g11006 ( 
.A1(n_9407),
.A2(n_7904),
.B(n_7792),
.Y(n_11006)
);

AO21x2_ASAP7_75t_L g11007 ( 
.A1(n_9978),
.A2(n_8931),
.B(n_8911),
.Y(n_11007)
);

HB1xp67_ASAP7_75t_L g11008 ( 
.A(n_9556),
.Y(n_11008)
);

AND2x4_ASAP7_75t_L g11009 ( 
.A(n_9672),
.B(n_8279),
.Y(n_11009)
);

NAND2xp5_ASAP7_75t_SL g11010 ( 
.A(n_9255),
.B(n_8475),
.Y(n_11010)
);

NAND2xp5_ASAP7_75t_L g11011 ( 
.A(n_9408),
.B(n_8872),
.Y(n_11011)
);

INVx5_ASAP7_75t_L g11012 ( 
.A(n_10148),
.Y(n_11012)
);

AO31x2_ASAP7_75t_L g11013 ( 
.A1(n_9414),
.A2(n_8240),
.A3(n_8229),
.B(n_8615),
.Y(n_11013)
);

A2O1A1Ixp33_ASAP7_75t_L g11014 ( 
.A1(n_10186),
.A2(n_7701),
.B(n_8329),
.C(n_8473),
.Y(n_11014)
);

INVx2_ASAP7_75t_L g11015 ( 
.A(n_9462),
.Y(n_11015)
);

AND2x4_ASAP7_75t_L g11016 ( 
.A(n_9672),
.B(n_9686),
.Y(n_11016)
);

NAND2xp5_ASAP7_75t_L g11017 ( 
.A(n_9111),
.B(n_8872),
.Y(n_11017)
);

INVx1_ASAP7_75t_L g11018 ( 
.A(n_9667),
.Y(n_11018)
);

INVx2_ASAP7_75t_L g11019 ( 
.A(n_9478),
.Y(n_11019)
);

INVx1_ASAP7_75t_L g11020 ( 
.A(n_9667),
.Y(n_11020)
);

AND2x2_ASAP7_75t_L g11021 ( 
.A(n_9487),
.B(n_7949),
.Y(n_11021)
);

AO31x2_ASAP7_75t_L g11022 ( 
.A1(n_9414),
.A2(n_8240),
.A3(n_8229),
.B(n_8615),
.Y(n_11022)
);

OAI21x1_ASAP7_75t_L g11023 ( 
.A1(n_9985),
.A2(n_8461),
.B(n_8415),
.Y(n_11023)
);

INVx2_ASAP7_75t_L g11024 ( 
.A(n_9478),
.Y(n_11024)
);

INVx1_ASAP7_75t_L g11025 ( 
.A(n_9667),
.Y(n_11025)
);

AO31x2_ASAP7_75t_L g11026 ( 
.A1(n_9579),
.A2(n_8240),
.A3(n_8229),
.B(n_8615),
.Y(n_11026)
);

INVx1_ASAP7_75t_L g11027 ( 
.A(n_9667),
.Y(n_11027)
);

NAND2x1p5_ASAP7_75t_L g11028 ( 
.A(n_9229),
.B(n_8420),
.Y(n_11028)
);

INVx2_ASAP7_75t_L g11029 ( 
.A(n_9478),
.Y(n_11029)
);

OAI21x1_ASAP7_75t_L g11030 ( 
.A1(n_9985),
.A2(n_8461),
.B(n_8415),
.Y(n_11030)
);

OAI21xp5_ASAP7_75t_L g11031 ( 
.A1(n_10099),
.A2(n_8350),
.B(n_8294),
.Y(n_11031)
);

INVx1_ASAP7_75t_L g11032 ( 
.A(n_9894),
.Y(n_11032)
);

OR2x2_ASAP7_75t_L g11033 ( 
.A(n_9190),
.B(n_8396),
.Y(n_11033)
);

AO31x2_ASAP7_75t_L g11034 ( 
.A1(n_9579),
.A2(n_8229),
.A3(n_8615),
.B(n_8649),
.Y(n_11034)
);

INVx1_ASAP7_75t_L g11035 ( 
.A(n_9894),
.Y(n_11035)
);

INVx1_ASAP7_75t_L g11036 ( 
.A(n_9894),
.Y(n_11036)
);

AO21x1_ASAP7_75t_L g11037 ( 
.A1(n_10092),
.A2(n_8511),
.B(n_8911),
.Y(n_11037)
);

NOR2x1_ASAP7_75t_R g11038 ( 
.A(n_9489),
.B(n_8338),
.Y(n_11038)
);

OAI21x1_ASAP7_75t_L g11039 ( 
.A1(n_9985),
.A2(n_8461),
.B(n_8415),
.Y(n_11039)
);

OAI21x1_ASAP7_75t_L g11040 ( 
.A1(n_9373),
.A2(n_8461),
.B(n_7754),
.Y(n_11040)
);

OAI21x1_ASAP7_75t_SL g11041 ( 
.A1(n_9407),
.A2(n_7904),
.B(n_7792),
.Y(n_11041)
);

OAI21x1_ASAP7_75t_L g11042 ( 
.A1(n_9373),
.A2(n_7754),
.B(n_7695),
.Y(n_11042)
);

INVx3_ASAP7_75t_L g11043 ( 
.A(n_9672),
.Y(n_11043)
);

NAND2xp5_ASAP7_75t_L g11044 ( 
.A(n_9111),
.B(n_8441),
.Y(n_11044)
);

AOI21xp5_ASAP7_75t_SL g11045 ( 
.A1(n_10146),
.A2(n_8298),
.B(n_8466),
.Y(n_11045)
);

AOI21xp5_ASAP7_75t_L g11046 ( 
.A1(n_9960),
.A2(n_8371),
.B(n_8365),
.Y(n_11046)
);

AOI21x1_ASAP7_75t_L g11047 ( 
.A1(n_9939),
.A2(n_8932),
.B(n_8891),
.Y(n_11047)
);

OA21x2_ASAP7_75t_L g11048 ( 
.A1(n_9695),
.A2(n_8917),
.B(n_8908),
.Y(n_11048)
);

NAND2xp5_ASAP7_75t_SL g11049 ( 
.A(n_9255),
.B(n_8475),
.Y(n_11049)
);

INVx1_ASAP7_75t_L g11050 ( 
.A(n_9894),
.Y(n_11050)
);

AOI21xp5_ASAP7_75t_L g11051 ( 
.A1(n_10099),
.A2(n_8371),
.B(n_8365),
.Y(n_11051)
);

NAND3xp33_ASAP7_75t_L g11052 ( 
.A(n_10151),
.B(n_8931),
.C(n_8147),
.Y(n_11052)
);

OAI21x1_ASAP7_75t_L g11053 ( 
.A1(n_9373),
.A2(n_7754),
.B(n_7695),
.Y(n_11053)
);

OAI21x1_ASAP7_75t_L g11054 ( 
.A1(n_9886),
.A2(n_7754),
.B(n_7695),
.Y(n_11054)
);

HB1xp67_ASAP7_75t_L g11055 ( 
.A(n_9556),
.Y(n_11055)
);

OAI21x1_ASAP7_75t_L g11056 ( 
.A1(n_9886),
.A2(n_7754),
.B(n_7695),
.Y(n_11056)
);

AO21x2_ASAP7_75t_L g11057 ( 
.A1(n_9978),
.A2(n_8931),
.B(n_8147),
.Y(n_11057)
);

OAI21xp5_ASAP7_75t_L g11058 ( 
.A1(n_10099),
.A2(n_8368),
.B(n_8350),
.Y(n_11058)
);

NAND2xp5_ASAP7_75t_SL g11059 ( 
.A(n_9201),
.B(n_9392),
.Y(n_11059)
);

INVx2_ASAP7_75t_L g11060 ( 
.A(n_9478),
.Y(n_11060)
);

INVx1_ASAP7_75t_L g11061 ( 
.A(n_9894),
.Y(n_11061)
);

OA21x2_ASAP7_75t_L g11062 ( 
.A1(n_9696),
.A2(n_8926),
.B(n_8921),
.Y(n_11062)
);

INVx2_ASAP7_75t_L g11063 ( 
.A(n_9478),
.Y(n_11063)
);

INVx1_ASAP7_75t_L g11064 ( 
.A(n_9919),
.Y(n_11064)
);

HB1xp67_ASAP7_75t_L g11065 ( 
.A(n_8998),
.Y(n_11065)
);

OR2x2_ASAP7_75t_L g11066 ( 
.A(n_9190),
.B(n_8396),
.Y(n_11066)
);

CKINVDCx20_ASAP7_75t_R g11067 ( 
.A(n_9225),
.Y(n_11067)
);

INVx1_ASAP7_75t_L g11068 ( 
.A(n_9919),
.Y(n_11068)
);

AOI21x1_ASAP7_75t_L g11069 ( 
.A1(n_9939),
.A2(n_8951),
.B(n_8932),
.Y(n_11069)
);

AND2x2_ASAP7_75t_L g11070 ( 
.A(n_9487),
.B(n_7949),
.Y(n_11070)
);

INVx1_ASAP7_75t_SL g11071 ( 
.A(n_9428),
.Y(n_11071)
);

OAI21x1_ASAP7_75t_L g11072 ( 
.A1(n_9471),
.A2(n_7870),
.B(n_7862),
.Y(n_11072)
);

BUFx2_ASAP7_75t_R g11073 ( 
.A(n_9219),
.Y(n_11073)
);

AND2x4_ASAP7_75t_L g11074 ( 
.A(n_9672),
.B(n_9686),
.Y(n_11074)
);

OAI21xp5_ASAP7_75t_L g11075 ( 
.A1(n_10005),
.A2(n_10025),
.B(n_10153),
.Y(n_11075)
);

INVx2_ASAP7_75t_L g11076 ( 
.A(n_9478),
.Y(n_11076)
);

BUFx3_ASAP7_75t_L g11077 ( 
.A(n_9131),
.Y(n_11077)
);

INVx1_ASAP7_75t_L g11078 ( 
.A(n_9919),
.Y(n_11078)
);

AOI21xp5_ASAP7_75t_L g11079 ( 
.A1(n_9625),
.A2(n_7740),
.B(n_7748),
.Y(n_11079)
);

HB1xp67_ASAP7_75t_L g11080 ( 
.A(n_8998),
.Y(n_11080)
);

NAND2xp5_ASAP7_75t_SL g11081 ( 
.A(n_9201),
.B(n_8475),
.Y(n_11081)
);

AO31x2_ASAP7_75t_L g11082 ( 
.A1(n_9552),
.A2(n_8649),
.A3(n_8961),
.B(n_8058),
.Y(n_11082)
);

INVx6_ASAP7_75t_L g11083 ( 
.A(n_9131),
.Y(n_11083)
);

OA21x2_ASAP7_75t_L g11084 ( 
.A1(n_9696),
.A2(n_8926),
.B(n_8921),
.Y(n_11084)
);

AO31x2_ASAP7_75t_L g11085 ( 
.A1(n_9552),
.A2(n_8649),
.A3(n_8961),
.B(n_8058),
.Y(n_11085)
);

INVx1_ASAP7_75t_L g11086 ( 
.A(n_9919),
.Y(n_11086)
);

AOI21x1_ASAP7_75t_L g11087 ( 
.A1(n_9939),
.A2(n_8951),
.B(n_8902),
.Y(n_11087)
);

NOR2xp33_ASAP7_75t_L g11088 ( 
.A(n_9050),
.B(n_7837),
.Y(n_11088)
);

OA21x2_ASAP7_75t_L g11089 ( 
.A1(n_9696),
.A2(n_8927),
.B(n_8936),
.Y(n_11089)
);

INVx2_ASAP7_75t_L g11090 ( 
.A(n_9478),
.Y(n_11090)
);

OAI21xp5_ASAP7_75t_L g11091 ( 
.A1(n_10005),
.A2(n_8368),
.B(n_8407),
.Y(n_11091)
);

INVx2_ASAP7_75t_L g11092 ( 
.A(n_9478),
.Y(n_11092)
);

AOI21xp5_ASAP7_75t_L g11093 ( 
.A1(n_9625),
.A2(n_7740),
.B(n_7748),
.Y(n_11093)
);

OA21x2_ASAP7_75t_L g11094 ( 
.A1(n_9696),
.A2(n_8927),
.B(n_8936),
.Y(n_11094)
);

OAI21x1_ASAP7_75t_L g11095 ( 
.A1(n_9674),
.A2(n_7876),
.B(n_7870),
.Y(n_11095)
);

INVx1_ASAP7_75t_L g11096 ( 
.A(n_9919),
.Y(n_11096)
);

NAND2xp5_ASAP7_75t_L g11097 ( 
.A(n_9168),
.B(n_8441),
.Y(n_11097)
);

INVx1_ASAP7_75t_L g11098 ( 
.A(n_9996),
.Y(n_11098)
);

BUFx2_ASAP7_75t_L g11099 ( 
.A(n_9686),
.Y(n_11099)
);

NOR2xp67_ASAP7_75t_SL g11100 ( 
.A(n_9161),
.B(n_7792),
.Y(n_11100)
);

INVx2_ASAP7_75t_L g11101 ( 
.A(n_9478),
.Y(n_11101)
);

NAND2xp5_ASAP7_75t_L g11102 ( 
.A(n_9168),
.B(n_8467),
.Y(n_11102)
);

INVx1_ASAP7_75t_L g11103 ( 
.A(n_9996),
.Y(n_11103)
);

INVx1_ASAP7_75t_L g11104 ( 
.A(n_9996),
.Y(n_11104)
);

INVx2_ASAP7_75t_L g11105 ( 
.A(n_9484),
.Y(n_11105)
);

INVx1_ASAP7_75t_L g11106 ( 
.A(n_9996),
.Y(n_11106)
);

AO31x2_ASAP7_75t_L g11107 ( 
.A1(n_9579),
.A2(n_8649),
.A3(n_8058),
.B(n_8537),
.Y(n_11107)
);

OA21x2_ASAP7_75t_L g11108 ( 
.A1(n_9703),
.A2(n_8940),
.B(n_8937),
.Y(n_11108)
);

INVx1_ASAP7_75t_L g11109 ( 
.A(n_9996),
.Y(n_11109)
);

INVx1_ASAP7_75t_L g11110 ( 
.A(n_10052),
.Y(n_11110)
);

INVx1_ASAP7_75t_L g11111 ( 
.A(n_10052),
.Y(n_11111)
);

AOI21xp5_ASAP7_75t_L g11112 ( 
.A1(n_9625),
.A2(n_8486),
.B(n_8407),
.Y(n_11112)
);

AND2x2_ASAP7_75t_L g11113 ( 
.A(n_9487),
.B(n_7749),
.Y(n_11113)
);

OA21x2_ASAP7_75t_L g11114 ( 
.A1(n_9703),
.A2(n_8940),
.B(n_8937),
.Y(n_11114)
);

OAI21x1_ASAP7_75t_SL g11115 ( 
.A1(n_8994),
.A2(n_7904),
.B(n_7761),
.Y(n_11115)
);

AND2x2_ASAP7_75t_L g11116 ( 
.A(n_9487),
.B(n_7749),
.Y(n_11116)
);

INVx1_ASAP7_75t_L g11117 ( 
.A(n_10052),
.Y(n_11117)
);

AO21x2_ASAP7_75t_L g11118 ( 
.A1(n_9986),
.A2(n_8437),
.B(n_8776),
.Y(n_11118)
);

INVx2_ASAP7_75t_L g11119 ( 
.A(n_9484),
.Y(n_11119)
);

AOI21xp5_ASAP7_75t_L g11120 ( 
.A1(n_9625),
.A2(n_8486),
.B(n_8407),
.Y(n_11120)
);

OAI21xp5_ASAP7_75t_L g11121 ( 
.A1(n_10025),
.A2(n_8407),
.B(n_8473),
.Y(n_11121)
);

OAI21x1_ASAP7_75t_L g11122 ( 
.A1(n_10183),
.A2(n_7884),
.B(n_7876),
.Y(n_11122)
);

CKINVDCx11_ASAP7_75t_R g11123 ( 
.A(n_9161),
.Y(n_11123)
);

INVx2_ASAP7_75t_L g11124 ( 
.A(n_9484),
.Y(n_11124)
);

INVx2_ASAP7_75t_L g11125 ( 
.A(n_9484),
.Y(n_11125)
);

NAND2xp5_ASAP7_75t_L g11126 ( 
.A(n_9168),
.B(n_8467),
.Y(n_11126)
);

OAI21x1_ASAP7_75t_L g11127 ( 
.A1(n_10183),
.A2(n_7895),
.B(n_7884),
.Y(n_11127)
);

INVx2_ASAP7_75t_L g11128 ( 
.A(n_9484),
.Y(n_11128)
);

OAI21x1_ASAP7_75t_L g11129 ( 
.A1(n_10183),
.A2(n_7903),
.B(n_7895),
.Y(n_11129)
);

AO22x2_ASAP7_75t_L g11130 ( 
.A1(n_9816),
.A2(n_7842),
.B1(n_7864),
.B2(n_7761),
.Y(n_11130)
);

OAI21xp5_ASAP7_75t_L g11131 ( 
.A1(n_10025),
.A2(n_8473),
.B(n_7699),
.Y(n_11131)
);

INVx1_ASAP7_75t_L g11132 ( 
.A(n_10052),
.Y(n_11132)
);

INVx2_ASAP7_75t_L g11133 ( 
.A(n_9484),
.Y(n_11133)
);

INVx2_ASAP7_75t_L g11134 ( 
.A(n_9484),
.Y(n_11134)
);

INVx4_ASAP7_75t_L g11135 ( 
.A(n_9161),
.Y(n_11135)
);

NAND2xp5_ASAP7_75t_L g11136 ( 
.A(n_9691),
.B(n_8781),
.Y(n_11136)
);

AO21x2_ASAP7_75t_L g11137 ( 
.A1(n_9986),
.A2(n_8437),
.B(n_8776),
.Y(n_11137)
);

NOR2xp33_ASAP7_75t_L g11138 ( 
.A(n_9050),
.B(n_8182),
.Y(n_11138)
);

OAI21x1_ASAP7_75t_L g11139 ( 
.A1(n_10185),
.A2(n_7903),
.B(n_7895),
.Y(n_11139)
);

OAI21x1_ASAP7_75t_L g11140 ( 
.A1(n_10185),
.A2(n_7903),
.B(n_7895),
.Y(n_11140)
);

AOI21xp5_ASAP7_75t_L g11141 ( 
.A1(n_9732),
.A2(n_7733),
.B(n_7719),
.Y(n_11141)
);

INVx1_ASAP7_75t_L g11142 ( 
.A(n_10052),
.Y(n_11142)
);

OAI21xp5_ASAP7_75t_L g11143 ( 
.A1(n_10153),
.A2(n_7699),
.B(n_8501),
.Y(n_11143)
);

BUFx8_ASAP7_75t_L g11144 ( 
.A(n_9185),
.Y(n_11144)
);

OAI21x1_ASAP7_75t_L g11145 ( 
.A1(n_10185),
.A2(n_7903),
.B(n_7895),
.Y(n_11145)
);

OA21x2_ASAP7_75t_L g11146 ( 
.A1(n_9703),
.A2(n_8953),
.B(n_8952),
.Y(n_11146)
);

INVx2_ASAP7_75t_L g11147 ( 
.A(n_9484),
.Y(n_11147)
);

AO31x2_ASAP7_75t_L g11148 ( 
.A1(n_9552),
.A2(n_8058),
.A3(n_8537),
.B(n_8480),
.Y(n_11148)
);

INVx2_ASAP7_75t_L g11149 ( 
.A(n_9484),
.Y(n_11149)
);

OAI21x1_ASAP7_75t_L g11150 ( 
.A1(n_9893),
.A2(n_7903),
.B(n_7895),
.Y(n_11150)
);

AND2x2_ASAP7_75t_L g11151 ( 
.A(n_9519),
.B(n_7761),
.Y(n_11151)
);

AOI21xp5_ASAP7_75t_SL g11152 ( 
.A1(n_10146),
.A2(n_8298),
.B(n_8471),
.Y(n_11152)
);

AND2x2_ASAP7_75t_L g11153 ( 
.A(n_9519),
.B(n_7761),
.Y(n_11153)
);

OAI21xp5_ASAP7_75t_L g11154 ( 
.A1(n_10153),
.A2(n_8501),
.B(n_7733),
.Y(n_11154)
);

INVx2_ASAP7_75t_L g11155 ( 
.A(n_9449),
.Y(n_11155)
);

INVx2_ASAP7_75t_L g11156 ( 
.A(n_9449),
.Y(n_11156)
);

AO21x2_ASAP7_75t_L g11157 ( 
.A1(n_9986),
.A2(n_8776),
.B(n_8606),
.Y(n_11157)
);

INVx1_ASAP7_75t_L g11158 ( 
.A(n_9028),
.Y(n_11158)
);

OAI21x1_ASAP7_75t_SL g11159 ( 
.A1(n_8994),
.A2(n_7904),
.B(n_7864),
.Y(n_11159)
);

OA21x2_ASAP7_75t_L g11160 ( 
.A1(n_9703),
.A2(n_8953),
.B(n_8952),
.Y(n_11160)
);

INVxp67_ASAP7_75t_SL g11161 ( 
.A(n_9579),
.Y(n_11161)
);

INVx1_ASAP7_75t_L g11162 ( 
.A(n_9028),
.Y(n_11162)
);

INVx3_ASAP7_75t_L g11163 ( 
.A(n_9686),
.Y(n_11163)
);

OAI21x1_ASAP7_75t_SL g11164 ( 
.A1(n_8994),
.A2(n_7864),
.B(n_7842),
.Y(n_11164)
);

OA21x2_ASAP7_75t_L g11165 ( 
.A1(n_9690),
.A2(n_8969),
.B(n_8960),
.Y(n_11165)
);

AO21x1_ASAP7_75t_L g11166 ( 
.A1(n_9879),
.A2(n_8512),
.B(n_7834),
.Y(n_11166)
);

INVx1_ASAP7_75t_L g11167 ( 
.A(n_9028),
.Y(n_11167)
);

INVx1_ASAP7_75t_L g11168 ( 
.A(n_9144),
.Y(n_11168)
);

AO21x2_ASAP7_75t_L g11169 ( 
.A1(n_9986),
.A2(n_8606),
.B(n_8946),
.Y(n_11169)
);

A2O1A1Ixp33_ASAP7_75t_L g11170 ( 
.A1(n_10151),
.A2(n_7751),
.B(n_7685),
.C(n_8626),
.Y(n_11170)
);

OAI21x1_ASAP7_75t_L g11171 ( 
.A1(n_10176),
.A2(n_8096),
.B(n_8009),
.Y(n_11171)
);

AO21x2_ASAP7_75t_L g11172 ( 
.A1(n_9986),
.A2(n_8606),
.B(n_8946),
.Y(n_11172)
);

INVx1_ASAP7_75t_L g11173 ( 
.A(n_9144),
.Y(n_11173)
);

AOI21xp5_ASAP7_75t_L g11174 ( 
.A1(n_9732),
.A2(n_7719),
.B(n_7736),
.Y(n_11174)
);

INVx3_ASAP7_75t_SL g11175 ( 
.A(n_9025),
.Y(n_11175)
);

AO21x2_ASAP7_75t_L g11176 ( 
.A1(n_9986),
.A2(n_8790),
.B(n_8788),
.Y(n_11176)
);

AOI22xp33_ASAP7_75t_L g11177 ( 
.A1(n_10058),
.A2(n_8501),
.B1(n_8219),
.B2(n_8325),
.Y(n_11177)
);

NOR3xp33_ASAP7_75t_L g11178 ( 
.A(n_9887),
.B(n_8263),
.C(n_8239),
.Y(n_11178)
);

BUFx2_ASAP7_75t_L g11179 ( 
.A(n_9686),
.Y(n_11179)
);

OR2x6_ASAP7_75t_L g11180 ( 
.A(n_9577),
.B(n_7744),
.Y(n_11180)
);

AOI21xp5_ASAP7_75t_L g11181 ( 
.A1(n_9732),
.A2(n_7736),
.B(n_8501),
.Y(n_11181)
);

AND2x2_ASAP7_75t_L g11182 ( 
.A(n_9519),
.B(n_7842),
.Y(n_11182)
);

NAND2x1p5_ASAP7_75t_L g11183 ( 
.A(n_9229),
.B(n_8420),
.Y(n_11183)
);

AO21x2_ASAP7_75t_L g11184 ( 
.A1(n_9986),
.A2(n_8790),
.B(n_8788),
.Y(n_11184)
);

NAND2xp5_ASAP7_75t_L g11185 ( 
.A(n_9691),
.B(n_8781),
.Y(n_11185)
);

INVx1_ASAP7_75t_L g11186 ( 
.A(n_9144),
.Y(n_11186)
);

NAND2x1_ASAP7_75t_L g11187 ( 
.A(n_9952),
.B(n_7842),
.Y(n_11187)
);

CKINVDCx11_ASAP7_75t_R g11188 ( 
.A(n_9185),
.Y(n_11188)
);

AOI21xp5_ASAP7_75t_L g11189 ( 
.A1(n_9732),
.A2(n_7689),
.B(n_8894),
.Y(n_11189)
);

INVx1_ASAP7_75t_L g11190 ( 
.A(n_9181),
.Y(n_11190)
);

INVx2_ASAP7_75t_L g11191 ( 
.A(n_9449),
.Y(n_11191)
);

INVx2_ASAP7_75t_L g11192 ( 
.A(n_9449),
.Y(n_11192)
);

BUFx2_ASAP7_75t_L g11193 ( 
.A(n_9686),
.Y(n_11193)
);

OAI21xp5_ASAP7_75t_L g11194 ( 
.A1(n_10058),
.A2(n_8626),
.B(n_8505),
.Y(n_11194)
);

BUFx2_ASAP7_75t_L g11195 ( 
.A(n_9733),
.Y(n_11195)
);

NAND2xp5_ASAP7_75t_SL g11196 ( 
.A(n_9201),
.B(n_8626),
.Y(n_11196)
);

AOI21xp5_ASAP7_75t_L g11197 ( 
.A1(n_9503),
.A2(n_7689),
.B(n_8894),
.Y(n_11197)
);

OR2x6_ASAP7_75t_L g11198 ( 
.A(n_9577),
.B(n_7744),
.Y(n_11198)
);

AOI22xp33_ASAP7_75t_L g11199 ( 
.A1(n_10058),
.A2(n_8219),
.B1(n_8325),
.B2(n_8263),
.Y(n_11199)
);

NAND2xp5_ASAP7_75t_SL g11200 ( 
.A(n_9392),
.B(n_9399),
.Y(n_11200)
);

OA21x2_ASAP7_75t_L g11201 ( 
.A1(n_9690),
.A2(n_8969),
.B(n_8960),
.Y(n_11201)
);

AO31x2_ASAP7_75t_L g11202 ( 
.A1(n_9879),
.A2(n_8537),
.A3(n_8607),
.B(n_8480),
.Y(n_11202)
);

CKINVDCx11_ASAP7_75t_R g11203 ( 
.A(n_9185),
.Y(n_11203)
);

INVx1_ASAP7_75t_L g11204 ( 
.A(n_9181),
.Y(n_11204)
);

INVx3_ASAP7_75t_L g11205 ( 
.A(n_9733),
.Y(n_11205)
);

AOI22xp5_ASAP7_75t_L g11206 ( 
.A1(n_10175),
.A2(n_8219),
.B1(n_8458),
.B2(n_8197),
.Y(n_11206)
);

INVx2_ASAP7_75t_L g11207 ( 
.A(n_9449),
.Y(n_11207)
);

INVx1_ASAP7_75t_SL g11208 ( 
.A(n_9428),
.Y(n_11208)
);

OA21x2_ASAP7_75t_L g11209 ( 
.A1(n_9690),
.A2(n_9693),
.B(n_10098),
.Y(n_11209)
);

HB1xp67_ASAP7_75t_L g11210 ( 
.A(n_8998),
.Y(n_11210)
);

INVx1_ASAP7_75t_L g11211 ( 
.A(n_9181),
.Y(n_11211)
);

OR2x6_ASAP7_75t_L g11212 ( 
.A(n_9577),
.B(n_9756),
.Y(n_11212)
);

OAI21xp5_ASAP7_75t_L g11213 ( 
.A1(n_9196),
.A2(n_8505),
.B(n_8499),
.Y(n_11213)
);

AOI22xp33_ASAP7_75t_L g11214 ( 
.A1(n_10105),
.A2(n_8239),
.B1(n_8468),
.B2(n_8323),
.Y(n_11214)
);

OR2x2_ASAP7_75t_L g11215 ( 
.A(n_9190),
.B(n_8396),
.Y(n_11215)
);

INVx2_ASAP7_75t_L g11216 ( 
.A(n_9449),
.Y(n_11216)
);

AND2x4_ASAP7_75t_L g11217 ( 
.A(n_9733),
.B(n_9773),
.Y(n_11217)
);

BUFx2_ASAP7_75t_L g11218 ( 
.A(n_9733),
.Y(n_11218)
);

INVxp67_ASAP7_75t_SL g11219 ( 
.A(n_9564),
.Y(n_11219)
);

INVx2_ASAP7_75t_L g11220 ( 
.A(n_9449),
.Y(n_11220)
);

AND2x2_ASAP7_75t_L g11221 ( 
.A(n_9519),
.B(n_7864),
.Y(n_11221)
);

AOI21xp5_ASAP7_75t_L g11222 ( 
.A1(n_9503),
.A2(n_7689),
.B(n_8358),
.Y(n_11222)
);

OAI21x1_ASAP7_75t_L g11223 ( 
.A1(n_9893),
.A2(n_9896),
.B(n_9895),
.Y(n_11223)
);

BUFx6f_ASAP7_75t_L g11224 ( 
.A(n_9060),
.Y(n_11224)
);

AND2x2_ASAP7_75t_SL g11225 ( 
.A(n_9959),
.B(n_7849),
.Y(n_11225)
);

NOR2x1_ASAP7_75t_L g11226 ( 
.A(n_8976),
.B(n_8754),
.Y(n_11226)
);

NAND2x1p5_ASAP7_75t_L g11227 ( 
.A(n_9229),
.B(n_8420),
.Y(n_11227)
);

AOI21xp5_ASAP7_75t_L g11228 ( 
.A1(n_9503),
.A2(n_7689),
.B(n_8358),
.Y(n_11228)
);

CKINVDCx5p33_ASAP7_75t_R g11229 ( 
.A(n_9794),
.Y(n_11229)
);

OAI21x1_ASAP7_75t_SL g11230 ( 
.A1(n_8994),
.A2(n_7880),
.B(n_8728),
.Y(n_11230)
);

AO21x2_ASAP7_75t_L g11231 ( 
.A1(n_9939),
.A2(n_8794),
.B(n_8791),
.Y(n_11231)
);

OA21x2_ASAP7_75t_L g11232 ( 
.A1(n_9690),
.A2(n_9693),
.B(n_10098),
.Y(n_11232)
);

INVx1_ASAP7_75t_L g11233 ( 
.A(n_9195),
.Y(n_11233)
);

INVx4_ASAP7_75t_L g11234 ( 
.A(n_9185),
.Y(n_11234)
);

CKINVDCx11_ASAP7_75t_R g11235 ( 
.A(n_9185),
.Y(n_11235)
);

AO21x2_ASAP7_75t_L g11236 ( 
.A1(n_9943),
.A2(n_8794),
.B(n_8791),
.Y(n_11236)
);

AO21x1_ASAP7_75t_L g11237 ( 
.A1(n_9369),
.A2(n_8512),
.B(n_7820),
.Y(n_11237)
);

INVx3_ASAP7_75t_L g11238 ( 
.A(n_9733),
.Y(n_11238)
);

HB1xp67_ASAP7_75t_L g11239 ( 
.A(n_8998),
.Y(n_11239)
);

NAND2xp5_ASAP7_75t_L g11240 ( 
.A(n_9691),
.B(n_9701),
.Y(n_11240)
);

NAND2xp5_ASAP7_75t_L g11241 ( 
.A(n_9701),
.B(n_8677),
.Y(n_11241)
);

NAND2x1p5_ASAP7_75t_L g11242 ( 
.A(n_9229),
.B(n_8420),
.Y(n_11242)
);

NAND3xp33_ASAP7_75t_L g11243 ( 
.A(n_10105),
.B(n_8510),
.C(n_8499),
.Y(n_11243)
);

INVx1_ASAP7_75t_L g11244 ( 
.A(n_9195),
.Y(n_11244)
);

OAI21x1_ASAP7_75t_L g11245 ( 
.A1(n_10176),
.A2(n_8146),
.B(n_8789),
.Y(n_11245)
);

CKINVDCx5p33_ASAP7_75t_R g11246 ( 
.A(n_9795),
.Y(n_11246)
);

INVx1_ASAP7_75t_L g11247 ( 
.A(n_9195),
.Y(n_11247)
);

OAI21x1_ASAP7_75t_L g11248 ( 
.A1(n_10176),
.A2(n_8146),
.B(n_8789),
.Y(n_11248)
);

AND2x2_ASAP7_75t_L g11249 ( 
.A(n_9708),
.B(n_9714),
.Y(n_11249)
);

NAND2xp5_ASAP7_75t_L g11250 ( 
.A(n_9701),
.B(n_8677),
.Y(n_11250)
);

OAI21x1_ASAP7_75t_L g11251 ( 
.A1(n_10176),
.A2(n_8146),
.B(n_8726),
.Y(n_11251)
);

OAI21x1_ASAP7_75t_L g11252 ( 
.A1(n_10176),
.A2(n_8146),
.B(n_8726),
.Y(n_11252)
);

OAI21x1_ASAP7_75t_L g11253 ( 
.A1(n_9895),
.A2(n_9899),
.B(n_9896),
.Y(n_11253)
);

NAND2xp5_ASAP7_75t_L g11254 ( 
.A(n_9179),
.B(n_8072),
.Y(n_11254)
);

OAI21x1_ASAP7_75t_L g11255 ( 
.A1(n_9895),
.A2(n_8146),
.B(n_8683),
.Y(n_11255)
);

INVx1_ASAP7_75t_L g11256 ( 
.A(n_9252),
.Y(n_11256)
);

OAI21xp5_ASAP7_75t_L g11257 ( 
.A1(n_9196),
.A2(n_8529),
.B(n_8510),
.Y(n_11257)
);

AO21x1_ASAP7_75t_L g11258 ( 
.A1(n_9369),
.A2(n_7820),
.B(n_7711),
.Y(n_11258)
);

NAND2xp5_ASAP7_75t_L g11259 ( 
.A(n_9179),
.B(n_9184),
.Y(n_11259)
);

OAI21x1_ASAP7_75t_L g11260 ( 
.A1(n_9895),
.A2(n_9899),
.B(n_9896),
.Y(n_11260)
);

OR2x2_ASAP7_75t_L g11261 ( 
.A(n_9190),
.B(n_8396),
.Y(n_11261)
);

OAI21x1_ASAP7_75t_L g11262 ( 
.A1(n_9895),
.A2(n_8684),
.B(n_8683),
.Y(n_11262)
);

AOI21xp5_ASAP7_75t_L g11263 ( 
.A1(n_9503),
.A2(n_9959),
.B(n_9380),
.Y(n_11263)
);

AO21x2_ASAP7_75t_L g11264 ( 
.A1(n_9943),
.A2(n_9955),
.B(n_9949),
.Y(n_11264)
);

AO21x2_ASAP7_75t_L g11265 ( 
.A1(n_9943),
.A2(n_9955),
.B(n_9949),
.Y(n_11265)
);

NAND2xp5_ASAP7_75t_L g11266 ( 
.A(n_9179),
.B(n_8072),
.Y(n_11266)
);

OAI21x1_ASAP7_75t_L g11267 ( 
.A1(n_9896),
.A2(n_8684),
.B(n_8683),
.Y(n_11267)
);

AOI21xp33_ASAP7_75t_SL g11268 ( 
.A1(n_9392),
.A2(n_8525),
.B(n_8523),
.Y(n_11268)
);

AND2x4_ASAP7_75t_L g11269 ( 
.A(n_9733),
.B(n_7880),
.Y(n_11269)
);

OAI21x1_ASAP7_75t_L g11270 ( 
.A1(n_9896),
.A2(n_8684),
.B(n_8683),
.Y(n_11270)
);

OAI21xp5_ASAP7_75t_L g11271 ( 
.A1(n_9196),
.A2(n_8535),
.B(n_8529),
.Y(n_11271)
);

AOI21xp5_ASAP7_75t_L g11272 ( 
.A1(n_9959),
.A2(n_7689),
.B(n_8730),
.Y(n_11272)
);

BUFx3_ASAP7_75t_L g11273 ( 
.A(n_9131),
.Y(n_11273)
);

INVx1_ASAP7_75t_SL g11274 ( 
.A(n_9497),
.Y(n_11274)
);

AND2x4_ASAP7_75t_L g11275 ( 
.A(n_9773),
.B(n_7880),
.Y(n_11275)
);

BUFx6f_ASAP7_75t_L g11276 ( 
.A(n_9060),
.Y(n_11276)
);

INVx2_ASAP7_75t_L g11277 ( 
.A(n_10179),
.Y(n_11277)
);

AOI21xp5_ASAP7_75t_L g11278 ( 
.A1(n_9959),
.A2(n_7689),
.B(n_8730),
.Y(n_11278)
);

OA21x2_ASAP7_75t_L g11279 ( 
.A1(n_9690),
.A2(n_8974),
.B(n_8679),
.Y(n_11279)
);

INVx8_ASAP7_75t_L g11280 ( 
.A(n_9185),
.Y(n_11280)
);

NOR2xp33_ASAP7_75t_L g11281 ( 
.A(n_9050),
.B(n_8182),
.Y(n_11281)
);

OA21x2_ASAP7_75t_L g11282 ( 
.A1(n_9693),
.A2(n_8974),
.B(n_8679),
.Y(n_11282)
);

INVx1_ASAP7_75t_L g11283 ( 
.A(n_9252),
.Y(n_11283)
);

AO31x2_ASAP7_75t_L g11284 ( 
.A1(n_9764),
.A2(n_8480),
.A3(n_8674),
.B(n_8607),
.Y(n_11284)
);

AOI21xp5_ASAP7_75t_L g11285 ( 
.A1(n_9959),
.A2(n_8736),
.B(n_8843),
.Y(n_11285)
);

INVx1_ASAP7_75t_L g11286 ( 
.A(n_9252),
.Y(n_11286)
);

NAND2x1p5_ASAP7_75t_L g11287 ( 
.A(n_9229),
.B(n_8420),
.Y(n_11287)
);

INVx1_ASAP7_75t_SL g11288 ( 
.A(n_9497),
.Y(n_11288)
);

INVx1_ASAP7_75t_L g11289 ( 
.A(n_9275),
.Y(n_11289)
);

OAI21xp33_ASAP7_75t_L g11290 ( 
.A1(n_10175),
.A2(n_8536),
.B(n_8535),
.Y(n_11290)
);

NAND2xp5_ASAP7_75t_L g11291 ( 
.A(n_9184),
.B(n_8073),
.Y(n_11291)
);

AOI21xp5_ASAP7_75t_L g11292 ( 
.A1(n_9959),
.A2(n_8736),
.B(n_8843),
.Y(n_11292)
);

INVx2_ASAP7_75t_L g11293 ( 
.A(n_10179),
.Y(n_11293)
);

NAND2xp5_ASAP7_75t_L g11294 ( 
.A(n_9184),
.B(n_8073),
.Y(n_11294)
);

CKINVDCx6p67_ASAP7_75t_R g11295 ( 
.A(n_9328),
.Y(n_11295)
);

OA21x2_ASAP7_75t_L g11296 ( 
.A1(n_9693),
.A2(n_8813),
.B(n_8812),
.Y(n_11296)
);

INVx1_ASAP7_75t_L g11297 ( 
.A(n_9275),
.Y(n_11297)
);

NAND2xp5_ASAP7_75t_L g11298 ( 
.A(n_9458),
.B(n_8838),
.Y(n_11298)
);

INVx3_ASAP7_75t_L g11299 ( 
.A(n_9773),
.Y(n_11299)
);

OA21x2_ASAP7_75t_L g11300 ( 
.A1(n_9693),
.A2(n_8813),
.B(n_8812),
.Y(n_11300)
);

INVx1_ASAP7_75t_L g11301 ( 
.A(n_9275),
.Y(n_11301)
);

NAND2xp5_ASAP7_75t_L g11302 ( 
.A(n_9458),
.B(n_8808),
.Y(n_11302)
);

OR2x2_ASAP7_75t_L g11303 ( 
.A(n_9190),
.B(n_8396),
.Y(n_11303)
);

NAND2xp5_ASAP7_75t_SL g11304 ( 
.A(n_9392),
.B(n_9399),
.Y(n_11304)
);

INVx2_ASAP7_75t_L g11305 ( 
.A(n_10179),
.Y(n_11305)
);

INVx1_ASAP7_75t_L g11306 ( 
.A(n_9290),
.Y(n_11306)
);

CKINVDCx16_ASAP7_75t_R g11307 ( 
.A(n_9399),
.Y(n_11307)
);

BUFx2_ASAP7_75t_SL g11308 ( 
.A(n_10017),
.Y(n_11308)
);

NAND2xp5_ASAP7_75t_L g11309 ( 
.A(n_9458),
.B(n_8808),
.Y(n_11309)
);

OAI21xp5_ASAP7_75t_L g11310 ( 
.A1(n_9196),
.A2(n_8540),
.B(n_8536),
.Y(n_11310)
);

AO21x2_ASAP7_75t_L g11311 ( 
.A1(n_9949),
.A2(n_8803),
.B(n_8798),
.Y(n_11311)
);

NAND2x1p5_ASAP7_75t_L g11312 ( 
.A(n_9229),
.B(n_8420),
.Y(n_11312)
);

INVx1_ASAP7_75t_L g11313 ( 
.A(n_9290),
.Y(n_11313)
);

HB1xp67_ASAP7_75t_L g11314 ( 
.A(n_8998),
.Y(n_11314)
);

INVx3_ASAP7_75t_L g11315 ( 
.A(n_9773),
.Y(n_11315)
);

NAND2xp5_ASAP7_75t_L g11316 ( 
.A(n_9498),
.B(n_9026),
.Y(n_11316)
);

OA21x2_ASAP7_75t_L g11317 ( 
.A1(n_10098),
.A2(n_8825),
.B(n_8803),
.Y(n_11317)
);

NAND2xp5_ASAP7_75t_L g11318 ( 
.A(n_9498),
.B(n_8258),
.Y(n_11318)
);

NAND2xp5_ASAP7_75t_L g11319 ( 
.A(n_9498),
.B(n_8258),
.Y(n_11319)
);

AND2x4_ASAP7_75t_L g11320 ( 
.A(n_9773),
.B(n_7880),
.Y(n_11320)
);

NAND2xp5_ASAP7_75t_L g11321 ( 
.A(n_9026),
.B(n_8312),
.Y(n_11321)
);

OA21x2_ASAP7_75t_L g11322 ( 
.A1(n_10098),
.A2(n_8825),
.B(n_8806),
.Y(n_11322)
);

NOR2xp33_ASAP7_75t_L g11323 ( 
.A(n_9369),
.B(n_8312),
.Y(n_11323)
);

INVxp67_ASAP7_75t_L g11324 ( 
.A(n_9530),
.Y(n_11324)
);

INVx2_ASAP7_75t_L g11325 ( 
.A(n_10179),
.Y(n_11325)
);

OA21x2_ASAP7_75t_L g11326 ( 
.A1(n_10098),
.A2(n_8806),
.B(n_8798),
.Y(n_11326)
);

NAND2x1p5_ASAP7_75t_L g11327 ( 
.A(n_9229),
.B(n_8420),
.Y(n_11327)
);

INVx1_ASAP7_75t_L g11328 ( 
.A(n_9290),
.Y(n_11328)
);

NAND2xp5_ASAP7_75t_L g11329 ( 
.A(n_9026),
.B(n_8641),
.Y(n_11329)
);

AO21x2_ASAP7_75t_L g11330 ( 
.A1(n_9949),
.A2(n_8811),
.B(n_8495),
.Y(n_11330)
);

INVx1_ASAP7_75t_L g11331 ( 
.A(n_9315),
.Y(n_11331)
);

INVx1_ASAP7_75t_L g11332 ( 
.A(n_9315),
.Y(n_11332)
);

INVx2_ASAP7_75t_SL g11333 ( 
.A(n_9577),
.Y(n_11333)
);

NOR2xp33_ASAP7_75t_L g11334 ( 
.A(n_9367),
.B(n_8468),
.Y(n_11334)
);

OA21x2_ASAP7_75t_L g11335 ( 
.A1(n_10108),
.A2(n_8811),
.B(n_8704),
.Y(n_11335)
);

AND2x2_ASAP7_75t_L g11336 ( 
.A(n_9708),
.B(n_8113),
.Y(n_11336)
);

OR2x6_ASAP7_75t_L g11337 ( 
.A(n_9577),
.B(n_7798),
.Y(n_11337)
);

BUFx2_ASAP7_75t_L g11338 ( 
.A(n_9773),
.Y(n_11338)
);

INVx1_ASAP7_75t_L g11339 ( 
.A(n_9315),
.Y(n_11339)
);

OR2x2_ASAP7_75t_L g11340 ( 
.A(n_9541),
.B(n_8396),
.Y(n_11340)
);

AO21x2_ASAP7_75t_L g11341 ( 
.A1(n_9955),
.A2(n_8495),
.B(n_8752),
.Y(n_11341)
);

AND2x2_ASAP7_75t_L g11342 ( 
.A(n_9708),
.B(n_8113),
.Y(n_11342)
);

AOI21xp5_ASAP7_75t_L g11343 ( 
.A1(n_9379),
.A2(n_9380),
.B(n_10018),
.Y(n_11343)
);

INVx3_ASAP7_75t_L g11344 ( 
.A(n_9783),
.Y(n_11344)
);

AOI21xp5_ASAP7_75t_L g11345 ( 
.A1(n_9379),
.A2(n_7691),
.B(n_7688),
.Y(n_11345)
);

INVx1_ASAP7_75t_L g11346 ( 
.A(n_9419),
.Y(n_11346)
);

OA21x2_ASAP7_75t_L g11347 ( 
.A1(n_10108),
.A2(n_8704),
.B(n_8644),
.Y(n_11347)
);

CKINVDCx6p67_ASAP7_75t_R g11348 ( 
.A(n_9328),
.Y(n_11348)
);

AO31x2_ASAP7_75t_L g11349 ( 
.A1(n_9714),
.A2(n_8674),
.A3(n_8760),
.B(n_8607),
.Y(n_11349)
);

OAI21xp5_ASAP7_75t_L g11350 ( 
.A1(n_8976),
.A2(n_8545),
.B(n_8540),
.Y(n_11350)
);

OAI21xp5_ASAP7_75t_L g11351 ( 
.A1(n_8976),
.A2(n_8550),
.B(n_8545),
.Y(n_11351)
);

NAND2x1p5_ASAP7_75t_L g11352 ( 
.A(n_9229),
.B(n_8420),
.Y(n_11352)
);

INVx1_ASAP7_75t_L g11353 ( 
.A(n_9419),
.Y(n_11353)
);

AO31x2_ASAP7_75t_L g11354 ( 
.A1(n_9890),
.A2(n_8674),
.A3(n_8764),
.B(n_8760),
.Y(n_11354)
);

OAI21xp5_ASAP7_75t_L g11355 ( 
.A1(n_8976),
.A2(n_8563),
.B(n_8550),
.Y(n_11355)
);

NAND2xp5_ASAP7_75t_L g11356 ( 
.A(n_9122),
.B(n_8641),
.Y(n_11356)
);

AND2x4_ASAP7_75t_L g11357 ( 
.A(n_9783),
.B(n_8420),
.Y(n_11357)
);

AO21x2_ASAP7_75t_L g11358 ( 
.A1(n_9955),
.A2(n_8495),
.B(n_8752),
.Y(n_11358)
);

AND2x4_ASAP7_75t_L g11359 ( 
.A(n_9783),
.B(n_8420),
.Y(n_11359)
);

NAND3xp33_ASAP7_75t_L g11360 ( 
.A(n_10105),
.B(n_8563),
.C(n_8613),
.Y(n_11360)
);

NAND2x1p5_ASAP7_75t_L g11361 ( 
.A(n_9587),
.B(n_8472),
.Y(n_11361)
);

NAND2x1p5_ASAP7_75t_L g11362 ( 
.A(n_9587),
.B(n_8472),
.Y(n_11362)
);

OA21x2_ASAP7_75t_L g11363 ( 
.A1(n_10108),
.A2(n_8704),
.B(n_8644),
.Y(n_11363)
);

INVx2_ASAP7_75t_L g11364 ( 
.A(n_10179),
.Y(n_11364)
);

AOI22xp33_ASAP7_75t_L g11365 ( 
.A1(n_10105),
.A2(n_8323),
.B1(n_8515),
.B2(n_8695),
.Y(n_11365)
);

INVx1_ASAP7_75t_L g11366 ( 
.A(n_9419),
.Y(n_11366)
);

AO21x2_ASAP7_75t_L g11367 ( 
.A1(n_9963),
.A2(n_9977),
.B(n_9957),
.Y(n_11367)
);

OAI21x1_ASAP7_75t_L g11368 ( 
.A1(n_9907),
.A2(n_8850),
.B(n_8857),
.Y(n_11368)
);

INVx2_ASAP7_75t_L g11369 ( 
.A(n_10179),
.Y(n_11369)
);

HB1xp67_ASAP7_75t_L g11370 ( 
.A(n_8998),
.Y(n_11370)
);

INVx2_ASAP7_75t_L g11371 ( 
.A(n_9449),
.Y(n_11371)
);

AO21x1_ASAP7_75t_L g11372 ( 
.A1(n_10175),
.A2(n_7820),
.B(n_7711),
.Y(n_11372)
);

OA21x2_ASAP7_75t_L g11373 ( 
.A1(n_10108),
.A2(n_8704),
.B(n_8644),
.Y(n_11373)
);

AND2x2_ASAP7_75t_L g11374 ( 
.A(n_9708),
.B(n_8113),
.Y(n_11374)
);

INVx1_ASAP7_75t_L g11375 ( 
.A(n_9427),
.Y(n_11375)
);

AOI22x1_ASAP7_75t_L g11376 ( 
.A1(n_9399),
.A2(n_8634),
.B1(n_8650),
.B2(n_8525),
.Y(n_11376)
);

INVx2_ASAP7_75t_L g11377 ( 
.A(n_9470),
.Y(n_11377)
);

INVx1_ASAP7_75t_L g11378 ( 
.A(n_9427),
.Y(n_11378)
);

OAI21x1_ASAP7_75t_L g11379 ( 
.A1(n_9907),
.A2(n_8850),
.B(n_8857),
.Y(n_11379)
);

OR2x2_ASAP7_75t_L g11380 ( 
.A(n_9541),
.B(n_8396),
.Y(n_11380)
);

OAI21x1_ASAP7_75t_L g11381 ( 
.A1(n_9907),
.A2(n_8850),
.B(n_8849),
.Y(n_11381)
);

INVx1_ASAP7_75t_L g11382 ( 
.A(n_9427),
.Y(n_11382)
);

NAND2x1_ASAP7_75t_L g11383 ( 
.A(n_9952),
.B(n_8728),
.Y(n_11383)
);

BUFx2_ASAP7_75t_L g11384 ( 
.A(n_9783),
.Y(n_11384)
);

OAI21xp5_ASAP7_75t_L g11385 ( 
.A1(n_8984),
.A2(n_8613),
.B(n_7751),
.Y(n_11385)
);

AND2x2_ASAP7_75t_L g11386 ( 
.A(n_9714),
.B(n_8113),
.Y(n_11386)
);

OAI21x1_ASAP7_75t_L g11387 ( 
.A1(n_9907),
.A2(n_8850),
.B(n_8849),
.Y(n_11387)
);

AOI22xp33_ASAP7_75t_L g11388 ( 
.A1(n_9887),
.A2(n_8515),
.B1(n_8695),
.B2(n_8613),
.Y(n_11388)
);

AND2x2_ASAP7_75t_L g11389 ( 
.A(n_9714),
.B(n_8138),
.Y(n_11389)
);

INVx6_ASAP7_75t_L g11390 ( 
.A(n_9131),
.Y(n_11390)
);

AO21x1_ASAP7_75t_L g11391 ( 
.A1(n_10175),
.A2(n_7834),
.B(n_7711),
.Y(n_11391)
);

HB1xp67_ASAP7_75t_L g11392 ( 
.A(n_8998),
.Y(n_11392)
);

INVx4_ASAP7_75t_L g11393 ( 
.A(n_9328),
.Y(n_11393)
);

NAND2xp5_ASAP7_75t_L g11394 ( 
.A(n_9122),
.B(n_8643),
.Y(n_11394)
);

NAND3xp33_ASAP7_75t_L g11395 ( 
.A(n_9887),
.B(n_8614),
.C(n_8148),
.Y(n_11395)
);

INVxp67_ASAP7_75t_SL g11396 ( 
.A(n_9564),
.Y(n_11396)
);

OAI22xp5_ASAP7_75t_L g11397 ( 
.A1(n_9689),
.A2(n_8620),
.B1(n_8816),
.B2(n_8632),
.Y(n_11397)
);

OAI21x1_ASAP7_75t_L g11398 ( 
.A1(n_10166),
.A2(n_8257),
.B(n_8050),
.Y(n_11398)
);

INVx6_ASAP7_75t_L g11399 ( 
.A(n_9175),
.Y(n_11399)
);

AND2x2_ASAP7_75t_L g11400 ( 
.A(n_9764),
.B(n_8138),
.Y(n_11400)
);

AOI21xp5_ASAP7_75t_L g11401 ( 
.A1(n_9379),
.A2(n_7691),
.B(n_7688),
.Y(n_11401)
);

INVx1_ASAP7_75t_L g11402 ( 
.A(n_9485),
.Y(n_11402)
);

NAND2xp5_ASAP7_75t_L g11403 ( 
.A(n_9122),
.B(n_8643),
.Y(n_11403)
);

AND2x2_ASAP7_75t_L g11404 ( 
.A(n_9764),
.B(n_8138),
.Y(n_11404)
);

BUFx3_ASAP7_75t_L g11405 ( 
.A(n_9175),
.Y(n_11405)
);

OAI21x1_ASAP7_75t_L g11406 ( 
.A1(n_10171),
.A2(n_8145),
.B(n_8080),
.Y(n_11406)
);

INVx1_ASAP7_75t_L g11407 ( 
.A(n_9485),
.Y(n_11407)
);

OR2x2_ASAP7_75t_L g11408 ( 
.A(n_9541),
.B(n_8287),
.Y(n_11408)
);

BUFx2_ASAP7_75t_R g11409 ( 
.A(n_9236),
.Y(n_11409)
);

INVx6_ASAP7_75t_L g11410 ( 
.A(n_9175),
.Y(n_11410)
);

OAI21x1_ASAP7_75t_L g11411 ( 
.A1(n_10171),
.A2(n_9926),
.B(n_9913),
.Y(n_11411)
);

AOI21xp5_ASAP7_75t_L g11412 ( 
.A1(n_9380),
.A2(n_7755),
.B(n_8148),
.Y(n_11412)
);

NAND2xp5_ASAP7_75t_L g11413 ( 
.A(n_9142),
.B(n_8666),
.Y(n_11413)
);

NAND2xp5_ASAP7_75t_L g11414 ( 
.A(n_9142),
.B(n_8666),
.Y(n_11414)
);

OAI21x1_ASAP7_75t_L g11415 ( 
.A1(n_9913),
.A2(n_8145),
.B(n_8080),
.Y(n_11415)
);

OAI21x1_ASAP7_75t_L g11416 ( 
.A1(n_9913),
.A2(n_9928),
.B(n_9926),
.Y(n_11416)
);

OAI21x1_ASAP7_75t_L g11417 ( 
.A1(n_9913),
.A2(n_8145),
.B(n_8080),
.Y(n_11417)
);

OAI22xp5_ASAP7_75t_L g11418 ( 
.A1(n_9689),
.A2(n_8620),
.B1(n_8816),
.B2(n_8632),
.Y(n_11418)
);

OAI22xp5_ASAP7_75t_L g11419 ( 
.A1(n_9689),
.A2(n_8620),
.B1(n_8816),
.B2(n_8632),
.Y(n_11419)
);

NAND2xp5_ASAP7_75t_L g11420 ( 
.A(n_9142),
.B(n_8666),
.Y(n_11420)
);

HB1xp67_ASAP7_75t_L g11421 ( 
.A(n_8998),
.Y(n_11421)
);

INVx1_ASAP7_75t_L g11422 ( 
.A(n_9485),
.Y(n_11422)
);

INVx1_ASAP7_75t_L g11423 ( 
.A(n_8979),
.Y(n_11423)
);

AOI21xp5_ASAP7_75t_L g11424 ( 
.A1(n_10018),
.A2(n_7755),
.B(n_8831),
.Y(n_11424)
);

OAI21x1_ASAP7_75t_L g11425 ( 
.A1(n_9913),
.A2(n_8050),
.B(n_8034),
.Y(n_11425)
);

OAI21x1_ASAP7_75t_L g11426 ( 
.A1(n_9926),
.A2(n_8050),
.B(n_8034),
.Y(n_11426)
);

AOI211xp5_ASAP7_75t_L g11427 ( 
.A1(n_9178),
.A2(n_8688),
.B(n_8568),
.C(n_8210),
.Y(n_11427)
);

OAI21xp5_ASAP7_75t_L g11428 ( 
.A1(n_8984),
.A2(n_7703),
.B(n_7700),
.Y(n_11428)
);

INVx1_ASAP7_75t_L g11429 ( 
.A(n_8979),
.Y(n_11429)
);

AOI22xp33_ASAP7_75t_L g11430 ( 
.A1(n_10018),
.A2(n_7703),
.B1(n_7700),
.B2(n_8513),
.Y(n_11430)
);

BUFx10_ASAP7_75t_L g11431 ( 
.A(n_9269),
.Y(n_11431)
);

INVx2_ASAP7_75t_L g11432 ( 
.A(n_9470),
.Y(n_11432)
);

OR2x6_ASAP7_75t_L g11433 ( 
.A(n_9577),
.B(n_7798),
.Y(n_11433)
);

OA21x2_ASAP7_75t_L g11434 ( 
.A1(n_10108),
.A2(n_8792),
.B(n_8729),
.Y(n_11434)
);

NAND2xp5_ASAP7_75t_L g11435 ( 
.A(n_9232),
.B(n_8565),
.Y(n_11435)
);

INVx2_ASAP7_75t_L g11436 ( 
.A(n_9470),
.Y(n_11436)
);

CKINVDCx5p33_ASAP7_75t_R g11437 ( 
.A(n_9795),
.Y(n_11437)
);

OAI21x1_ASAP7_75t_L g11438 ( 
.A1(n_9926),
.A2(n_8034),
.B(n_8050),
.Y(n_11438)
);

OAI21x1_ASAP7_75t_L g11439 ( 
.A1(n_9926),
.A2(n_8034),
.B(n_8080),
.Y(n_11439)
);

NAND2xp5_ASAP7_75t_L g11440 ( 
.A(n_9232),
.B(n_8565),
.Y(n_11440)
);

INVx1_ASAP7_75t_L g11441 ( 
.A(n_8979),
.Y(n_11441)
);

NAND2xp5_ASAP7_75t_L g11442 ( 
.A(n_9232),
.B(n_7916),
.Y(n_11442)
);

NOR2x1_ASAP7_75t_SL g11443 ( 
.A(n_9272),
.B(n_9296),
.Y(n_11443)
);

INVx1_ASAP7_75t_SL g11444 ( 
.A(n_9497),
.Y(n_11444)
);

INVx1_ASAP7_75t_L g11445 ( 
.A(n_8979),
.Y(n_11445)
);

OAI21x1_ASAP7_75t_L g11446 ( 
.A1(n_9928),
.A2(n_9930),
.B(n_9929),
.Y(n_11446)
);

BUFx3_ASAP7_75t_L g11447 ( 
.A(n_9175),
.Y(n_11447)
);

OAI21x1_ASAP7_75t_L g11448 ( 
.A1(n_9928),
.A2(n_8034),
.B(n_8080),
.Y(n_11448)
);

OAI21x1_ASAP7_75t_L g11449 ( 
.A1(n_9928),
.A2(n_8429),
.B(n_8243),
.Y(n_11449)
);

INVx1_ASAP7_75t_L g11450 ( 
.A(n_8987),
.Y(n_11450)
);

INVx1_ASAP7_75t_L g11451 ( 
.A(n_8987),
.Y(n_11451)
);

AO31x2_ASAP7_75t_L g11452 ( 
.A1(n_9764),
.A2(n_9890),
.A3(n_10161),
.B(n_10065),
.Y(n_11452)
);

CKINVDCx20_ASAP7_75t_R g11453 ( 
.A(n_9225),
.Y(n_11453)
);

INVx1_ASAP7_75t_L g11454 ( 
.A(n_8987),
.Y(n_11454)
);

AND2x4_ASAP7_75t_L g11455 ( 
.A(n_9783),
.B(n_8472),
.Y(n_11455)
);

INVx1_ASAP7_75t_L g11456 ( 
.A(n_8987),
.Y(n_11456)
);

INVx1_ASAP7_75t_SL g11457 ( 
.A(n_9511),
.Y(n_11457)
);

AND2x2_ASAP7_75t_L g11458 ( 
.A(n_9890),
.B(n_8138),
.Y(n_11458)
);

INVx1_ASAP7_75t_L g11459 ( 
.A(n_8989),
.Y(n_11459)
);

CKINVDCx20_ASAP7_75t_R g11460 ( 
.A(n_9423),
.Y(n_11460)
);

AND2x2_ASAP7_75t_L g11461 ( 
.A(n_9890),
.B(n_8904),
.Y(n_11461)
);

INVx1_ASAP7_75t_L g11462 ( 
.A(n_8989),
.Y(n_11462)
);

BUFx8_ASAP7_75t_L g11463 ( 
.A(n_9328),
.Y(n_11463)
);

AOI21xp5_ASAP7_75t_L g11464 ( 
.A1(n_10018),
.A2(n_8836),
.B(n_8831),
.Y(n_11464)
);

AOI21xp5_ASAP7_75t_L g11465 ( 
.A1(n_10018),
.A2(n_8842),
.B(n_8836),
.Y(n_11465)
);

AOI22xp33_ASAP7_75t_SL g11466 ( 
.A1(n_9689),
.A2(n_7831),
.B1(n_8124),
.B2(n_7849),
.Y(n_11466)
);

OAI21x1_ASAP7_75t_L g11467 ( 
.A1(n_10171),
.A2(n_8243),
.B(n_8145),
.Y(n_11467)
);

INVx1_ASAP7_75t_L g11468 ( 
.A(n_8989),
.Y(n_11468)
);

BUFx6f_ASAP7_75t_L g11469 ( 
.A(n_9060),
.Y(n_11469)
);

AND2x2_ASAP7_75t_L g11470 ( 
.A(n_9706),
.B(n_8904),
.Y(n_11470)
);

BUFx3_ASAP7_75t_L g11471 ( 
.A(n_9175),
.Y(n_11471)
);

NAND2xp5_ASAP7_75t_L g11472 ( 
.A(n_9118),
.B(n_7916),
.Y(n_11472)
);

NAND2xp5_ASAP7_75t_L g11473 ( 
.A(n_9118),
.B(n_9580),
.Y(n_11473)
);

INVx1_ASAP7_75t_L g11474 ( 
.A(n_8989),
.Y(n_11474)
);

OAI21xp5_ASAP7_75t_L g11475 ( 
.A1(n_8984),
.A2(n_8548),
.B(n_8485),
.Y(n_11475)
);

AOI21xp5_ASAP7_75t_L g11476 ( 
.A1(n_10018),
.A2(n_8842),
.B(n_7690),
.Y(n_11476)
);

AOI21x1_ASAP7_75t_L g11477 ( 
.A1(n_9963),
.A2(n_8951),
.B(n_8902),
.Y(n_11477)
);

BUFx6f_ASAP7_75t_L g11478 ( 
.A(n_9060),
.Y(n_11478)
);

OAI21x1_ASAP7_75t_L g11479 ( 
.A1(n_9928),
.A2(n_8145),
.B(n_8243),
.Y(n_11479)
);

OAI21xp5_ASAP7_75t_L g11480 ( 
.A1(n_8984),
.A2(n_9882),
.B(n_9258),
.Y(n_11480)
);

INVxp67_ASAP7_75t_SL g11481 ( 
.A(n_9564),
.Y(n_11481)
);

OA21x2_ASAP7_75t_L g11482 ( 
.A1(n_10119),
.A2(n_8792),
.B(n_8729),
.Y(n_11482)
);

OAI21x1_ASAP7_75t_L g11483 ( 
.A1(n_9929),
.A2(n_8257),
.B(n_8243),
.Y(n_11483)
);

OAI21xp5_ASAP7_75t_L g11484 ( 
.A1(n_9882),
.A2(n_9258),
.B(n_9254),
.Y(n_11484)
);

BUFx3_ASAP7_75t_L g11485 ( 
.A(n_9175),
.Y(n_11485)
);

O2A1O1Ixp33_ASAP7_75t_L g11486 ( 
.A1(n_9882),
.A2(n_9178),
.B(n_9220),
.C(n_9365),
.Y(n_11486)
);

OAI22xp5_ASAP7_75t_SL g11487 ( 
.A1(n_10148),
.A2(n_9626),
.B1(n_9423),
.B2(n_9178),
.Y(n_11487)
);

INVx1_ASAP7_75t_L g11488 ( 
.A(n_8993),
.Y(n_11488)
);

AND2x2_ASAP7_75t_L g11489 ( 
.A(n_9706),
.B(n_8904),
.Y(n_11489)
);

AND2x2_ASAP7_75t_L g11490 ( 
.A(n_9706),
.B(n_8904),
.Y(n_11490)
);

AOI21xp5_ASAP7_75t_L g11491 ( 
.A1(n_10018),
.A2(n_7690),
.B(n_7684),
.Y(n_11491)
);

INVx2_ASAP7_75t_L g11492 ( 
.A(n_9470),
.Y(n_11492)
);

OAI21x1_ASAP7_75t_L g11493 ( 
.A1(n_9929),
.A2(n_8509),
.B(n_8257),
.Y(n_11493)
);

BUFx2_ASAP7_75t_L g11494 ( 
.A(n_9783),
.Y(n_11494)
);

OAI21xp5_ASAP7_75t_L g11495 ( 
.A1(n_9254),
.A2(n_8548),
.B(n_8485),
.Y(n_11495)
);

OAI21xp5_ASAP7_75t_L g11496 ( 
.A1(n_9254),
.A2(n_8492),
.B(n_8471),
.Y(n_11496)
);

OAI21xp5_ASAP7_75t_L g11497 ( 
.A1(n_9258),
.A2(n_8492),
.B(n_8614),
.Y(n_11497)
);

INVx3_ASAP7_75t_L g11498 ( 
.A(n_9831),
.Y(n_11498)
);

AO31x2_ASAP7_75t_L g11499 ( 
.A1(n_10065),
.A2(n_8764),
.A3(n_8774),
.B(n_8760),
.Y(n_11499)
);

OA21x2_ASAP7_75t_L g11500 ( 
.A1(n_10119),
.A2(n_8792),
.B(n_8729),
.Y(n_11500)
);

INVx1_ASAP7_75t_L g11501 ( 
.A(n_8993),
.Y(n_11501)
);

AO21x2_ASAP7_75t_L g11502 ( 
.A1(n_9963),
.A2(n_8495),
.B(n_8752),
.Y(n_11502)
);

AND2x2_ASAP7_75t_L g11503 ( 
.A(n_9706),
.B(n_8756),
.Y(n_11503)
);

AOI21x1_ASAP7_75t_L g11504 ( 
.A1(n_9963),
.A2(n_8967),
.B(n_8957),
.Y(n_11504)
);

OAI21x1_ASAP7_75t_L g11505 ( 
.A1(n_9929),
.A2(n_8257),
.B(n_8243),
.Y(n_11505)
);

AOI21x1_ASAP7_75t_L g11506 ( 
.A1(n_9977),
.A2(n_8957),
.B(n_8967),
.Y(n_11506)
);

BUFx2_ASAP7_75t_L g11507 ( 
.A(n_9831),
.Y(n_11507)
);

OAI21x1_ASAP7_75t_L g11508 ( 
.A1(n_9929),
.A2(n_8429),
.B(n_8257),
.Y(n_11508)
);

AND2x4_ASAP7_75t_L g11509 ( 
.A(n_9831),
.B(n_8472),
.Y(n_11509)
);

INVx1_ASAP7_75t_SL g11510 ( 
.A(n_9511),
.Y(n_11510)
);

OAI21x1_ASAP7_75t_L g11511 ( 
.A1(n_9930),
.A2(n_8509),
.B(n_8429),
.Y(n_11511)
);

NAND2xp5_ASAP7_75t_L g11512 ( 
.A(n_9118),
.B(n_7917),
.Y(n_11512)
);

INVx2_ASAP7_75t_L g11513 ( 
.A(n_9470),
.Y(n_11513)
);

AO31x2_ASAP7_75t_L g11514 ( 
.A1(n_10065),
.A2(n_8774),
.A3(n_8780),
.B(n_8764),
.Y(n_11514)
);

OAI21x1_ASAP7_75t_L g11515 ( 
.A1(n_9930),
.A2(n_8509),
.B(n_8429),
.Y(n_11515)
);

OAI21x1_ASAP7_75t_L g11516 ( 
.A1(n_9930),
.A2(n_8509),
.B(n_8429),
.Y(n_11516)
);

INVx1_ASAP7_75t_L g11517 ( 
.A(n_8993),
.Y(n_11517)
);

CKINVDCx11_ASAP7_75t_R g11518 ( 
.A(n_9328),
.Y(n_11518)
);

OAI21x1_ASAP7_75t_L g11519 ( 
.A1(n_9951),
.A2(n_8274),
.B(n_8178),
.Y(n_11519)
);

BUFx8_ASAP7_75t_L g11520 ( 
.A(n_9328),
.Y(n_11520)
);

INVx2_ASAP7_75t_SL g11521 ( 
.A(n_9577),
.Y(n_11521)
);

AO31x2_ASAP7_75t_L g11522 ( 
.A1(n_10065),
.A2(n_8780),
.A3(n_8799),
.B(n_8774),
.Y(n_11522)
);

OR2x6_ASAP7_75t_L g11523 ( 
.A(n_9756),
.B(n_10027),
.Y(n_11523)
);

INVx1_ASAP7_75t_L g11524 ( 
.A(n_8993),
.Y(n_11524)
);

OAI21x1_ASAP7_75t_L g11525 ( 
.A1(n_10166),
.A2(n_8274),
.B(n_8178),
.Y(n_11525)
);

OAI21xp5_ASAP7_75t_L g11526 ( 
.A1(n_9258),
.A2(n_8754),
.B(n_8055),
.Y(n_11526)
);

HB1xp67_ASAP7_75t_L g11527 ( 
.A(n_8998),
.Y(n_11527)
);

OAI21x1_ASAP7_75t_L g11528 ( 
.A1(n_9951),
.A2(n_8274),
.B(n_8178),
.Y(n_11528)
);

CKINVDCx5p33_ASAP7_75t_R g11529 ( 
.A(n_9795),
.Y(n_11529)
);

INVx1_ASAP7_75t_L g11530 ( 
.A(n_8996),
.Y(n_11530)
);

OAI21x1_ASAP7_75t_L g11531 ( 
.A1(n_9951),
.A2(n_8274),
.B(n_8178),
.Y(n_11531)
);

INVx3_ASAP7_75t_L g11532 ( 
.A(n_9831),
.Y(n_11532)
);

OAI21x1_ASAP7_75t_L g11533 ( 
.A1(n_9951),
.A2(n_9961),
.B(n_9958),
.Y(n_11533)
);

OA21x2_ASAP7_75t_L g11534 ( 
.A1(n_10119),
.A2(n_9817),
.B(n_9812),
.Y(n_11534)
);

AO31x2_ASAP7_75t_L g11535 ( 
.A1(n_10161),
.A2(n_8780),
.A3(n_8799),
.B(n_8919),
.Y(n_11535)
);

INVx2_ASAP7_75t_SL g11536 ( 
.A(n_9756),
.Y(n_11536)
);

INVx1_ASAP7_75t_L g11537 ( 
.A(n_8996),
.Y(n_11537)
);

INVx1_ASAP7_75t_L g11538 ( 
.A(n_8996),
.Y(n_11538)
);

INVx3_ASAP7_75t_L g11539 ( 
.A(n_9831),
.Y(n_11539)
);

AOI22xp33_ASAP7_75t_L g11540 ( 
.A1(n_10018),
.A2(n_8513),
.B1(n_7831),
.B2(n_8124),
.Y(n_11540)
);

NOR2x1_ASAP7_75t_SL g11541 ( 
.A(n_9296),
.B(n_8542),
.Y(n_11541)
);

OAI21x1_ASAP7_75t_L g11542 ( 
.A1(n_9951),
.A2(n_8274),
.B(n_8178),
.Y(n_11542)
);

HB1xp67_ASAP7_75t_L g11543 ( 
.A(n_8998),
.Y(n_11543)
);

OR2x2_ASAP7_75t_L g11544 ( 
.A(n_9541),
.B(n_8287),
.Y(n_11544)
);

INVx1_ASAP7_75t_L g11545 ( 
.A(n_8996),
.Y(n_11545)
);

OAI21x1_ASAP7_75t_SL g11546 ( 
.A1(n_8994),
.A2(n_8728),
.B(n_8709),
.Y(n_11546)
);

INVx1_ASAP7_75t_L g11547 ( 
.A(n_9000),
.Y(n_11547)
);

INVx1_ASAP7_75t_L g11548 ( 
.A(n_9000),
.Y(n_11548)
);

INVx3_ASAP7_75t_L g11549 ( 
.A(n_9831),
.Y(n_11549)
);

INVx2_ASAP7_75t_L g11550 ( 
.A(n_9470),
.Y(n_11550)
);

OAI21x1_ASAP7_75t_L g11551 ( 
.A1(n_9958),
.A2(n_8299),
.B(n_8178),
.Y(n_11551)
);

OAI21x1_ASAP7_75t_L g11552 ( 
.A1(n_9958),
.A2(n_8315),
.B(n_8299),
.Y(n_11552)
);

OAI21x1_ASAP7_75t_L g11553 ( 
.A1(n_9958),
.A2(n_8315),
.B(n_8299),
.Y(n_11553)
);

OR2x2_ASAP7_75t_L g11554 ( 
.A(n_9541),
.B(n_9597),
.Y(n_11554)
);

OAI21x1_ASAP7_75t_L g11555 ( 
.A1(n_9958),
.A2(n_8315),
.B(n_8299),
.Y(n_11555)
);

INVx5_ASAP7_75t_L g11556 ( 
.A(n_10148),
.Y(n_11556)
);

AOI22xp33_ASAP7_75t_L g11557 ( 
.A1(n_10070),
.A2(n_8513),
.B1(n_7831),
.B2(n_8124),
.Y(n_11557)
);

AOI21xp5_ASAP7_75t_L g11558 ( 
.A1(n_10070),
.A2(n_7694),
.B(n_7684),
.Y(n_11558)
);

INVx2_ASAP7_75t_L g11559 ( 
.A(n_9470),
.Y(n_11559)
);

INVx2_ASAP7_75t_L g11560 ( 
.A(n_9470),
.Y(n_11560)
);

OAI21x1_ASAP7_75t_L g11561 ( 
.A1(n_9961),
.A2(n_8315),
.B(n_8299),
.Y(n_11561)
);

AOI21x1_ASAP7_75t_L g11562 ( 
.A1(n_9977),
.A2(n_7729),
.B(n_7727),
.Y(n_11562)
);

AO31x2_ASAP7_75t_L g11563 ( 
.A1(n_10161),
.A2(n_8799),
.A3(n_8919),
.B(n_8841),
.Y(n_11563)
);

AOI21x1_ASAP7_75t_L g11564 ( 
.A1(n_9977),
.A2(n_7729),
.B(n_7727),
.Y(n_11564)
);

INVx3_ASAP7_75t_L g11565 ( 
.A(n_10036),
.Y(n_11565)
);

HB1xp67_ASAP7_75t_L g11566 ( 
.A(n_8998),
.Y(n_11566)
);

NAND2xp5_ASAP7_75t_L g11567 ( 
.A(n_9580),
.B(n_7917),
.Y(n_11567)
);

NAND2xp5_ASAP7_75t_L g11568 ( 
.A(n_9580),
.B(n_7898),
.Y(n_11568)
);

AO21x2_ASAP7_75t_L g11569 ( 
.A1(n_9957),
.A2(n_8495),
.B(n_8820),
.Y(n_11569)
);

OAI21x1_ASAP7_75t_L g11570 ( 
.A1(n_10166),
.A2(n_8315),
.B(n_8750),
.Y(n_11570)
);

OAI21x1_ASAP7_75t_L g11571 ( 
.A1(n_10166),
.A2(n_8771),
.B(n_8750),
.Y(n_11571)
);

OAI21x1_ASAP7_75t_L g11572 ( 
.A1(n_10166),
.A2(n_8772),
.B(n_8771),
.Y(n_11572)
);

OAI21x1_ASAP7_75t_L g11573 ( 
.A1(n_9961),
.A2(n_8773),
.B(n_8772),
.Y(n_11573)
);

INVx1_ASAP7_75t_L g11574 ( 
.A(n_9000),
.Y(n_11574)
);

NAND2x1p5_ASAP7_75t_L g11575 ( 
.A(n_9587),
.B(n_8472),
.Y(n_11575)
);

INVx4_ASAP7_75t_L g11576 ( 
.A(n_9025),
.Y(n_11576)
);

AND2x4_ASAP7_75t_L g11577 ( 
.A(n_9715),
.B(n_8472),
.Y(n_11577)
);

INVx2_ASAP7_75t_L g11578 ( 
.A(n_9548),
.Y(n_11578)
);

AO21x2_ASAP7_75t_L g11579 ( 
.A1(n_9957),
.A2(n_8495),
.B(n_8820),
.Y(n_11579)
);

OAI21x1_ASAP7_75t_L g11580 ( 
.A1(n_9961),
.A2(n_8778),
.B(n_8773),
.Y(n_11580)
);

NOR2xp33_ASAP7_75t_L g11581 ( 
.A(n_9367),
.B(n_8100),
.Y(n_11581)
);

INVx1_ASAP7_75t_L g11582 ( 
.A(n_9000),
.Y(n_11582)
);

OAI21x1_ASAP7_75t_L g11583 ( 
.A1(n_9964),
.A2(n_8800),
.B(n_8778),
.Y(n_11583)
);

OAI21xp5_ASAP7_75t_L g11584 ( 
.A1(n_9202),
.A2(n_8754),
.B(n_8055),
.Y(n_11584)
);

AO21x2_ASAP7_75t_L g11585 ( 
.A1(n_9957),
.A2(n_8820),
.B(n_8846),
.Y(n_11585)
);

INVx3_ASAP7_75t_L g11586 ( 
.A(n_10036),
.Y(n_11586)
);

BUFx3_ASAP7_75t_L g11587 ( 
.A(n_9175),
.Y(n_11587)
);

BUFx2_ASAP7_75t_L g11588 ( 
.A(n_9845),
.Y(n_11588)
);

INVx1_ASAP7_75t_L g11589 ( 
.A(n_9020),
.Y(n_11589)
);

HB1xp67_ASAP7_75t_L g11590 ( 
.A(n_8998),
.Y(n_11590)
);

AND2x4_ASAP7_75t_L g11591 ( 
.A(n_9715),
.B(n_8472),
.Y(n_11591)
);

INVx1_ASAP7_75t_L g11592 ( 
.A(n_9020),
.Y(n_11592)
);

OR3x4_ASAP7_75t_SL g11593 ( 
.A(n_10041),
.B(n_8688),
.C(n_8210),
.Y(n_11593)
);

AO31x2_ASAP7_75t_L g11594 ( 
.A1(n_10161),
.A2(n_8919),
.A3(n_8841),
.B(n_8818),
.Y(n_11594)
);

OAI21x1_ASAP7_75t_L g11595 ( 
.A1(n_9964),
.A2(n_8802),
.B(n_8800),
.Y(n_11595)
);

OAI21x1_ASAP7_75t_L g11596 ( 
.A1(n_9964),
.A2(n_8805),
.B(n_8802),
.Y(n_11596)
);

AND2x4_ASAP7_75t_L g11597 ( 
.A(n_9715),
.B(n_9750),
.Y(n_11597)
);

OAI21x1_ASAP7_75t_SL g11598 ( 
.A1(n_9233),
.A2(n_8709),
.B(n_8702),
.Y(n_11598)
);

INVxp67_ASAP7_75t_L g11599 ( 
.A(n_9530),
.Y(n_11599)
);

AOI21xp5_ASAP7_75t_L g11600 ( 
.A1(n_10070),
.A2(n_7698),
.B(n_7694),
.Y(n_11600)
);

NAND2xp5_ASAP7_75t_L g11601 ( 
.A(n_9599),
.B(n_7898),
.Y(n_11601)
);

AOI21xp5_ASAP7_75t_L g11602 ( 
.A1(n_10070),
.A2(n_7713),
.B(n_7698),
.Y(n_11602)
);

AO21x2_ASAP7_75t_L g11603 ( 
.A1(n_9957),
.A2(n_8846),
.B(n_8955),
.Y(n_11603)
);

OAI21x1_ASAP7_75t_L g11604 ( 
.A1(n_9964),
.A2(n_8829),
.B(n_8805),
.Y(n_11604)
);

AO31x2_ASAP7_75t_L g11605 ( 
.A1(n_10172),
.A2(n_10190),
.A3(n_10173),
.B(n_9474),
.Y(n_11605)
);

BUFx8_ASAP7_75t_L g11606 ( 
.A(n_9798),
.Y(n_11606)
);

OAI21x1_ASAP7_75t_L g11607 ( 
.A1(n_9964),
.A2(n_8829),
.B(n_8839),
.Y(n_11607)
);

INVx1_ASAP7_75t_SL g11608 ( 
.A(n_9511),
.Y(n_11608)
);

OAI21x1_ASAP7_75t_L g11609 ( 
.A1(n_10062),
.A2(n_8839),
.B(n_8661),
.Y(n_11609)
);

NAND2x1p5_ASAP7_75t_L g11610 ( 
.A(n_9587),
.B(n_8472),
.Y(n_11610)
);

AOI21xp5_ASAP7_75t_L g11611 ( 
.A1(n_10070),
.A2(n_7724),
.B(n_7713),
.Y(n_11611)
);

HB1xp67_ASAP7_75t_L g11612 ( 
.A(n_8998),
.Y(n_11612)
);

AO21x1_ASAP7_75t_L g11613 ( 
.A1(n_9854),
.A2(n_7872),
.B(n_7834),
.Y(n_11613)
);

INVx2_ASAP7_75t_L g11614 ( 
.A(n_9548),
.Y(n_11614)
);

BUFx10_ASAP7_75t_L g11615 ( 
.A(n_9269),
.Y(n_11615)
);

NAND2x1p5_ASAP7_75t_L g11616 ( 
.A(n_9587),
.B(n_8472),
.Y(n_11616)
);

AO31x2_ASAP7_75t_L g11617 ( 
.A1(n_10172),
.A2(n_8818),
.A3(n_8929),
.B(n_8833),
.Y(n_11617)
);

INVx1_ASAP7_75t_L g11618 ( 
.A(n_9020),
.Y(n_11618)
);

AO31x2_ASAP7_75t_L g11619 ( 
.A1(n_10172),
.A2(n_8971),
.A3(n_8948),
.B(n_8912),
.Y(n_11619)
);

NAND2xp5_ASAP7_75t_L g11620 ( 
.A(n_9599),
.B(n_7899),
.Y(n_11620)
);

NAND2xp5_ASAP7_75t_SL g11621 ( 
.A(n_9175),
.B(n_7782),
.Y(n_11621)
);

A2O1A1Ixp33_ASAP7_75t_L g11622 ( 
.A1(n_9365),
.A2(n_9202),
.B(n_9061),
.C(n_9248),
.Y(n_11622)
);

AND2x4_ASAP7_75t_L g11623 ( 
.A(n_9715),
.B(n_8472),
.Y(n_11623)
);

AND2x4_ASAP7_75t_L g11624 ( 
.A(n_9750),
.B(n_7901),
.Y(n_11624)
);

BUFx2_ASAP7_75t_L g11625 ( 
.A(n_9845),
.Y(n_11625)
);

OAI21x1_ASAP7_75t_L g11626 ( 
.A1(n_10062),
.A2(n_8839),
.B(n_8661),
.Y(n_11626)
);

AO21x2_ASAP7_75t_L g11627 ( 
.A1(n_9957),
.A2(n_8846),
.B(n_8955),
.Y(n_11627)
);

AND2x4_ASAP7_75t_L g11628 ( 
.A(n_9750),
.B(n_8405),
.Y(n_11628)
);

INVx1_ASAP7_75t_L g11629 ( 
.A(n_10196),
.Y(n_11629)
);

OR2x2_ASAP7_75t_L g11630 ( 
.A(n_10324),
.B(n_9901),
.Y(n_11630)
);

OAI22xp5_ASAP7_75t_L g11631 ( 
.A1(n_10981),
.A2(n_9202),
.B1(n_9061),
.B2(n_9262),
.Y(n_11631)
);

OR2x2_ASAP7_75t_L g11632 ( 
.A(n_10324),
.B(n_9901),
.Y(n_11632)
);

AND2x2_ASAP7_75t_L g11633 ( 
.A(n_10708),
.B(n_9538),
.Y(n_11633)
);

NAND2xp5_ASAP7_75t_L g11634 ( 
.A(n_10816),
.B(n_9374),
.Y(n_11634)
);

CKINVDCx16_ASAP7_75t_R g11635 ( 
.A(n_10263),
.Y(n_11635)
);

AOI21xp5_ASAP7_75t_SL g11636 ( 
.A1(n_10329),
.A2(n_9585),
.B(n_9440),
.Y(n_11636)
);

HB1xp67_ASAP7_75t_L g11637 ( 
.A(n_10470),
.Y(n_11637)
);

O2A1O1Ixp33_ASAP7_75t_L g11638 ( 
.A1(n_10694),
.A2(n_9178),
.B(n_9177),
.C(n_9036),
.Y(n_11638)
);

AND2x2_ASAP7_75t_L g11639 ( 
.A(n_10708),
.B(n_9538),
.Y(n_11639)
);

AOI21xp5_ASAP7_75t_SL g11640 ( 
.A1(n_10329),
.A2(n_9585),
.B(n_9440),
.Y(n_11640)
);

NOR2xp67_ASAP7_75t_L g11641 ( 
.A(n_10247),
.B(n_11012),
.Y(n_11641)
);

O2A1O1Ixp33_ASAP7_75t_L g11642 ( 
.A1(n_10694),
.A2(n_10752),
.B(n_10291),
.C(n_10886),
.Y(n_11642)
);

INVx1_ASAP7_75t_L g11643 ( 
.A(n_10196),
.Y(n_11643)
);

AND2x2_ASAP7_75t_L g11644 ( 
.A(n_11307),
.B(n_9538),
.Y(n_11644)
);

AOI221x1_ASAP7_75t_SL g11645 ( 
.A1(n_10886),
.A2(n_9506),
.B1(n_9565),
.B2(n_9474),
.C(n_9469),
.Y(n_11645)
);

INVx2_ASAP7_75t_L g11646 ( 
.A(n_10226),
.Y(n_11646)
);

AND2x4_ASAP7_75t_L g11647 ( 
.A(n_10246),
.B(n_9750),
.Y(n_11647)
);

NOR3xp33_ASAP7_75t_L g11648 ( 
.A(n_10981),
.B(n_9262),
.C(n_9755),
.Y(n_11648)
);

A2O1A1Ixp33_ASAP7_75t_L g11649 ( 
.A1(n_10498),
.A2(n_9365),
.B(n_9837),
.C(n_9202),
.Y(n_11649)
);

CKINVDCx5p33_ASAP7_75t_R g11650 ( 
.A(n_10369),
.Y(n_11650)
);

OAI22xp5_ASAP7_75t_L g11651 ( 
.A1(n_10726),
.A2(n_9061),
.B1(n_9262),
.B2(n_9767),
.Y(n_11651)
);

INVx1_ASAP7_75t_L g11652 ( 
.A(n_10197),
.Y(n_11652)
);

INVx1_ASAP7_75t_L g11653 ( 
.A(n_10197),
.Y(n_11653)
);

OAI22xp5_ASAP7_75t_L g11654 ( 
.A1(n_10726),
.A2(n_9061),
.B1(n_9800),
.B2(n_9767),
.Y(n_11654)
);

NAND2xp5_ASAP7_75t_L g11655 ( 
.A(n_10816),
.B(n_9374),
.Y(n_11655)
);

AOI21xp5_ASAP7_75t_SL g11656 ( 
.A1(n_10396),
.A2(n_9585),
.B(n_9440),
.Y(n_11656)
);

HB1xp67_ASAP7_75t_L g11657 ( 
.A(n_10470),
.Y(n_11657)
);

HB1xp67_ASAP7_75t_L g11658 ( 
.A(n_10476),
.Y(n_11658)
);

INVx2_ASAP7_75t_L g11659 ( 
.A(n_10226),
.Y(n_11659)
);

OA21x2_ASAP7_75t_L g11660 ( 
.A1(n_10291),
.A2(n_10015),
.B(n_10014),
.Y(n_11660)
);

AOI21xp5_ASAP7_75t_L g11661 ( 
.A1(n_10498),
.A2(n_10070),
.B(n_9837),
.Y(n_11661)
);

AND2x4_ASAP7_75t_L g11662 ( 
.A(n_10246),
.B(n_10160),
.Y(n_11662)
);

OAI22xp5_ASAP7_75t_L g11663 ( 
.A1(n_10983),
.A2(n_9800),
.B1(n_9767),
.B2(n_9707),
.Y(n_11663)
);

INVx1_ASAP7_75t_L g11664 ( 
.A(n_10207),
.Y(n_11664)
);

AND2x4_ASAP7_75t_L g11665 ( 
.A(n_10246),
.B(n_10043),
.Y(n_11665)
);

OA22x2_ASAP7_75t_L g11666 ( 
.A1(n_10983),
.A2(n_9178),
.B1(n_9236),
.B2(n_9477),
.Y(n_11666)
);

HB1xp67_ASAP7_75t_L g11667 ( 
.A(n_10476),
.Y(n_11667)
);

INVx2_ASAP7_75t_L g11668 ( 
.A(n_10226),
.Y(n_11668)
);

AND2x4_ASAP7_75t_L g11669 ( 
.A(n_10246),
.B(n_10043),
.Y(n_11669)
);

AND2x2_ASAP7_75t_L g11670 ( 
.A(n_11307),
.B(n_9538),
.Y(n_11670)
);

NAND2xp5_ASAP7_75t_L g11671 ( 
.A(n_10683),
.B(n_9374),
.Y(n_11671)
);

AND2x2_ASAP7_75t_L g11672 ( 
.A(n_10247),
.B(n_11012),
.Y(n_11672)
);

INVx1_ASAP7_75t_L g11673 ( 
.A(n_10207),
.Y(n_11673)
);

INVx2_ASAP7_75t_SL g11674 ( 
.A(n_10423),
.Y(n_11674)
);

HB1xp67_ASAP7_75t_L g11675 ( 
.A(n_10484),
.Y(n_11675)
);

OAI22xp5_ASAP7_75t_L g11676 ( 
.A1(n_10918),
.A2(n_9800),
.B1(n_9707),
.B2(n_9745),
.Y(n_11676)
);

AOI21x1_ASAP7_75t_SL g11677 ( 
.A1(n_10994),
.A2(n_9565),
.B(n_9506),
.Y(n_11677)
);

NAND2x1p5_ASAP7_75t_L g11678 ( 
.A(n_10247),
.B(n_9837),
.Y(n_11678)
);

OA21x2_ASAP7_75t_L g11679 ( 
.A1(n_10252),
.A2(n_10015),
.B(n_10014),
.Y(n_11679)
);

INVx2_ASAP7_75t_L g11680 ( 
.A(n_10226),
.Y(n_11680)
);

AND2x4_ASAP7_75t_L g11681 ( 
.A(n_10246),
.B(n_10043),
.Y(n_11681)
);

AND2x4_ASAP7_75t_L g11682 ( 
.A(n_10246),
.B(n_10043),
.Y(n_11682)
);

AOI221x1_ASAP7_75t_SL g11683 ( 
.A1(n_10289),
.A2(n_10952),
.B1(n_10994),
.B2(n_11259),
.C(n_10618),
.Y(n_11683)
);

INVx2_ASAP7_75t_L g11684 ( 
.A(n_10226),
.Y(n_11684)
);

AND2x2_ASAP7_75t_L g11685 ( 
.A(n_10247),
.B(n_9538),
.Y(n_11685)
);

NAND2xp5_ASAP7_75t_L g11686 ( 
.A(n_10683),
.B(n_10806),
.Y(n_11686)
);

OAI22xp5_ASAP7_75t_L g11687 ( 
.A1(n_10918),
.A2(n_9707),
.B1(n_9745),
.B2(n_9738),
.Y(n_11687)
);

CKINVDCx12_ASAP7_75t_R g11688 ( 
.A(n_10684),
.Y(n_11688)
);

AOI21x1_ASAP7_75t_SL g11689 ( 
.A1(n_11259),
.A2(n_9565),
.B(n_9506),
.Y(n_11689)
);

AOI21x1_ASAP7_75t_SL g11690 ( 
.A1(n_10809),
.A2(n_9157),
.B(n_9150),
.Y(n_11690)
);

INVx2_ASAP7_75t_L g11691 ( 
.A(n_10226),
.Y(n_11691)
);

OAI22xp5_ASAP7_75t_L g11692 ( 
.A1(n_10396),
.A2(n_9745),
.B1(n_9738),
.B2(n_9178),
.Y(n_11692)
);

OAI22xp5_ASAP7_75t_L g11693 ( 
.A1(n_10229),
.A2(n_9738),
.B1(n_9178),
.B2(n_9830),
.Y(n_11693)
);

INVx2_ASAP7_75t_L g11694 ( 
.A(n_10226),
.Y(n_11694)
);

NOR2x1_ASAP7_75t_SL g11695 ( 
.A(n_11081),
.B(n_9296),
.Y(n_11695)
);

OAI22xp5_ASAP7_75t_L g11696 ( 
.A1(n_10229),
.A2(n_9738),
.B1(n_9830),
.B2(n_9099),
.Y(n_11696)
);

AOI21xp5_ASAP7_75t_L g11697 ( 
.A1(n_10400),
.A2(n_10070),
.B(n_9837),
.Y(n_11697)
);

OA21x2_ASAP7_75t_L g11698 ( 
.A1(n_10252),
.A2(n_10015),
.B(n_10014),
.Y(n_11698)
);

AND2x2_ASAP7_75t_L g11699 ( 
.A(n_10247),
.B(n_11012),
.Y(n_11699)
);

NOR2xp67_ASAP7_75t_L g11700 ( 
.A(n_10247),
.B(n_9854),
.Y(n_11700)
);

OR2x2_ASAP7_75t_L g11701 ( 
.A(n_10342),
.B(n_9901),
.Y(n_11701)
);

INVx1_ASAP7_75t_L g11702 ( 
.A(n_10213),
.Y(n_11702)
);

AOI221x1_ASAP7_75t_SL g11703 ( 
.A1(n_10289),
.A2(n_9474),
.B1(n_9469),
.B2(n_9150),
.C(n_9157),
.Y(n_11703)
);

OAI22xp5_ASAP7_75t_L g11704 ( 
.A1(n_10240),
.A2(n_9738),
.B1(n_9830),
.B2(n_9099),
.Y(n_11704)
);

INVx1_ASAP7_75t_L g11705 ( 
.A(n_10213),
.Y(n_11705)
);

INVxp67_ASAP7_75t_SL g11706 ( 
.A(n_10378),
.Y(n_11706)
);

OAI22xp5_ASAP7_75t_L g11707 ( 
.A1(n_10240),
.A2(n_9738),
.B1(n_9099),
.B2(n_9287),
.Y(n_11707)
);

NAND2xp5_ASAP7_75t_L g11708 ( 
.A(n_10806),
.B(n_9384),
.Y(n_11708)
);

HB1xp67_ASAP7_75t_L g11709 ( 
.A(n_10484),
.Y(n_11709)
);

AOI21x1_ASAP7_75t_SL g11710 ( 
.A1(n_10809),
.A2(n_9157),
.B(n_9150),
.Y(n_11710)
);

AND2x2_ASAP7_75t_L g11711 ( 
.A(n_10247),
.B(n_9547),
.Y(n_11711)
);

NAND2xp5_ASAP7_75t_L g11712 ( 
.A(n_10567),
.B(n_9384),
.Y(n_11712)
);

CKINVDCx20_ASAP7_75t_R g11713 ( 
.A(n_10377),
.Y(n_11713)
);

AND2x4_ASAP7_75t_L g11714 ( 
.A(n_10234),
.B(n_10189),
.Y(n_11714)
);

INVx2_ASAP7_75t_L g11715 ( 
.A(n_10226),
.Y(n_11715)
);

HB1xp67_ASAP7_75t_L g11716 ( 
.A(n_10487),
.Y(n_11716)
);

NAND2xp5_ASAP7_75t_L g11717 ( 
.A(n_10567),
.B(n_9384),
.Y(n_11717)
);

NAND2xp5_ASAP7_75t_L g11718 ( 
.A(n_10620),
.B(n_9615),
.Y(n_11718)
);

NOR2xp67_ASAP7_75t_L g11719 ( 
.A(n_10247),
.B(n_9854),
.Y(n_11719)
);

NAND2xp5_ASAP7_75t_L g11720 ( 
.A(n_10620),
.B(n_9615),
.Y(n_11720)
);

AOI21xp5_ASAP7_75t_SL g11721 ( 
.A1(n_10209),
.A2(n_9585),
.B(n_9440),
.Y(n_11721)
);

AND2x2_ASAP7_75t_L g11722 ( 
.A(n_11012),
.B(n_9547),
.Y(n_11722)
);

AOI21xp5_ASAP7_75t_L g11723 ( 
.A1(n_10400),
.A2(n_10070),
.B(n_9177),
.Y(n_11723)
);

O2A1O1Ixp33_ASAP7_75t_L g11724 ( 
.A1(n_10752),
.A2(n_10463),
.B(n_10705),
.C(n_11075),
.Y(n_11724)
);

OR2x2_ASAP7_75t_L g11725 ( 
.A(n_10342),
.B(n_9901),
.Y(n_11725)
);

OAI22xp5_ASAP7_75t_L g11726 ( 
.A1(n_10705),
.A2(n_9738),
.B1(n_9099),
.B2(n_9287),
.Y(n_11726)
);

AO21x2_ASAP7_75t_L g11727 ( 
.A1(n_10392),
.A2(n_9631),
.B(n_10117),
.Y(n_11727)
);

AND2x2_ASAP7_75t_L g11728 ( 
.A(n_11012),
.B(n_9547),
.Y(n_11728)
);

AND2x2_ASAP7_75t_L g11729 ( 
.A(n_11012),
.B(n_9547),
.Y(n_11729)
);

INVx3_ASAP7_75t_SL g11730 ( 
.A(n_10233),
.Y(n_11730)
);

NAND2xp5_ASAP7_75t_L g11731 ( 
.A(n_10558),
.B(n_9615),
.Y(n_11731)
);

AND2x2_ASAP7_75t_L g11732 ( 
.A(n_11012),
.B(n_11556),
.Y(n_11732)
);

OAI22xp5_ASAP7_75t_L g11733 ( 
.A1(n_10909),
.A2(n_9099),
.B1(n_9287),
.B2(n_9025),
.Y(n_11733)
);

INVx2_ASAP7_75t_SL g11734 ( 
.A(n_10423),
.Y(n_11734)
);

OAI22xp5_ASAP7_75t_L g11735 ( 
.A1(n_10909),
.A2(n_10530),
.B1(n_10463),
.B2(n_10325),
.Y(n_11735)
);

INVx1_ASAP7_75t_L g11736 ( 
.A(n_10222),
.Y(n_11736)
);

AND2x4_ASAP7_75t_L g11737 ( 
.A(n_10234),
.B(n_10189),
.Y(n_11737)
);

NAND2xp5_ASAP7_75t_L g11738 ( 
.A(n_10558),
.B(n_9822),
.Y(n_11738)
);

O2A1O1Ixp33_ASAP7_75t_L g11739 ( 
.A1(n_11075),
.A2(n_9177),
.B(n_9036),
.C(n_9631),
.Y(n_11739)
);

INVx1_ASAP7_75t_L g11740 ( 
.A(n_10222),
.Y(n_11740)
);

AOI21xp5_ASAP7_75t_SL g11741 ( 
.A1(n_10209),
.A2(n_9770),
.B(n_9063),
.Y(n_11741)
);

OR2x6_ASAP7_75t_L g11742 ( 
.A(n_11152),
.B(n_9798),
.Y(n_11742)
);

OAI22xp5_ASAP7_75t_L g11743 ( 
.A1(n_10530),
.A2(n_9287),
.B1(n_9025),
.B2(n_9076),
.Y(n_11743)
);

OAI22xp5_ASAP7_75t_L g11744 ( 
.A1(n_10325),
.A2(n_9287),
.B1(n_9076),
.B2(n_10041),
.Y(n_11744)
);

OAI22xp5_ASAP7_75t_L g11745 ( 
.A1(n_10828),
.A2(n_10402),
.B1(n_10647),
.B2(n_10697),
.Y(n_11745)
);

OA21x2_ASAP7_75t_L g11746 ( 
.A1(n_10367),
.A2(n_11484),
.B(n_10392),
.Y(n_11746)
);

INVx1_ASAP7_75t_L g11747 ( 
.A(n_10228),
.Y(n_11747)
);

AOI21x1_ASAP7_75t_SL g11748 ( 
.A1(n_10200),
.A2(n_9599),
.B(n_9607),
.Y(n_11748)
);

INVx2_ASAP7_75t_L g11749 ( 
.A(n_10308),
.Y(n_11749)
);

OR2x2_ASAP7_75t_L g11750 ( 
.A(n_10215),
.B(n_9901),
.Y(n_11750)
);

AOI21xp5_ASAP7_75t_L g11751 ( 
.A1(n_10894),
.A2(n_9036),
.B(n_9220),
.Y(n_11751)
);

AND2x2_ASAP7_75t_L g11752 ( 
.A(n_11012),
.B(n_9547),
.Y(n_11752)
);

HB1xp67_ASAP7_75t_L g11753 ( 
.A(n_10487),
.Y(n_11753)
);

AND2x2_ASAP7_75t_L g11754 ( 
.A(n_11556),
.B(n_9567),
.Y(n_11754)
);

NAND2xp5_ASAP7_75t_L g11755 ( 
.A(n_10413),
.B(n_9822),
.Y(n_11755)
);

OAI22xp5_ASAP7_75t_L g11756 ( 
.A1(n_10828),
.A2(n_9076),
.B1(n_10088),
.B2(n_9612),
.Y(n_11756)
);

A2O1A1Ixp33_ASAP7_75t_L g11757 ( 
.A1(n_10952),
.A2(n_9248),
.B(n_9415),
.C(n_9362),
.Y(n_11757)
);

AND2x2_ASAP7_75t_L g11758 ( 
.A(n_11556),
.B(n_9567),
.Y(n_11758)
);

AOI21xp5_ASAP7_75t_L g11759 ( 
.A1(n_10894),
.A2(n_9220),
.B(n_9362),
.Y(n_11759)
);

INVx1_ASAP7_75t_L g11760 ( 
.A(n_10228),
.Y(n_11760)
);

OR2x2_ASAP7_75t_L g11761 ( 
.A(n_10215),
.B(n_9901),
.Y(n_11761)
);

AOI21xp5_ASAP7_75t_SL g11762 ( 
.A1(n_10684),
.A2(n_9770),
.B(n_9063),
.Y(n_11762)
);

AOI21xp5_ASAP7_75t_SL g11763 ( 
.A1(n_11038),
.A2(n_9770),
.B(n_9063),
.Y(n_11763)
);

INVx1_ASAP7_75t_L g11764 ( 
.A(n_10235),
.Y(n_11764)
);

AOI21x1_ASAP7_75t_SL g11765 ( 
.A1(n_10200),
.A2(n_9617),
.B(n_9607),
.Y(n_11765)
);

OA21x2_ASAP7_75t_L g11766 ( 
.A1(n_10367),
.A2(n_10015),
.B(n_10014),
.Y(n_11766)
);

AOI21x1_ASAP7_75t_SL g11767 ( 
.A1(n_10208),
.A2(n_9617),
.B(n_9607),
.Y(n_11767)
);

OR2x2_ASAP7_75t_L g11768 ( 
.A(n_10309),
.B(n_9901),
.Y(n_11768)
);

AND2x2_ASAP7_75t_L g11769 ( 
.A(n_11556),
.B(n_9567),
.Y(n_11769)
);

NAND2xp5_ASAP7_75t_L g11770 ( 
.A(n_10413),
.B(n_9822),
.Y(n_11770)
);

NAND2xp5_ASAP7_75t_L g11771 ( 
.A(n_10635),
.B(n_9850),
.Y(n_11771)
);

NAND2xp5_ASAP7_75t_L g11772 ( 
.A(n_10635),
.B(n_9850),
.Y(n_11772)
);

INVx1_ASAP7_75t_L g11773 ( 
.A(n_10235),
.Y(n_11773)
);

INVx1_ASAP7_75t_L g11774 ( 
.A(n_10241),
.Y(n_11774)
);

O2A1O1Ixp33_ASAP7_75t_L g11775 ( 
.A1(n_10409),
.A2(n_9631),
.B(n_9469),
.C(n_9248),
.Y(n_11775)
);

AND2x2_ASAP7_75t_L g11776 ( 
.A(n_11556),
.B(n_9567),
.Y(n_11776)
);

INVx1_ASAP7_75t_L g11777 ( 
.A(n_10241),
.Y(n_11777)
);

INVx2_ASAP7_75t_L g11778 ( 
.A(n_10308),
.Y(n_11778)
);

INVx1_ASAP7_75t_L g11779 ( 
.A(n_10250),
.Y(n_11779)
);

O2A1O1Ixp33_ASAP7_75t_L g11780 ( 
.A1(n_10409),
.A2(n_9631),
.B(n_9248),
.C(n_9617),
.Y(n_11780)
);

AND2x4_ASAP7_75t_L g11781 ( 
.A(n_10234),
.B(n_10189),
.Y(n_11781)
);

AND2x2_ASAP7_75t_L g11782 ( 
.A(n_11556),
.B(n_9567),
.Y(n_11782)
);

AND2x2_ASAP7_75t_L g11783 ( 
.A(n_11556),
.B(n_9581),
.Y(n_11783)
);

AND2x2_ASAP7_75t_L g11784 ( 
.A(n_11556),
.B(n_9581),
.Y(n_11784)
);

INVx2_ASAP7_75t_SL g11785 ( 
.A(n_10423),
.Y(n_11785)
);

INVx2_ASAP7_75t_L g11786 ( 
.A(n_10308),
.Y(n_11786)
);

NAND2xp5_ASAP7_75t_L g11787 ( 
.A(n_10309),
.B(n_9850),
.Y(n_11787)
);

AND2x2_ASAP7_75t_L g11788 ( 
.A(n_10678),
.B(n_10911),
.Y(n_11788)
);

INVx1_ASAP7_75t_L g11789 ( 
.A(n_10250),
.Y(n_11789)
);

HB1xp67_ASAP7_75t_L g11790 ( 
.A(n_10493),
.Y(n_11790)
);

OAI22xp5_ASAP7_75t_L g11791 ( 
.A1(n_10402),
.A2(n_10647),
.B1(n_10697),
.B2(n_11177),
.Y(n_11791)
);

OR2x2_ASAP7_75t_L g11792 ( 
.A(n_10313),
.B(n_9901),
.Y(n_11792)
);

AND2x2_ASAP7_75t_L g11793 ( 
.A(n_10678),
.B(n_9581),
.Y(n_11793)
);

INVx3_ASAP7_75t_L g11794 ( 
.A(n_11597),
.Y(n_11794)
);

A2O1A1Ixp33_ASAP7_75t_L g11795 ( 
.A1(n_11046),
.A2(n_9415),
.B(n_9362),
.C(n_9755),
.Y(n_11795)
);

AND2x2_ASAP7_75t_L g11796 ( 
.A(n_10678),
.B(n_9581),
.Y(n_11796)
);

O2A1O1Ixp5_ASAP7_75t_L g11797 ( 
.A1(n_10392),
.A2(n_9263),
.B(n_9416),
.C(n_9409),
.Y(n_11797)
);

OR2x2_ASAP7_75t_L g11798 ( 
.A(n_10313),
.B(n_9901),
.Y(n_11798)
);

CKINVDCx11_ASAP7_75t_R g11799 ( 
.A(n_10263),
.Y(n_11799)
);

AND2x2_ASAP7_75t_L g11800 ( 
.A(n_10911),
.B(n_9581),
.Y(n_11800)
);

INVxp67_ASAP7_75t_L g11801 ( 
.A(n_10448),
.Y(n_11801)
);

BUFx2_ASAP7_75t_L g11802 ( 
.A(n_10736),
.Y(n_11802)
);

AND2x4_ASAP7_75t_L g11803 ( 
.A(n_10234),
.B(n_10160),
.Y(n_11803)
);

AND2x2_ASAP7_75t_L g11804 ( 
.A(n_10911),
.B(n_9175),
.Y(n_11804)
);

OAI22xp5_ASAP7_75t_L g11805 ( 
.A1(n_11177),
.A2(n_10088),
.B1(n_9612),
.B2(n_9610),
.Y(n_11805)
);

AND2x4_ASAP7_75t_L g11806 ( 
.A(n_10239),
.B(n_10160),
.Y(n_11806)
);

INVx2_ASAP7_75t_L g11807 ( 
.A(n_10308),
.Y(n_11807)
);

INVx1_ASAP7_75t_L g11808 ( 
.A(n_10257),
.Y(n_11808)
);

AOI21xp5_ASAP7_75t_L g11809 ( 
.A1(n_11046),
.A2(n_10013),
.B(n_10010),
.Y(n_11809)
);

AND2x4_ASAP7_75t_L g11810 ( 
.A(n_10239),
.B(n_10160),
.Y(n_11810)
);

INVx1_ASAP7_75t_L g11811 ( 
.A(n_10257),
.Y(n_11811)
);

NAND2xp5_ASAP7_75t_L g11812 ( 
.A(n_11088),
.B(n_9729),
.Y(n_11812)
);

A2O1A1Ixp33_ASAP7_75t_L g11813 ( 
.A1(n_10945),
.A2(n_9415),
.B(n_9755),
.C(n_9816),
.Y(n_11813)
);

CKINVDCx12_ASAP7_75t_R g11814 ( 
.A(n_11038),
.Y(n_11814)
);

HB1xp67_ASAP7_75t_L g11815 ( 
.A(n_10493),
.Y(n_11815)
);

AND2x6_ASAP7_75t_L g11816 ( 
.A(n_10239),
.B(n_10063),
.Y(n_11816)
);

INVx2_ASAP7_75t_L g11817 ( 
.A(n_10308),
.Y(n_11817)
);

HB1xp67_ASAP7_75t_SL g11818 ( 
.A(n_10581),
.Y(n_11818)
);

AOI21x1_ASAP7_75t_SL g11819 ( 
.A1(n_10208),
.A2(n_9646),
.B(n_9640),
.Y(n_11819)
);

AND2x2_ASAP7_75t_L g11820 ( 
.A(n_11099),
.B(n_8756),
.Y(n_11820)
);

NAND2xp5_ASAP7_75t_L g11821 ( 
.A(n_11088),
.B(n_9729),
.Y(n_11821)
);

OA21x2_ASAP7_75t_L g11822 ( 
.A1(n_11484),
.A2(n_10015),
.B(n_10014),
.Y(n_11822)
);

INVx2_ASAP7_75t_SL g11823 ( 
.A(n_10423),
.Y(n_11823)
);

AOI21x1_ASAP7_75t_SL g11824 ( 
.A1(n_11318),
.A2(n_9646),
.B(n_9640),
.Y(n_11824)
);

INVx1_ASAP7_75t_SL g11825 ( 
.A(n_10788),
.Y(n_11825)
);

O2A1O1Ixp5_ASAP7_75t_L g11826 ( 
.A1(n_10866),
.A2(n_9263),
.B(n_9416),
.C(n_9409),
.Y(n_11826)
);

AOI21xp5_ASAP7_75t_L g11827 ( 
.A1(n_11051),
.A2(n_10013),
.B(n_10010),
.Y(n_11827)
);

CKINVDCx20_ASAP7_75t_R g11828 ( 
.A(n_10377),
.Y(n_11828)
);

OAI22xp5_ASAP7_75t_L g11829 ( 
.A1(n_11052),
.A2(n_10088),
.B1(n_9612),
.B2(n_9610),
.Y(n_11829)
);

OAI22xp5_ASAP7_75t_L g11830 ( 
.A1(n_11052),
.A2(n_9610),
.B1(n_9626),
.B2(n_9423),
.Y(n_11830)
);

OAI22xp5_ASAP7_75t_L g11831 ( 
.A1(n_11014),
.A2(n_9626),
.B1(n_9085),
.B2(n_9009),
.Y(n_11831)
);

OAI22x1_ASAP7_75t_L g11832 ( 
.A1(n_10366),
.A2(n_9321),
.B1(n_9443),
.B2(n_9406),
.Y(n_11832)
);

OA21x2_ASAP7_75t_L g11833 ( 
.A1(n_10556),
.A2(n_10016),
.B(n_10120),
.Y(n_11833)
);

INVxp67_ASAP7_75t_L g11834 ( 
.A(n_10448),
.Y(n_11834)
);

NAND2xp5_ASAP7_75t_L g11835 ( 
.A(n_11138),
.B(n_9729),
.Y(n_11835)
);

INVx1_ASAP7_75t_L g11836 ( 
.A(n_10258),
.Y(n_11836)
);

OA21x2_ASAP7_75t_L g11837 ( 
.A1(n_10556),
.A2(n_10016),
.B(n_10120),
.Y(n_11837)
);

NAND2xp5_ASAP7_75t_L g11838 ( 
.A(n_11138),
.B(n_11281),
.Y(n_11838)
);

CKINVDCx5p33_ASAP7_75t_R g11839 ( 
.A(n_10369),
.Y(n_11839)
);

AOI211xp5_ASAP7_75t_L g11840 ( 
.A1(n_10690),
.A2(n_9263),
.B(n_9416),
.C(n_9409),
.Y(n_11840)
);

O2A1O1Ixp5_ASAP7_75t_L g11841 ( 
.A1(n_10866),
.A2(n_9140),
.B(n_9413),
.C(n_9259),
.Y(n_11841)
);

AOI21xp5_ASAP7_75t_L g11842 ( 
.A1(n_11051),
.A2(n_10013),
.B(n_10010),
.Y(n_11842)
);

AOI21xp5_ASAP7_75t_SL g11843 ( 
.A1(n_10588),
.A2(n_9770),
.B(n_9063),
.Y(n_11843)
);

A2O1A1Ixp33_ASAP7_75t_L g11844 ( 
.A1(n_10945),
.A2(n_9755),
.B(n_9816),
.C(n_9446),
.Y(n_11844)
);

OAI22xp5_ASAP7_75t_SL g11845 ( 
.A1(n_10465),
.A2(n_9477),
.B1(n_9601),
.B2(n_9507),
.Y(n_11845)
);

AND2x2_ASAP7_75t_L g11846 ( 
.A(n_11099),
.B(n_9018),
.Y(n_11846)
);

AOI21x1_ASAP7_75t_SL g11847 ( 
.A1(n_11318),
.A2(n_9646),
.B(n_9640),
.Y(n_11847)
);

INVx1_ASAP7_75t_L g11848 ( 
.A(n_10258),
.Y(n_11848)
);

AND2x2_ASAP7_75t_L g11849 ( 
.A(n_11099),
.B(n_9018),
.Y(n_11849)
);

OAI22xp5_ASAP7_75t_L g11850 ( 
.A1(n_11014),
.A2(n_9085),
.B1(n_9009),
.B2(n_9030),
.Y(n_11850)
);

AND2x4_ASAP7_75t_L g11851 ( 
.A(n_10239),
.B(n_10189),
.Y(n_11851)
);

INVx1_ASAP7_75t_L g11852 ( 
.A(n_10261),
.Y(n_11852)
);

AOI21xp5_ASAP7_75t_L g11853 ( 
.A1(n_10652),
.A2(n_10013),
.B(n_10010),
.Y(n_11853)
);

INVx1_ASAP7_75t_L g11854 ( 
.A(n_10261),
.Y(n_11854)
);

AOI21xp5_ASAP7_75t_L g11855 ( 
.A1(n_10652),
.A2(n_10013),
.B(n_10010),
.Y(n_11855)
);

HB1xp67_ASAP7_75t_L g11856 ( 
.A(n_10308),
.Y(n_11856)
);

OAI22xp5_ASAP7_75t_L g11857 ( 
.A1(n_11214),
.A2(n_9085),
.B1(n_9009),
.B2(n_9030),
.Y(n_11857)
);

OAI22xp5_ASAP7_75t_L g11858 ( 
.A1(n_11214),
.A2(n_10732),
.B1(n_11199),
.B2(n_10827),
.Y(n_11858)
);

NOR2xp33_ASAP7_75t_L g11859 ( 
.A(n_10465),
.B(n_9367),
.Y(n_11859)
);

OA21x2_ASAP7_75t_L g11860 ( 
.A1(n_10529),
.A2(n_10016),
.B(n_10120),
.Y(n_11860)
);

INVx1_ASAP7_75t_L g11861 ( 
.A(n_10262),
.Y(n_11861)
);

OA21x2_ASAP7_75t_L g11862 ( 
.A1(n_10529),
.A2(n_10559),
.B(n_11343),
.Y(n_11862)
);

NAND2xp5_ASAP7_75t_L g11863 ( 
.A(n_11281),
.B(n_9530),
.Y(n_11863)
);

AND2x2_ASAP7_75t_L g11864 ( 
.A(n_11179),
.B(n_9018),
.Y(n_11864)
);

O2A1O1Ixp5_ASAP7_75t_L g11865 ( 
.A1(n_10588),
.A2(n_10361),
.B(n_10363),
.C(n_10566),
.Y(n_11865)
);

INVx2_ASAP7_75t_L g11866 ( 
.A(n_10308),
.Y(n_11866)
);

OA21x2_ASAP7_75t_L g11867 ( 
.A1(n_10559),
.A2(n_10016),
.B(n_10120),
.Y(n_11867)
);

OA22x2_ASAP7_75t_L g11868 ( 
.A1(n_10275),
.A2(n_10692),
.B1(n_10566),
.B2(n_10259),
.Y(n_11868)
);

OR2x2_ASAP7_75t_L g11869 ( 
.A(n_10338),
.B(n_9901),
.Y(n_11869)
);

NAND2xp5_ASAP7_75t_L g11870 ( 
.A(n_10253),
.B(n_9534),
.Y(n_11870)
);

OA22x2_ASAP7_75t_L g11871 ( 
.A1(n_10275),
.A2(n_9236),
.B1(n_9477),
.B2(n_9401),
.Y(n_11871)
);

HB1xp67_ASAP7_75t_L g11872 ( 
.A(n_10308),
.Y(n_11872)
);

NAND2xp5_ASAP7_75t_L g11873 ( 
.A(n_10253),
.B(n_9534),
.Y(n_11873)
);

NAND2xp5_ASAP7_75t_L g11874 ( 
.A(n_10277),
.B(n_9534),
.Y(n_11874)
);

AND2x2_ASAP7_75t_L g11875 ( 
.A(n_11179),
.B(n_9018),
.Y(n_11875)
);

O2A1O1Ixp5_ASAP7_75t_L g11876 ( 
.A1(n_10361),
.A2(n_9140),
.B(n_9413),
.C(n_9259),
.Y(n_11876)
);

BUFx8_ASAP7_75t_SL g11877 ( 
.A(n_10736),
.Y(n_11877)
);

OR2x2_ASAP7_75t_L g11878 ( 
.A(n_10338),
.B(n_9901),
.Y(n_11878)
);

AOI21xp5_ASAP7_75t_SL g11879 ( 
.A1(n_10739),
.A2(n_9059),
.B(n_9401),
.Y(n_11879)
);

OR2x2_ASAP7_75t_L g11880 ( 
.A(n_10783),
.B(n_9901),
.Y(n_11880)
);

AOI21xp5_ASAP7_75t_L g11881 ( 
.A1(n_10633),
.A2(n_10013),
.B(n_10010),
.Y(n_11881)
);

AND2x2_ASAP7_75t_L g11882 ( 
.A(n_11179),
.B(n_9018),
.Y(n_11882)
);

O2A1O1Ixp33_ASAP7_75t_L g11883 ( 
.A1(n_10453),
.A2(n_10117),
.B(n_9246),
.C(n_9140),
.Y(n_11883)
);

AND2x2_ASAP7_75t_L g11884 ( 
.A(n_11193),
.B(n_9104),
.Y(n_11884)
);

OAI22xp5_ASAP7_75t_L g11885 ( 
.A1(n_10732),
.A2(n_9030),
.B1(n_9515),
.B2(n_9106),
.Y(n_11885)
);

AND2x2_ASAP7_75t_L g11886 ( 
.A(n_11193),
.B(n_9104),
.Y(n_11886)
);

CKINVDCx6p67_ASAP7_75t_R g11887 ( 
.A(n_10454),
.Y(n_11887)
);

INVx1_ASAP7_75t_L g11888 ( 
.A(n_10262),
.Y(n_11888)
);

HB1xp67_ASAP7_75t_L g11889 ( 
.A(n_10328),
.Y(n_11889)
);

HB1xp67_ASAP7_75t_L g11890 ( 
.A(n_10328),
.Y(n_11890)
);

NOR2xp33_ASAP7_75t_L g11891 ( 
.A(n_10465),
.B(n_9509),
.Y(n_11891)
);

AOI21x1_ASAP7_75t_SL g11892 ( 
.A1(n_11319),
.A2(n_11185),
.B(n_11136),
.Y(n_11892)
);

A2O1A1Ixp33_ASAP7_75t_L g11893 ( 
.A1(n_10502),
.A2(n_10544),
.B(n_10739),
.C(n_10720),
.Y(n_11893)
);

AND2x2_ASAP7_75t_L g11894 ( 
.A(n_11193),
.B(n_9104),
.Y(n_11894)
);

OR2x2_ASAP7_75t_L g11895 ( 
.A(n_10783),
.B(n_9901),
.Y(n_11895)
);

AND2x2_ASAP7_75t_L g11896 ( 
.A(n_11195),
.B(n_9104),
.Y(n_11896)
);

INVx2_ASAP7_75t_L g11897 ( 
.A(n_10328),
.Y(n_11897)
);

AOI21xp5_ASAP7_75t_L g11898 ( 
.A1(n_10633),
.A2(n_10013),
.B(n_10010),
.Y(n_11898)
);

NAND2xp5_ASAP7_75t_L g11899 ( 
.A(n_10277),
.B(n_9536),
.Y(n_11899)
);

INVx1_ASAP7_75t_L g11900 ( 
.A(n_10270),
.Y(n_11900)
);

OAI22xp5_ASAP7_75t_L g11901 ( 
.A1(n_11199),
.A2(n_9515),
.B1(n_9106),
.B2(n_9657),
.Y(n_11901)
);

INVx2_ASAP7_75t_L g11902 ( 
.A(n_10328),
.Y(n_11902)
);

AND2x2_ASAP7_75t_L g11903 ( 
.A(n_11195),
.B(n_9104),
.Y(n_11903)
);

OA21x2_ASAP7_75t_L g11904 ( 
.A1(n_11343),
.A2(n_10016),
.B(n_10120),
.Y(n_11904)
);

NAND2xp5_ASAP7_75t_L g11905 ( 
.A(n_10284),
.B(n_9536),
.Y(n_11905)
);

INVxp67_ASAP7_75t_L g11906 ( 
.A(n_10581),
.Y(n_11906)
);

OR2x2_ASAP7_75t_L g11907 ( 
.A(n_10797),
.B(n_8335),
.Y(n_11907)
);

NAND2xp5_ASAP7_75t_L g11908 ( 
.A(n_10284),
.B(n_9536),
.Y(n_11908)
);

AND2x2_ASAP7_75t_L g11909 ( 
.A(n_11195),
.B(n_9105),
.Y(n_11909)
);

OAI22xp5_ASAP7_75t_L g11910 ( 
.A1(n_10827),
.A2(n_9515),
.B1(n_9106),
.B2(n_9657),
.Y(n_11910)
);

AOI21x1_ASAP7_75t_SL g11911 ( 
.A1(n_11319),
.A2(n_9192),
.B(n_9191),
.Y(n_11911)
);

O2A1O1Ixp33_ASAP7_75t_L g11912 ( 
.A1(n_10453),
.A2(n_10117),
.B(n_9246),
.C(n_9902),
.Y(n_11912)
);

INVx2_ASAP7_75t_L g11913 ( 
.A(n_10328),
.Y(n_11913)
);

OR2x2_ASAP7_75t_L g11914 ( 
.A(n_10797),
.B(n_8335),
.Y(n_11914)
);

AND2x2_ASAP7_75t_L g11915 ( 
.A(n_11218),
.B(n_9105),
.Y(n_11915)
);

INVx1_ASAP7_75t_L g11916 ( 
.A(n_10270),
.Y(n_11916)
);

OAI22xp5_ASAP7_75t_L g11917 ( 
.A1(n_10346),
.A2(n_9515),
.B1(n_9657),
.B2(n_9127),
.Y(n_11917)
);

AOI21x1_ASAP7_75t_SL g11918 ( 
.A1(n_11136),
.A2(n_11185),
.B(n_10360),
.Y(n_11918)
);

AND2x2_ASAP7_75t_L g11919 ( 
.A(n_11218),
.B(n_9105),
.Y(n_11919)
);

NAND2xp5_ASAP7_75t_L g11920 ( 
.A(n_10552),
.B(n_9545),
.Y(n_11920)
);

O2A1O1Ixp33_ASAP7_75t_L g11921 ( 
.A1(n_10962),
.A2(n_10117),
.B(n_9246),
.C(n_9902),
.Y(n_11921)
);

NAND2xp5_ASAP7_75t_L g11922 ( 
.A(n_10552),
.B(n_9545),
.Y(n_11922)
);

O2A1O1Ixp33_ASAP7_75t_L g11923 ( 
.A1(n_10962),
.A2(n_10117),
.B(n_9902),
.C(n_9957),
.Y(n_11923)
);

O2A1O1Ixp5_ASAP7_75t_L g11924 ( 
.A1(n_10361),
.A2(n_9413),
.B(n_9259),
.C(n_9250),
.Y(n_11924)
);

AND2x4_ASAP7_75t_L g11925 ( 
.A(n_10299),
.B(n_9869),
.Y(n_11925)
);

INVx2_ASAP7_75t_L g11926 ( 
.A(n_10328),
.Y(n_11926)
);

OA21x2_ASAP7_75t_L g11927 ( 
.A1(n_11480),
.A2(n_10001),
.B(n_10000),
.Y(n_11927)
);

AND2x2_ASAP7_75t_L g11928 ( 
.A(n_11218),
.B(n_9105),
.Y(n_11928)
);

AOI21xp5_ASAP7_75t_SL g11929 ( 
.A1(n_11170),
.A2(n_9059),
.B(n_9507),
.Y(n_11929)
);

OAI22xp5_ASAP7_75t_L g11930 ( 
.A1(n_10346),
.A2(n_9127),
.B1(n_9793),
.B2(n_9555),
.Y(n_11930)
);

NAND2xp5_ASAP7_75t_L g11931 ( 
.A(n_10692),
.B(n_9545),
.Y(n_11931)
);

OAI22xp5_ASAP7_75t_L g11932 ( 
.A1(n_11388),
.A2(n_9127),
.B1(n_9793),
.B2(n_9555),
.Y(n_11932)
);

CKINVDCx5p33_ASAP7_75t_R g11933 ( 
.A(n_10454),
.Y(n_11933)
);

OR2x2_ASAP7_75t_L g11934 ( 
.A(n_10841),
.B(n_8335),
.Y(n_11934)
);

NAND2xp5_ASAP7_75t_L g11935 ( 
.A(n_10382),
.B(n_9753),
.Y(n_11935)
);

AOI21x1_ASAP7_75t_SL g11936 ( 
.A1(n_10360),
.A2(n_9192),
.B(n_9191),
.Y(n_11936)
);

NAND2xp5_ASAP7_75t_L g11937 ( 
.A(n_10382),
.B(n_9753),
.Y(n_11937)
);

NAND2xp5_ASAP7_75t_L g11938 ( 
.A(n_10292),
.B(n_9753),
.Y(n_11938)
);

AOI21xp5_ASAP7_75t_L g11939 ( 
.A1(n_10490),
.A2(n_10690),
.B(n_10763),
.Y(n_11939)
);

INVx1_ASAP7_75t_L g11940 ( 
.A(n_10274),
.Y(n_11940)
);

AND2x2_ASAP7_75t_L g11941 ( 
.A(n_11338),
.B(n_9105),
.Y(n_11941)
);

INVx1_ASAP7_75t_L g11942 ( 
.A(n_10274),
.Y(n_11942)
);

NAND2xp5_ASAP7_75t_L g11943 ( 
.A(n_10292),
.B(n_9758),
.Y(n_11943)
);

AOI221xp5_ASAP7_75t_L g11944 ( 
.A1(n_10618),
.A2(n_9192),
.B1(n_9279),
.B2(n_9218),
.C(n_9191),
.Y(n_11944)
);

INVx1_ASAP7_75t_L g11945 ( 
.A(n_10301),
.Y(n_11945)
);

AOI221xp5_ASAP7_75t_L g11946 ( 
.A1(n_10269),
.A2(n_9280),
.B1(n_9291),
.B2(n_9279),
.C(n_9218),
.Y(n_11946)
);

O2A1O1Ixp33_ASAP7_75t_L g11947 ( 
.A1(n_10489),
.A2(n_10117),
.B(n_9902),
.C(n_9957),
.Y(n_11947)
);

OA21x2_ASAP7_75t_L g11948 ( 
.A1(n_11480),
.A2(n_10001),
.B(n_10000),
.Y(n_11948)
);

AOI21xp5_ASAP7_75t_L g11949 ( 
.A1(n_10490),
.A2(n_10013),
.B(n_10010),
.Y(n_11949)
);

AOI21xp5_ASAP7_75t_L g11950 ( 
.A1(n_10763),
.A2(n_9953),
.B(n_9446),
.Y(n_11950)
);

NAND2xp5_ASAP7_75t_L g11951 ( 
.A(n_10841),
.B(n_9758),
.Y(n_11951)
);

BUFx2_ASAP7_75t_L g11952 ( 
.A(n_10736),
.Y(n_11952)
);

AND2x2_ASAP7_75t_L g11953 ( 
.A(n_11338),
.B(n_9728),
.Y(n_11953)
);

BUFx3_ASAP7_75t_L g11954 ( 
.A(n_10379),
.Y(n_11954)
);

OR2x6_ASAP7_75t_L g11955 ( 
.A(n_11280),
.B(n_9798),
.Y(n_11955)
);

BUFx2_ASAP7_75t_L g11956 ( 
.A(n_10877),
.Y(n_11956)
);

NAND2xp5_ASAP7_75t_L g11957 ( 
.A(n_10845),
.B(n_9758),
.Y(n_11957)
);

NAND2xp5_ASAP7_75t_L g11958 ( 
.A(n_10845),
.B(n_9761),
.Y(n_11958)
);

INVx3_ASAP7_75t_SL g11959 ( 
.A(n_10233),
.Y(n_11959)
);

INVx2_ASAP7_75t_L g11960 ( 
.A(n_10328),
.Y(n_11960)
);

O2A1O1Ixp5_ASAP7_75t_L g11961 ( 
.A1(n_10363),
.A2(n_9250),
.B(n_9253),
.C(n_9334),
.Y(n_11961)
);

AND2x2_ASAP7_75t_L g11962 ( 
.A(n_11338),
.B(n_9728),
.Y(n_11962)
);

HB1xp67_ASAP7_75t_L g11963 ( 
.A(n_10328),
.Y(n_11963)
);

AOI21xp5_ASAP7_75t_L g11964 ( 
.A1(n_10658),
.A2(n_10502),
.B(n_10664),
.Y(n_11964)
);

OR2x2_ASAP7_75t_L g11965 ( 
.A(n_10851),
.B(n_8434),
.Y(n_11965)
);

INVx1_ASAP7_75t_L g11966 ( 
.A(n_10301),
.Y(n_11966)
);

INVx3_ASAP7_75t_L g11967 ( 
.A(n_11597),
.Y(n_11967)
);

OAI22xp5_ASAP7_75t_L g11968 ( 
.A1(n_11388),
.A2(n_9555),
.B1(n_9793),
.B2(n_9242),
.Y(n_11968)
);

AOI211xp5_ASAP7_75t_L g11969 ( 
.A1(n_10996),
.A2(n_9344),
.B(n_9334),
.C(n_9546),
.Y(n_11969)
);

OAI22xp5_ASAP7_75t_L g11970 ( 
.A1(n_10627),
.A2(n_9242),
.B1(n_9260),
.B2(n_9082),
.Y(n_11970)
);

OAI22xp5_ASAP7_75t_L g11971 ( 
.A1(n_10627),
.A2(n_9242),
.B1(n_9260),
.B2(n_9082),
.Y(n_11971)
);

AND2x2_ASAP7_75t_L g11972 ( 
.A(n_11384),
.B(n_9728),
.Y(n_11972)
);

AND2x2_ASAP7_75t_L g11973 ( 
.A(n_11384),
.B(n_11494),
.Y(n_11973)
);

NAND2xp5_ASAP7_75t_L g11974 ( 
.A(n_10611),
.B(n_9761),
.Y(n_11974)
);

BUFx3_ASAP7_75t_L g11975 ( 
.A(n_10379),
.Y(n_11975)
);

OA22x2_ASAP7_75t_L g11976 ( 
.A1(n_10275),
.A2(n_9601),
.B1(n_9507),
.B2(n_9814),
.Y(n_11976)
);

O2A1O1Ixp33_ASAP7_75t_L g11977 ( 
.A1(n_10489),
.A2(n_10117),
.B(n_9902),
.C(n_9057),
.Y(n_11977)
);

CKINVDCx5p33_ASAP7_75t_R g11978 ( 
.A(n_10788),
.Y(n_11978)
);

AND2x2_ASAP7_75t_L g11979 ( 
.A(n_11384),
.B(n_9728),
.Y(n_11979)
);

OR2x6_ASAP7_75t_L g11980 ( 
.A(n_11280),
.B(n_9798),
.Y(n_11980)
);

CKINVDCx6p67_ASAP7_75t_R g11981 ( 
.A(n_10465),
.Y(n_11981)
);

AND2x2_ASAP7_75t_L g11982 ( 
.A(n_11494),
.B(n_11507),
.Y(n_11982)
);

INVx2_ASAP7_75t_L g11983 ( 
.A(n_10378),
.Y(n_11983)
);

OR2x2_ASAP7_75t_L g11984 ( 
.A(n_10851),
.B(n_8434),
.Y(n_11984)
);

OA21x2_ASAP7_75t_L g11985 ( 
.A1(n_10768),
.A2(n_10001),
.B(n_10000),
.Y(n_11985)
);

CKINVDCx6p67_ASAP7_75t_R g11986 ( 
.A(n_10233),
.Y(n_11986)
);

OR2x2_ASAP7_75t_L g11987 ( 
.A(n_10885),
.B(n_10920),
.Y(n_11987)
);

AND2x2_ASAP7_75t_L g11988 ( 
.A(n_11494),
.B(n_9728),
.Y(n_11988)
);

AOI21xp5_ASAP7_75t_SL g11989 ( 
.A1(n_11170),
.A2(n_9059),
.B(n_9601),
.Y(n_11989)
);

HB1xp67_ASAP7_75t_L g11990 ( 
.A(n_10315),
.Y(n_11990)
);

AND2x4_ASAP7_75t_L g11991 ( 
.A(n_10299),
.B(n_9381),
.Y(n_11991)
);

INVx1_ASAP7_75t_L g11992 ( 
.A(n_10305),
.Y(n_11992)
);

AND2x2_ASAP7_75t_L g11993 ( 
.A(n_11507),
.B(n_9740),
.Y(n_11993)
);

OAI22xp5_ASAP7_75t_L g11994 ( 
.A1(n_10216),
.A2(n_9260),
.B1(n_9082),
.B2(n_9094),
.Y(n_11994)
);

AND2x2_ASAP7_75t_L g11995 ( 
.A(n_11507),
.B(n_11212),
.Y(n_11995)
);

INVx2_ASAP7_75t_L g11996 ( 
.A(n_10378),
.Y(n_11996)
);

INVx1_ASAP7_75t_L g11997 ( 
.A(n_10305),
.Y(n_11997)
);

OR2x2_ASAP7_75t_L g11998 ( 
.A(n_10885),
.B(n_8434),
.Y(n_11998)
);

NAND2xp5_ASAP7_75t_L g11999 ( 
.A(n_10611),
.B(n_9761),
.Y(n_11999)
);

HB1xp67_ASAP7_75t_L g12000 ( 
.A(n_10315),
.Y(n_12000)
);

AND2x2_ASAP7_75t_L g12001 ( 
.A(n_11212),
.B(n_9740),
.Y(n_12001)
);

INVx3_ASAP7_75t_L g12002 ( 
.A(n_11597),
.Y(n_12002)
);

INVx2_ASAP7_75t_L g12003 ( 
.A(n_10378),
.Y(n_12003)
);

OR2x2_ASAP7_75t_L g12004 ( 
.A(n_10920),
.B(n_8823),
.Y(n_12004)
);

BUFx2_ASAP7_75t_L g12005 ( 
.A(n_10877),
.Y(n_12005)
);

NAND2xp33_ASAP7_75t_SL g12006 ( 
.A(n_10331),
.B(n_9668),
.Y(n_12006)
);

BUFx2_ASAP7_75t_L g12007 ( 
.A(n_10877),
.Y(n_12007)
);

INVx3_ASAP7_75t_L g12008 ( 
.A(n_11597),
.Y(n_12008)
);

NAND2xp5_ASAP7_75t_L g12009 ( 
.A(n_11323),
.B(n_8100),
.Y(n_12009)
);

NAND2xp5_ASAP7_75t_L g12010 ( 
.A(n_11323),
.B(n_8104),
.Y(n_12010)
);

HB1xp67_ASAP7_75t_L g12011 ( 
.A(n_10315),
.Y(n_12011)
);

HB1xp67_ASAP7_75t_L g12012 ( 
.A(n_10315),
.Y(n_12012)
);

BUFx3_ASAP7_75t_L g12013 ( 
.A(n_10423),
.Y(n_12013)
);

INVx2_ASAP7_75t_L g12014 ( 
.A(n_10378),
.Y(n_12014)
);

OA21x2_ASAP7_75t_L g12015 ( 
.A1(n_10768),
.A2(n_10001),
.B(n_10000),
.Y(n_12015)
);

AOI21x1_ASAP7_75t_SL g12016 ( 
.A1(n_11001),
.A2(n_9279),
.B(n_9218),
.Y(n_12016)
);

OAI22xp5_ASAP7_75t_L g12017 ( 
.A1(n_10216),
.A2(n_9082),
.B1(n_9495),
.B2(n_9094),
.Y(n_12017)
);

AND2x2_ASAP7_75t_L g12018 ( 
.A(n_11212),
.B(n_11523),
.Y(n_12018)
);

NAND2xp5_ASAP7_75t_L g12019 ( 
.A(n_10921),
.B(n_8104),
.Y(n_12019)
);

AOI21x1_ASAP7_75t_SL g12020 ( 
.A1(n_11001),
.A2(n_9291),
.B(n_9280),
.Y(n_12020)
);

NAND2xp5_ASAP7_75t_L g12021 ( 
.A(n_10921),
.B(n_8176),
.Y(n_12021)
);

HB1xp67_ASAP7_75t_L g12022 ( 
.A(n_10315),
.Y(n_12022)
);

INVx1_ASAP7_75t_L g12023 ( 
.A(n_10312),
.Y(n_12023)
);

INVx2_ASAP7_75t_L g12024 ( 
.A(n_10378),
.Y(n_12024)
);

AND2x2_ASAP7_75t_L g12025 ( 
.A(n_11212),
.B(n_9740),
.Y(n_12025)
);

AOI221x1_ASAP7_75t_SL g12026 ( 
.A1(n_10269),
.A2(n_9180),
.B1(n_9139),
.B2(n_9459),
.C(n_9457),
.Y(n_12026)
);

INVx1_ASAP7_75t_L g12027 ( 
.A(n_10312),
.Y(n_12027)
);

AND2x4_ASAP7_75t_L g12028 ( 
.A(n_10299),
.B(n_9381),
.Y(n_12028)
);

OAI22xp5_ASAP7_75t_SL g12029 ( 
.A1(n_10638),
.A2(n_10017),
.B1(n_9884),
.B2(n_9765),
.Y(n_12029)
);

OR2x2_ASAP7_75t_L g12030 ( 
.A(n_10368),
.B(n_8823),
.Y(n_12030)
);

NAND2xp5_ASAP7_75t_L g12031 ( 
.A(n_10943),
.B(n_8176),
.Y(n_12031)
);

OAI22xp5_ASAP7_75t_L g12032 ( 
.A1(n_10251),
.A2(n_9082),
.B1(n_9495),
.B2(n_9094),
.Y(n_12032)
);

AND2x2_ASAP7_75t_L g12033 ( 
.A(n_11212),
.B(n_9740),
.Y(n_12033)
);

AOI21xp5_ASAP7_75t_SL g12034 ( 
.A1(n_10959),
.A2(n_9059),
.B(n_9814),
.Y(n_12034)
);

AOI21xp5_ASAP7_75t_L g12035 ( 
.A1(n_10658),
.A2(n_9953),
.B(n_9446),
.Y(n_12035)
);

INVx1_ASAP7_75t_L g12036 ( 
.A(n_10317),
.Y(n_12036)
);

O2A1O1Ixp5_ASAP7_75t_L g12037 ( 
.A1(n_10363),
.A2(n_9250),
.B(n_9253),
.C(n_9334),
.Y(n_12037)
);

INVx2_ASAP7_75t_L g12038 ( 
.A(n_10378),
.Y(n_12038)
);

INVx1_ASAP7_75t_L g12039 ( 
.A(n_10317),
.Y(n_12039)
);

INVxp67_ASAP7_75t_L g12040 ( 
.A(n_10919),
.Y(n_12040)
);

NAND2x1p5_ASAP7_75t_L g12041 ( 
.A(n_11226),
.B(n_9587),
.Y(n_12041)
);

BUFx3_ASAP7_75t_L g12042 ( 
.A(n_10586),
.Y(n_12042)
);

NOR2x1_ASAP7_75t_SL g12043 ( 
.A(n_11081),
.B(n_9296),
.Y(n_12043)
);

AND2x2_ASAP7_75t_L g12044 ( 
.A(n_11212),
.B(n_9740),
.Y(n_12044)
);

AOI21xp5_ASAP7_75t_SL g12045 ( 
.A1(n_10959),
.A2(n_9933),
.B(n_9814),
.Y(n_12045)
);

INVx1_ASAP7_75t_L g12046 ( 
.A(n_10321),
.Y(n_12046)
);

AOI21xp5_ASAP7_75t_SL g12047 ( 
.A1(n_10467),
.A2(n_10090),
.B(n_9933),
.Y(n_12047)
);

NAND2xp5_ASAP7_75t_L g12048 ( 
.A(n_10943),
.B(n_8179),
.Y(n_12048)
);

AND2x2_ASAP7_75t_L g12049 ( 
.A(n_11212),
.B(n_9746),
.Y(n_12049)
);

OAI22xp5_ASAP7_75t_L g12050 ( 
.A1(n_10251),
.A2(n_9082),
.B1(n_9495),
.B2(n_9094),
.Y(n_12050)
);

NAND2xp5_ASAP7_75t_L g12051 ( 
.A(n_10949),
.B(n_8179),
.Y(n_12051)
);

O2A1O1Ixp33_ASAP7_75t_L g12052 ( 
.A1(n_10491),
.A2(n_10117),
.B(n_9902),
.C(n_9057),
.Y(n_12052)
);

OR2x2_ASAP7_75t_L g12053 ( 
.A(n_10368),
.B(n_8177),
.Y(n_12053)
);

AOI21x1_ASAP7_75t_SL g12054 ( 
.A1(n_11011),
.A2(n_9291),
.B(n_9280),
.Y(n_12054)
);

BUFx3_ASAP7_75t_L g12055 ( 
.A(n_10586),
.Y(n_12055)
);

AOI31xp33_ASAP7_75t_L g12056 ( 
.A1(n_10467),
.A2(n_10090),
.A3(n_9933),
.B(n_9353),
.Y(n_12056)
);

INVx2_ASAP7_75t_L g12057 ( 
.A(n_10378),
.Y(n_12057)
);

INVx1_ASAP7_75t_L g12058 ( 
.A(n_10321),
.Y(n_12058)
);

NAND2xp5_ASAP7_75t_L g12059 ( 
.A(n_10949),
.B(n_8189),
.Y(n_12059)
);

OR2x2_ASAP7_75t_L g12060 ( 
.A(n_10386),
.B(n_8177),
.Y(n_12060)
);

INVx6_ASAP7_75t_L g12061 ( 
.A(n_10271),
.Y(n_12061)
);

OAI22xp5_ASAP7_75t_L g12062 ( 
.A1(n_10410),
.A2(n_9082),
.B1(n_9495),
.B2(n_9094),
.Y(n_12062)
);

AOI221x1_ASAP7_75t_SL g12063 ( 
.A1(n_10939),
.A2(n_10765),
.B1(n_11243),
.B2(n_10901),
.C(n_11011),
.Y(n_12063)
);

INVxp67_ASAP7_75t_L g12064 ( 
.A(n_10919),
.Y(n_12064)
);

INVx3_ASAP7_75t_L g12065 ( 
.A(n_11597),
.Y(n_12065)
);

AND2x2_ASAP7_75t_L g12066 ( 
.A(n_11523),
.B(n_10365),
.Y(n_12066)
);

A2O1A1Ixp33_ASAP7_75t_L g12067 ( 
.A1(n_10544),
.A2(n_9619),
.B(n_9811),
.C(n_9344),
.Y(n_12067)
);

O2A1O1Ixp5_ASAP7_75t_L g12068 ( 
.A1(n_11037),
.A2(n_9253),
.B(n_9344),
.C(n_9057),
.Y(n_12068)
);

INVx1_ASAP7_75t_L g12069 ( 
.A(n_10330),
.Y(n_12069)
);

AND2x2_ASAP7_75t_L g12070 ( 
.A(n_11523),
.B(n_9746),
.Y(n_12070)
);

HB1xp67_ASAP7_75t_L g12071 ( 
.A(n_10315),
.Y(n_12071)
);

NAND2xp5_ASAP7_75t_L g12072 ( 
.A(n_10950),
.B(n_8189),
.Y(n_12072)
);

AND2x4_ASAP7_75t_L g12073 ( 
.A(n_10299),
.B(n_9381),
.Y(n_12073)
);

O2A1O1Ixp5_ASAP7_75t_L g12074 ( 
.A1(n_11037),
.A2(n_10996),
.B(n_11058),
.C(n_11031),
.Y(n_12074)
);

AND2x2_ASAP7_75t_L g12075 ( 
.A(n_11523),
.B(n_9746),
.Y(n_12075)
);

INVx2_ASAP7_75t_SL g12076 ( 
.A(n_11431),
.Y(n_12076)
);

OA21x2_ASAP7_75t_L g12077 ( 
.A1(n_10561),
.A2(n_10001),
.B(n_10000),
.Y(n_12077)
);

BUFx2_ASAP7_75t_R g12078 ( 
.A(n_11308),
.Y(n_12078)
);

AND2x2_ASAP7_75t_L g12079 ( 
.A(n_11523),
.B(n_9746),
.Y(n_12079)
);

INVx1_ASAP7_75t_L g12080 ( 
.A(n_10330),
.Y(n_12080)
);

INVx1_ASAP7_75t_L g12081 ( 
.A(n_10352),
.Y(n_12081)
);

AOI21x1_ASAP7_75t_SL g12082 ( 
.A1(n_11017),
.A2(n_9437),
.B(n_9331),
.Y(n_12082)
);

AOI221x1_ASAP7_75t_SL g12083 ( 
.A1(n_10939),
.A2(n_9139),
.B1(n_9180),
.B2(n_9459),
.C(n_9457),
.Y(n_12083)
);

AND2x4_ASAP7_75t_L g12084 ( 
.A(n_10393),
.B(n_9381),
.Y(n_12084)
);

BUFx2_ASAP7_75t_L g12085 ( 
.A(n_10638),
.Y(n_12085)
);

O2A1O1Ixp5_ASAP7_75t_L g12086 ( 
.A1(n_11037),
.A2(n_9570),
.B(n_9546),
.C(n_9501),
.Y(n_12086)
);

OA21x2_ASAP7_75t_L g12087 ( 
.A1(n_10561),
.A2(n_8986),
.B(n_8985),
.Y(n_12087)
);

CKINVDCx5p33_ASAP7_75t_R g12088 ( 
.A(n_11073),
.Y(n_12088)
);

AOI21xp5_ASAP7_75t_L g12089 ( 
.A1(n_10664),
.A2(n_9953),
.B(n_9074),
.Y(n_12089)
);

NAND2xp5_ASAP7_75t_L g12090 ( 
.A(n_10950),
.B(n_8214),
.Y(n_12090)
);

OAI22xp5_ASAP7_75t_L g12091 ( 
.A1(n_10410),
.A2(n_9082),
.B1(n_9495),
.B2(n_9094),
.Y(n_12091)
);

HB1xp67_ASAP7_75t_L g12092 ( 
.A(n_10796),
.Y(n_12092)
);

OA21x2_ASAP7_75t_L g12093 ( 
.A1(n_10343),
.A2(n_8986),
.B(n_8985),
.Y(n_12093)
);

NAND2xp5_ASAP7_75t_L g12094 ( 
.A(n_10977),
.B(n_8214),
.Y(n_12094)
);

AOI21xp5_ASAP7_75t_SL g12095 ( 
.A1(n_10648),
.A2(n_10090),
.B(n_10140),
.Y(n_12095)
);

AND2x4_ASAP7_75t_L g12096 ( 
.A(n_10393),
.B(n_9381),
.Y(n_12096)
);

HB1xp67_ASAP7_75t_L g12097 ( 
.A(n_10796),
.Y(n_12097)
);

AOI21xp5_ASAP7_75t_L g12098 ( 
.A1(n_10491),
.A2(n_9953),
.B(n_9074),
.Y(n_12098)
);

CKINVDCx12_ASAP7_75t_R g12099 ( 
.A(n_11487),
.Y(n_12099)
);

AOI21xp5_ASAP7_75t_SL g12100 ( 
.A1(n_10648),
.A2(n_10162),
.B(n_10140),
.Y(n_12100)
);

OA22x2_ASAP7_75t_L g12101 ( 
.A1(n_10259),
.A2(n_9368),
.B1(n_9347),
.B2(n_9353),
.Y(n_12101)
);

OR2x2_ASAP7_75t_L g12102 ( 
.A(n_10386),
.B(n_8177),
.Y(n_12102)
);

CKINVDCx20_ASAP7_75t_R g12103 ( 
.A(n_10445),
.Y(n_12103)
);

AOI21xp5_ASAP7_75t_SL g12104 ( 
.A1(n_10564),
.A2(n_10162),
.B(n_10140),
.Y(n_12104)
);

INVx1_ASAP7_75t_L g12105 ( 
.A(n_10352),
.Y(n_12105)
);

INVx2_ASAP7_75t_L g12106 ( 
.A(n_10458),
.Y(n_12106)
);

AND2x4_ASAP7_75t_L g12107 ( 
.A(n_10393),
.B(n_9381),
.Y(n_12107)
);

O2A1O1Ixp5_ASAP7_75t_L g12108 ( 
.A1(n_11031),
.A2(n_9570),
.B(n_9546),
.C(n_9501),
.Y(n_12108)
);

O2A1O1Ixp5_ASAP7_75t_L g12109 ( 
.A1(n_11058),
.A2(n_9570),
.B(n_9501),
.C(n_9769),
.Y(n_12109)
);

OA21x2_ASAP7_75t_L g12110 ( 
.A1(n_10343),
.A2(n_8986),
.B(n_8985),
.Y(n_12110)
);

O2A1O1Ixp5_ASAP7_75t_L g12111 ( 
.A1(n_10887),
.A2(n_9769),
.B(n_9187),
.C(n_9786),
.Y(n_12111)
);

AND2x2_ASAP7_75t_L g12112 ( 
.A(n_11523),
.B(n_9746),
.Y(n_12112)
);

AND2x2_ASAP7_75t_L g12113 ( 
.A(n_11523),
.B(n_9762),
.Y(n_12113)
);

OA22x2_ASAP7_75t_L g12114 ( 
.A1(n_10259),
.A2(n_9368),
.B1(n_9347),
.B2(n_9353),
.Y(n_12114)
);

O2A1O1Ixp5_ASAP7_75t_L g12115 ( 
.A1(n_10887),
.A2(n_9769),
.B(n_9187),
.C(n_9786),
.Y(n_12115)
);

INVx1_ASAP7_75t_L g12116 ( 
.A(n_10354),
.Y(n_12116)
);

AND2x2_ASAP7_75t_L g12117 ( 
.A(n_10365),
.B(n_9762),
.Y(n_12117)
);

AND2x2_ASAP7_75t_L g12118 ( 
.A(n_10365),
.B(n_9762),
.Y(n_12118)
);

INVx2_ASAP7_75t_L g12119 ( 
.A(n_10458),
.Y(n_12119)
);

AND2x2_ASAP7_75t_L g12120 ( 
.A(n_10365),
.B(n_10628),
.Y(n_12120)
);

AND2x2_ASAP7_75t_L g12121 ( 
.A(n_10365),
.B(n_10628),
.Y(n_12121)
);

AOI211xp5_ASAP7_75t_L g12122 ( 
.A1(n_11178),
.A2(n_9628),
.B(n_9655),
.C(n_9638),
.Y(n_12122)
);

NAND2xp5_ASAP7_75t_L g12123 ( 
.A(n_10977),
.B(n_8215),
.Y(n_12123)
);

INVx2_ASAP7_75t_SL g12124 ( 
.A(n_11431),
.Y(n_12124)
);

OR2x2_ASAP7_75t_L g12125 ( 
.A(n_10349),
.B(n_8198),
.Y(n_12125)
);

AOI21x1_ASAP7_75t_SL g12126 ( 
.A1(n_11017),
.A2(n_9437),
.B(n_9331),
.Y(n_12126)
);

INVx2_ASAP7_75t_L g12127 ( 
.A(n_10458),
.Y(n_12127)
);

O2A1O1Ixp5_ASAP7_75t_L g12128 ( 
.A1(n_11091),
.A2(n_9187),
.B(n_9786),
.C(n_9327),
.Y(n_12128)
);

INVx1_ASAP7_75t_L g12129 ( 
.A(n_10354),
.Y(n_12129)
);

AND2x2_ASAP7_75t_L g12130 ( 
.A(n_10628),
.B(n_9762),
.Y(n_12130)
);

INVx2_ASAP7_75t_L g12131 ( 
.A(n_10458),
.Y(n_12131)
);

OAI22xp5_ASAP7_75t_L g12132 ( 
.A1(n_10422),
.A2(n_9094),
.B1(n_9542),
.B2(n_9495),
.Y(n_12132)
);

OAI22xp5_ASAP7_75t_L g12133 ( 
.A1(n_10422),
.A2(n_9094),
.B1(n_9542),
.B2(n_9495),
.Y(n_12133)
);

AOI221x1_ASAP7_75t_SL g12134 ( 
.A1(n_10765),
.A2(n_9139),
.B1(n_9180),
.B2(n_9459),
.C(n_9457),
.Y(n_12134)
);

NAND2xp5_ASAP7_75t_L g12135 ( 
.A(n_10978),
.B(n_8215),
.Y(n_12135)
);

NAND2xp5_ASAP7_75t_L g12136 ( 
.A(n_10978),
.B(n_10727),
.Y(n_12136)
);

OAI22xp5_ASAP7_75t_L g12137 ( 
.A1(n_10585),
.A2(n_9542),
.B1(n_10079),
.B2(n_9495),
.Y(n_12137)
);

INVx1_ASAP7_75t_L g12138 ( 
.A(n_10356),
.Y(n_12138)
);

INVx2_ASAP7_75t_SL g12139 ( 
.A(n_11431),
.Y(n_12139)
);

NAND2xp5_ASAP7_75t_L g12140 ( 
.A(n_10727),
.B(n_8218),
.Y(n_12140)
);

AND2x2_ASAP7_75t_L g12141 ( 
.A(n_10628),
.B(n_9762),
.Y(n_12141)
);

INVx1_ASAP7_75t_L g12142 ( 
.A(n_10356),
.Y(n_12142)
);

HB1xp67_ASAP7_75t_L g12143 ( 
.A(n_10825),
.Y(n_12143)
);

AND2x2_ASAP7_75t_L g12144 ( 
.A(n_10628),
.B(n_9908),
.Y(n_12144)
);

A2O1A1Ixp33_ASAP7_75t_L g12145 ( 
.A1(n_10720),
.A2(n_9619),
.B(n_9811),
.C(n_9425),
.Y(n_12145)
);

INVx1_ASAP7_75t_L g12146 ( 
.A(n_10357),
.Y(n_12146)
);

O2A1O1Ixp33_ASAP7_75t_L g12147 ( 
.A1(n_11091),
.A2(n_9902),
.B(n_9368),
.C(n_9347),
.Y(n_12147)
);

AND2x2_ASAP7_75t_L g12148 ( 
.A(n_11016),
.B(n_9908),
.Y(n_12148)
);

BUFx6f_ASAP7_75t_L g12149 ( 
.A(n_10729),
.Y(n_12149)
);

INVx1_ASAP7_75t_L g12150 ( 
.A(n_10357),
.Y(n_12150)
);

INVx1_ASAP7_75t_L g12151 ( 
.A(n_10371),
.Y(n_12151)
);

INVx1_ASAP7_75t_L g12152 ( 
.A(n_10371),
.Y(n_12152)
);

AND2x2_ASAP7_75t_L g12153 ( 
.A(n_11016),
.B(n_9908),
.Y(n_12153)
);

INVx1_ASAP7_75t_L g12154 ( 
.A(n_10385),
.Y(n_12154)
);

NAND2xp5_ASAP7_75t_SL g12155 ( 
.A(n_10214),
.B(n_9668),
.Y(n_12155)
);

AND2x2_ASAP7_75t_L g12156 ( 
.A(n_11016),
.B(n_9908),
.Y(n_12156)
);

AND2x2_ASAP7_75t_L g12157 ( 
.A(n_11016),
.B(n_9908),
.Y(n_12157)
);

OAI22xp5_ASAP7_75t_SL g12158 ( 
.A1(n_10770),
.A2(n_10017),
.B1(n_9884),
.B2(n_9765),
.Y(n_12158)
);

OAI22xp5_ASAP7_75t_L g12159 ( 
.A1(n_10585),
.A2(n_10079),
.B1(n_9542),
.B2(n_9325),
.Y(n_12159)
);

AND2x2_ASAP7_75t_L g12160 ( 
.A(n_11016),
.B(n_9908),
.Y(n_12160)
);

AOI21x1_ASAP7_75t_SL g12161 ( 
.A1(n_10265),
.A2(n_9437),
.B(n_9331),
.Y(n_12161)
);

BUFx3_ASAP7_75t_L g12162 ( 
.A(n_10729),
.Y(n_12162)
);

AOI21xp5_ASAP7_75t_SL g12163 ( 
.A1(n_10564),
.A2(n_10162),
.B(n_10140),
.Y(n_12163)
);

NAND2x1p5_ASAP7_75t_L g12164 ( 
.A(n_11226),
.B(n_9587),
.Y(n_12164)
);

BUFx2_ASAP7_75t_L g12165 ( 
.A(n_10770),
.Y(n_12165)
);

AOI21xp5_ASAP7_75t_SL g12166 ( 
.A1(n_10617),
.A2(n_10162),
.B(n_10140),
.Y(n_12166)
);

AND2x4_ASAP7_75t_L g12167 ( 
.A(n_10393),
.B(n_9382),
.Y(n_12167)
);

AOI21x1_ASAP7_75t_SL g12168 ( 
.A1(n_10265),
.A2(n_11309),
.B(n_11302),
.Y(n_12168)
);

AOI21xp5_ASAP7_75t_SL g12169 ( 
.A1(n_10617),
.A2(n_10162),
.B(n_10140),
.Y(n_12169)
);

HB1xp67_ASAP7_75t_L g12170 ( 
.A(n_10825),
.Y(n_12170)
);

O2A1O1Ixp5_ASAP7_75t_L g12171 ( 
.A1(n_10214),
.A2(n_9327),
.B(n_9228),
.C(n_9223),
.Y(n_12171)
);

CKINVDCx5p33_ASAP7_75t_R g12172 ( 
.A(n_11073),
.Y(n_12172)
);

INVx2_ASAP7_75t_L g12173 ( 
.A(n_10458),
.Y(n_12173)
);

NAND2xp5_ASAP7_75t_L g12174 ( 
.A(n_10730),
.B(n_8218),
.Y(n_12174)
);

AOI21xp5_ASAP7_75t_L g12175 ( 
.A1(n_10850),
.A2(n_9953),
.B(n_9074),
.Y(n_12175)
);

OA21x2_ASAP7_75t_L g12176 ( 
.A1(n_10343),
.A2(n_8986),
.B(n_8985),
.Y(n_12176)
);

AND2x2_ASAP7_75t_L g12177 ( 
.A(n_11074),
.B(n_9908),
.Y(n_12177)
);

INVxp67_ASAP7_75t_SL g12178 ( 
.A(n_10458),
.Y(n_12178)
);

CKINVDCx20_ASAP7_75t_R g12179 ( 
.A(n_10445),
.Y(n_12179)
);

AOI21xp5_ASAP7_75t_SL g12180 ( 
.A1(n_11290),
.A2(n_10162),
.B(n_10140),
.Y(n_12180)
);

AND2x2_ASAP7_75t_L g12181 ( 
.A(n_11074),
.B(n_9908),
.Y(n_12181)
);

AND2x2_ASAP7_75t_L g12182 ( 
.A(n_11074),
.B(n_9908),
.Y(n_12182)
);

OAI22xp5_ASAP7_75t_L g12183 ( 
.A1(n_10667),
.A2(n_10079),
.B1(n_9542),
.B2(n_9325),
.Y(n_12183)
);

OAI22xp5_ASAP7_75t_L g12184 ( 
.A1(n_10667),
.A2(n_10079),
.B1(n_9542),
.B2(n_9325),
.Y(n_12184)
);

NAND2xp5_ASAP7_75t_L g12185 ( 
.A(n_10730),
.B(n_8220),
.Y(n_12185)
);

NAND2xp5_ASAP7_75t_L g12186 ( 
.A(n_11213),
.B(n_8220),
.Y(n_12186)
);

AOI21x1_ASAP7_75t_SL g12187 ( 
.A1(n_11302),
.A2(n_9298),
.B(n_9676),
.Y(n_12187)
);

AND2x4_ASAP7_75t_L g12188 ( 
.A(n_10597),
.B(n_9382),
.Y(n_12188)
);

NAND2x1p5_ASAP7_75t_L g12189 ( 
.A(n_10535),
.B(n_9587),
.Y(n_12189)
);

A2O1A1Ixp33_ASAP7_75t_SL g12190 ( 
.A1(n_11178),
.A2(n_8611),
.B(n_9095),
.C(n_9372),
.Y(n_12190)
);

AOI21xp5_ASAP7_75t_L g12191 ( 
.A1(n_10850),
.A2(n_9953),
.B(n_9074),
.Y(n_12191)
);

AND2x2_ASAP7_75t_L g12192 ( 
.A(n_11074),
.B(n_9915),
.Y(n_12192)
);

AOI21xp5_ASAP7_75t_L g12193 ( 
.A1(n_10940),
.A2(n_9953),
.B(n_9944),
.Y(n_12193)
);

INVx2_ASAP7_75t_L g12194 ( 
.A(n_10458),
.Y(n_12194)
);

AND2x2_ASAP7_75t_L g12195 ( 
.A(n_11074),
.B(n_9915),
.Y(n_12195)
);

BUFx12f_ASAP7_75t_L g12196 ( 
.A(n_10793),
.Y(n_12196)
);

AOI21xp5_ASAP7_75t_L g12197 ( 
.A1(n_10940),
.A2(n_9953),
.B(n_9944),
.Y(n_12197)
);

A2O1A1Ixp33_ASAP7_75t_L g12198 ( 
.A1(n_11290),
.A2(n_9619),
.B(n_9811),
.C(n_9425),
.Y(n_12198)
);

NAND2xp5_ASAP7_75t_L g12199 ( 
.A(n_11213),
.B(n_11257),
.Y(n_12199)
);

O2A1O1Ixp5_ASAP7_75t_L g12200 ( 
.A1(n_10214),
.A2(n_9327),
.B(n_9223),
.C(n_9228),
.Y(n_12200)
);

AOI21xp5_ASAP7_75t_L g12201 ( 
.A1(n_10716),
.A2(n_9944),
.B(n_9936),
.Y(n_12201)
);

OR2x2_ASAP7_75t_L g12202 ( 
.A(n_10349),
.B(n_8198),
.Y(n_12202)
);

OAI22xp5_ASAP7_75t_L g12203 ( 
.A1(n_10934),
.A2(n_10079),
.B1(n_9542),
.B2(n_9433),
.Y(n_12203)
);

HB1xp67_ASAP7_75t_L g12204 ( 
.A(n_10864),
.Y(n_12204)
);

A2O1A1Ixp33_ASAP7_75t_L g12205 ( 
.A1(n_11112),
.A2(n_9811),
.B(n_9425),
.C(n_9699),
.Y(n_12205)
);

OA22x2_ASAP7_75t_L g12206 ( 
.A1(n_11121),
.A2(n_10925),
.B1(n_11497),
.B2(n_10800),
.Y(n_12206)
);

A2O1A1Ixp33_ASAP7_75t_L g12207 ( 
.A1(n_11112),
.A2(n_9425),
.B(n_9699),
.C(n_9431),
.Y(n_12207)
);

OAI22xp5_ASAP7_75t_L g12208 ( 
.A1(n_10934),
.A2(n_10079),
.B1(n_9542),
.B2(n_9433),
.Y(n_12208)
);

HB1xp67_ASAP7_75t_L g12209 ( 
.A(n_10864),
.Y(n_12209)
);

NAND2xp5_ASAP7_75t_L g12210 ( 
.A(n_11257),
.B(n_8230),
.Y(n_12210)
);

HB1xp67_ASAP7_75t_L g12211 ( 
.A(n_10878),
.Y(n_12211)
);

INVx1_ASAP7_75t_L g12212 ( 
.A(n_10385),
.Y(n_12212)
);

BUFx3_ASAP7_75t_L g12213 ( 
.A(n_10793),
.Y(n_12213)
);

AND2x2_ASAP7_75t_L g12214 ( 
.A(n_11217),
.B(n_10203),
.Y(n_12214)
);

AOI21x1_ASAP7_75t_SL g12215 ( 
.A1(n_11309),
.A2(n_9298),
.B(n_9676),
.Y(n_12215)
);

INVx2_ASAP7_75t_L g12216 ( 
.A(n_10458),
.Y(n_12216)
);

BUFx3_ASAP7_75t_L g12217 ( 
.A(n_11431),
.Y(n_12217)
);

OR2x2_ASAP7_75t_L g12218 ( 
.A(n_10416),
.B(n_8198),
.Y(n_12218)
);

NAND2xp5_ASAP7_75t_L g12219 ( 
.A(n_11271),
.B(n_8230),
.Y(n_12219)
);

OAI22xp5_ASAP7_75t_L g12220 ( 
.A1(n_11071),
.A2(n_10079),
.B1(n_9433),
.B2(n_8888),
.Y(n_12220)
);

INVx1_ASAP7_75t_L g12221 ( 
.A(n_10394),
.Y(n_12221)
);

HB1xp67_ASAP7_75t_L g12222 ( 
.A(n_10878),
.Y(n_12222)
);

OAI211xp5_ASAP7_75t_L g12223 ( 
.A1(n_10366),
.A2(n_10162),
.B(n_10140),
.C(n_9228),
.Y(n_12223)
);

AND2x2_ASAP7_75t_L g12224 ( 
.A(n_11217),
.B(n_9915),
.Y(n_12224)
);

OAI22xp5_ASAP7_75t_L g12225 ( 
.A1(n_11071),
.A2(n_10079),
.B1(n_8888),
.B2(n_9285),
.Y(n_12225)
);

AOI21x1_ASAP7_75t_SL g12226 ( 
.A1(n_11321),
.A2(n_9298),
.B(n_9676),
.Y(n_12226)
);

HB1xp67_ASAP7_75t_L g12227 ( 
.A(n_10888),
.Y(n_12227)
);

AND2x2_ASAP7_75t_L g12228 ( 
.A(n_11217),
.B(n_10203),
.Y(n_12228)
);

AND2x4_ASAP7_75t_L g12229 ( 
.A(n_10597),
.B(n_9382),
.Y(n_12229)
);

AOI21xp5_ASAP7_75t_L g12230 ( 
.A1(n_10716),
.A2(n_9944),
.B(n_9936),
.Y(n_12230)
);

AOI21xp5_ASAP7_75t_L g12231 ( 
.A1(n_10811),
.A2(n_9944),
.B(n_9936),
.Y(n_12231)
);

OR2x2_ASAP7_75t_L g12232 ( 
.A(n_10416),
.B(n_8855),
.Y(n_12232)
);

OAI22xp5_ASAP7_75t_L g12233 ( 
.A1(n_11208),
.A2(n_8888),
.B1(n_9285),
.B2(n_9884),
.Y(n_12233)
);

NAND2xp5_ASAP7_75t_L g12234 ( 
.A(n_11271),
.B(n_11310),
.Y(n_12234)
);

AOI21xp5_ASAP7_75t_L g12235 ( 
.A1(n_10811),
.A2(n_9944),
.B(n_9936),
.Y(n_12235)
);

HB1xp67_ASAP7_75t_L g12236 ( 
.A(n_10888),
.Y(n_12236)
);

NAND2xp5_ASAP7_75t_L g12237 ( 
.A(n_11310),
.B(n_8231),
.Y(n_12237)
);

AOI21x1_ASAP7_75t_SL g12238 ( 
.A1(n_11321),
.A2(n_9680),
.B(n_9749),
.Y(n_12238)
);

AND2x2_ASAP7_75t_L g12239 ( 
.A(n_11217),
.B(n_9915),
.Y(n_12239)
);

HB1xp67_ASAP7_75t_L g12240 ( 
.A(n_10914),
.Y(n_12240)
);

AOI21x1_ASAP7_75t_SL g12241 ( 
.A1(n_11044),
.A2(n_11102),
.B(n_11097),
.Y(n_12241)
);

AOI21xp5_ASAP7_75t_L g12242 ( 
.A1(n_10925),
.A2(n_9944),
.B(n_9936),
.Y(n_12242)
);

AOI22xp5_ASAP7_75t_L g12243 ( 
.A1(n_10488),
.A2(n_11487),
.B1(n_10901),
.B2(n_10237),
.Y(n_12243)
);

INVx1_ASAP7_75t_SL g12244 ( 
.A(n_11409),
.Y(n_12244)
);

AOI21xp5_ASAP7_75t_L g12245 ( 
.A1(n_10800),
.A2(n_9944),
.B(n_9936),
.Y(n_12245)
);

AND2x2_ASAP7_75t_L g12246 ( 
.A(n_11217),
.B(n_9915),
.Y(n_12246)
);

NAND2xp5_ASAP7_75t_L g12247 ( 
.A(n_10554),
.B(n_8231),
.Y(n_12247)
);

OA21x2_ASAP7_75t_L g12248 ( 
.A1(n_10376),
.A2(n_8986),
.B(n_8985),
.Y(n_12248)
);

NAND2xp5_ASAP7_75t_L g12249 ( 
.A(n_10554),
.B(n_8233),
.Y(n_12249)
);

HB1xp67_ASAP7_75t_L g12250 ( 
.A(n_10914),
.Y(n_12250)
);

INVx1_ASAP7_75t_L g12251 ( 
.A(n_10394),
.Y(n_12251)
);

AOI21xp5_ASAP7_75t_L g12252 ( 
.A1(n_11121),
.A2(n_9936),
.B(n_10111),
.Y(n_12252)
);

AND2x2_ASAP7_75t_L g12253 ( 
.A(n_10203),
.B(n_9915),
.Y(n_12253)
);

CKINVDCx5p33_ASAP7_75t_R g12254 ( 
.A(n_11409),
.Y(n_12254)
);

HB1xp67_ASAP7_75t_L g12255 ( 
.A(n_10916),
.Y(n_12255)
);

AOI21x1_ASAP7_75t_SL g12256 ( 
.A1(n_11044),
.A2(n_9680),
.B(n_9749),
.Y(n_12256)
);

OA21x2_ASAP7_75t_L g12257 ( 
.A1(n_10376),
.A2(n_8986),
.B(n_8985),
.Y(n_12257)
);

OAI22xp5_ASAP7_75t_L g12258 ( 
.A1(n_11208),
.A2(n_9285),
.B1(n_9152),
.B2(n_8972),
.Y(n_12258)
);

NOR2x1_ASAP7_75t_L g12259 ( 
.A(n_11045),
.B(n_9765),
.Y(n_12259)
);

AND2x2_ASAP7_75t_L g12260 ( 
.A(n_10212),
.B(n_9915),
.Y(n_12260)
);

OR2x2_ASAP7_75t_L g12261 ( 
.A(n_11442),
.B(n_8855),
.Y(n_12261)
);

INVx1_ASAP7_75t_L g12262 ( 
.A(n_10395),
.Y(n_12262)
);

O2A1O1Ixp33_ASAP7_75t_L g12263 ( 
.A1(n_10869),
.A2(n_9902),
.B(n_9368),
.C(n_9347),
.Y(n_12263)
);

AOI21x1_ASAP7_75t_SL g12264 ( 
.A1(n_11097),
.A2(n_11126),
.B(n_11102),
.Y(n_12264)
);

INVx2_ASAP7_75t_L g12265 ( 
.A(n_10980),
.Y(n_12265)
);

O2A1O1Ixp5_ASAP7_75t_L g12266 ( 
.A1(n_10780),
.A2(n_9223),
.B(n_9638),
.C(n_9628),
.Y(n_12266)
);

INVx1_ASAP7_75t_L g12267 ( 
.A(n_10395),
.Y(n_12267)
);

AND2x4_ASAP7_75t_L g12268 ( 
.A(n_10597),
.B(n_9869),
.Y(n_12268)
);

INVx2_ASAP7_75t_SL g12269 ( 
.A(n_11431),
.Y(n_12269)
);

INVx1_ASAP7_75t_L g12270 ( 
.A(n_10401),
.Y(n_12270)
);

INVx1_ASAP7_75t_L g12271 ( 
.A(n_10401),
.Y(n_12271)
);

HB1xp67_ASAP7_75t_L g12272 ( 
.A(n_10916),
.Y(n_12272)
);

NOR2xp67_ASAP7_75t_L g12273 ( 
.A(n_11059),
.B(n_9669),
.Y(n_12273)
);

OA21x2_ASAP7_75t_L g12274 ( 
.A1(n_10376),
.A2(n_9006),
.B(n_9593),
.Y(n_12274)
);

HB1xp67_ASAP7_75t_L g12275 ( 
.A(n_11008),
.Y(n_12275)
);

O2A1O1Ixp33_ASAP7_75t_L g12276 ( 
.A1(n_10869),
.A2(n_9684),
.B(n_9771),
.C(n_9687),
.Y(n_12276)
);

AOI21xp5_ASAP7_75t_SL g12277 ( 
.A1(n_11059),
.A2(n_10162),
.B(n_10140),
.Y(n_12277)
);

AND2x2_ASAP7_75t_L g12278 ( 
.A(n_10212),
.B(n_9915),
.Y(n_12278)
);

AND2x4_ASAP7_75t_L g12279 ( 
.A(n_10597),
.B(n_9869),
.Y(n_12279)
);

OAI22xp5_ASAP7_75t_L g12280 ( 
.A1(n_11274),
.A2(n_9152),
.B1(n_8972),
.B2(n_8942),
.Y(n_12280)
);

O2A1O1Ixp5_ASAP7_75t_L g12281 ( 
.A1(n_10780),
.A2(n_9628),
.B(n_9655),
.C(n_9638),
.Y(n_12281)
);

O2A1O1Ixp5_ASAP7_75t_L g12282 ( 
.A1(n_10780),
.A2(n_9655),
.B(n_9790),
.C(n_9711),
.Y(n_12282)
);

OR2x2_ASAP7_75t_L g12283 ( 
.A(n_11442),
.B(n_8855),
.Y(n_12283)
);

INVx1_ASAP7_75t_SL g12284 ( 
.A(n_11308),
.Y(n_12284)
);

O2A1O1Ixp5_ASAP7_75t_L g12285 ( 
.A1(n_11200),
.A2(n_9711),
.B(n_9808),
.C(n_9790),
.Y(n_12285)
);

AND2x2_ASAP7_75t_L g12286 ( 
.A(n_10212),
.B(n_9915),
.Y(n_12286)
);

BUFx2_ASAP7_75t_L g12287 ( 
.A(n_10514),
.Y(n_12287)
);

O2A1O1Ixp33_ASAP7_75t_L g12288 ( 
.A1(n_11131),
.A2(n_9684),
.B(n_9771),
.C(n_9687),
.Y(n_12288)
);

INVx3_ASAP7_75t_L g12289 ( 
.A(n_10619),
.Y(n_12289)
);

CKINVDCx5p33_ASAP7_75t_R g12290 ( 
.A(n_10272),
.Y(n_12290)
);

AOI21xp5_ASAP7_75t_L g12291 ( 
.A1(n_10702),
.A2(n_9936),
.B(n_10111),
.Y(n_12291)
);

BUFx2_ASAP7_75t_L g12292 ( 
.A(n_10514),
.Y(n_12292)
);

O2A1O1Ixp33_ASAP7_75t_L g12293 ( 
.A1(n_11131),
.A2(n_11497),
.B(n_11622),
.C(n_11143),
.Y(n_12293)
);

OR2x2_ASAP7_75t_L g12294 ( 
.A(n_10714),
.B(n_10115),
.Y(n_12294)
);

AND2x2_ASAP7_75t_L g12295 ( 
.A(n_10218),
.B(n_9934),
.Y(n_12295)
);

OA21x2_ASAP7_75t_L g12296 ( 
.A1(n_11237),
.A2(n_11003),
.B(n_10957),
.Y(n_12296)
);

CKINVDCx20_ASAP7_75t_R g12297 ( 
.A(n_10812),
.Y(n_12297)
);

A2O1A1Ixp33_ASAP7_75t_L g12298 ( 
.A1(n_11120),
.A2(n_9699),
.B(n_9431),
.C(n_9737),
.Y(n_12298)
);

NAND2xp5_ASAP7_75t_L g12299 ( 
.A(n_10573),
.B(n_8233),
.Y(n_12299)
);

INVx1_ASAP7_75t_L g12300 ( 
.A(n_10406),
.Y(n_12300)
);

AND2x4_ASAP7_75t_L g12301 ( 
.A(n_10602),
.B(n_9869),
.Y(n_12301)
);

AND2x2_ASAP7_75t_L g12302 ( 
.A(n_10218),
.B(n_9934),
.Y(n_12302)
);

AND2x2_ASAP7_75t_L g12303 ( 
.A(n_10218),
.B(n_9934),
.Y(n_12303)
);

NOR2x1_ASAP7_75t_SL g12304 ( 
.A(n_11200),
.B(n_9574),
.Y(n_12304)
);

O2A1O1Ixp33_ASAP7_75t_L g12305 ( 
.A1(n_11622),
.A2(n_9684),
.B(n_9771),
.C(n_9687),
.Y(n_12305)
);

NAND2x1p5_ASAP7_75t_L g12306 ( 
.A(n_10535),
.B(n_9587),
.Y(n_12306)
);

INVx1_ASAP7_75t_L g12307 ( 
.A(n_10406),
.Y(n_12307)
);

AND2x2_ASAP7_75t_L g12308 ( 
.A(n_10607),
.B(n_9934),
.Y(n_12308)
);

OAI22xp5_ASAP7_75t_L g12309 ( 
.A1(n_11274),
.A2(n_9152),
.B1(n_8972),
.B2(n_8942),
.Y(n_12309)
);

O2A1O1Ixp33_ASAP7_75t_L g12310 ( 
.A1(n_11143),
.A2(n_9684),
.B(n_9771),
.C(n_9687),
.Y(n_12310)
);

AND2x2_ASAP7_75t_L g12311 ( 
.A(n_10607),
.B(n_9934),
.Y(n_12311)
);

INVx3_ASAP7_75t_L g12312 ( 
.A(n_10619),
.Y(n_12312)
);

HB1xp67_ASAP7_75t_L g12313 ( 
.A(n_11008),
.Y(n_12313)
);

OAI22xp5_ASAP7_75t_L g12314 ( 
.A1(n_11288),
.A2(n_8858),
.B1(n_7720),
.B2(n_9681),
.Y(n_12314)
);

AND2x2_ASAP7_75t_L g12315 ( 
.A(n_10607),
.B(n_9934),
.Y(n_12315)
);

NAND2xp5_ASAP7_75t_L g12316 ( 
.A(n_10573),
.B(n_8241),
.Y(n_12316)
);

O2A1O1Ixp5_ASAP7_75t_L g12317 ( 
.A1(n_11304),
.A2(n_9711),
.B(n_9808),
.C(n_9790),
.Y(n_12317)
);

AND2x2_ASAP7_75t_L g12318 ( 
.A(n_10790),
.B(n_9934),
.Y(n_12318)
);

AND2x2_ASAP7_75t_L g12319 ( 
.A(n_10790),
.B(n_9934),
.Y(n_12319)
);

INVx1_ASAP7_75t_L g12320 ( 
.A(n_10414),
.Y(n_12320)
);

OA21x2_ASAP7_75t_L g12321 ( 
.A1(n_11237),
.A2(n_9006),
.B(n_9593),
.Y(n_12321)
);

OA21x2_ASAP7_75t_L g12322 ( 
.A1(n_11237),
.A2(n_9006),
.B(n_9593),
.Y(n_12322)
);

AND2x2_ASAP7_75t_L g12323 ( 
.A(n_10790),
.B(n_9934),
.Y(n_12323)
);

O2A1O1Ixp33_ASAP7_75t_L g12324 ( 
.A1(n_11495),
.A2(n_9684),
.B(n_9771),
.C(n_9687),
.Y(n_12324)
);

AND2x2_ASAP7_75t_L g12325 ( 
.A(n_10801),
.B(n_9393),
.Y(n_12325)
);

AOI21xp5_ASAP7_75t_SL g12326 ( 
.A1(n_11304),
.A2(n_10162),
.B(n_9269),
.Y(n_12326)
);

INVx1_ASAP7_75t_L g12327 ( 
.A(n_10414),
.Y(n_12327)
);

O2A1O1Ixp33_ASAP7_75t_L g12328 ( 
.A1(n_11495),
.A2(n_11196),
.B(n_11475),
.C(n_10504),
.Y(n_12328)
);

AND2x2_ASAP7_75t_L g12329 ( 
.A(n_10801),
.B(n_9393),
.Y(n_12329)
);

INVx2_ASAP7_75t_L g12330 ( 
.A(n_10980),
.Y(n_12330)
);

INVx1_ASAP7_75t_L g12331 ( 
.A(n_10415),
.Y(n_12331)
);

NAND2xp5_ASAP7_75t_L g12332 ( 
.A(n_10714),
.B(n_8241),
.Y(n_12332)
);

INVxp33_ASAP7_75t_SL g12333 ( 
.A(n_10331),
.Y(n_12333)
);

OAI22xp5_ASAP7_75t_L g12334 ( 
.A1(n_11288),
.A2(n_8858),
.B1(n_7720),
.B2(n_9681),
.Y(n_12334)
);

INVx1_ASAP7_75t_L g12335 ( 
.A(n_10415),
.Y(n_12335)
);

AOI21x1_ASAP7_75t_SL g12336 ( 
.A1(n_11126),
.A2(n_9680),
.B(n_9749),
.Y(n_12336)
);

BUFx3_ASAP7_75t_L g12337 ( 
.A(n_11615),
.Y(n_12337)
);

O2A1O1Ixp33_ASAP7_75t_L g12338 ( 
.A1(n_11196),
.A2(n_9776),
.B(n_9095),
.C(n_10111),
.Y(n_12338)
);

AND2x2_ASAP7_75t_L g12339 ( 
.A(n_10801),
.B(n_9393),
.Y(n_12339)
);

NAND2xp5_ASAP7_75t_L g12340 ( 
.A(n_10505),
.B(n_8244),
.Y(n_12340)
);

AND2x4_ASAP7_75t_L g12341 ( 
.A(n_10602),
.B(n_9869),
.Y(n_12341)
);

NAND2xp5_ASAP7_75t_L g12342 ( 
.A(n_10505),
.B(n_8244),
.Y(n_12342)
);

OA21x2_ASAP7_75t_L g12343 ( 
.A1(n_11003),
.A2(n_9006),
.B(n_9593),
.Y(n_12343)
);

AOI21xp5_ASAP7_75t_L g12344 ( 
.A1(n_10702),
.A2(n_10111),
.B(n_9372),
.Y(n_12344)
);

INVxp67_ASAP7_75t_L g12345 ( 
.A(n_10535),
.Y(n_12345)
);

NOR3xp33_ASAP7_75t_L g12346 ( 
.A(n_11395),
.B(n_9180),
.C(n_9139),
.Y(n_12346)
);

BUFx6f_ASAP7_75t_L g12347 ( 
.A(n_11123),
.Y(n_12347)
);

O2A1O1Ixp33_ASAP7_75t_L g12348 ( 
.A1(n_11475),
.A2(n_9776),
.B(n_9095),
.C(n_10111),
.Y(n_12348)
);

NAND2xp5_ASAP7_75t_L g12349 ( 
.A(n_11435),
.B(n_8261),
.Y(n_12349)
);

OAI22xp5_ASAP7_75t_L g12350 ( 
.A1(n_11444),
.A2(n_8858),
.B1(n_7720),
.B2(n_9681),
.Y(n_12350)
);

O2A1O1Ixp5_ASAP7_75t_L g12351 ( 
.A1(n_11166),
.A2(n_9808),
.B(n_9861),
.C(n_9823),
.Y(n_12351)
);

INVx2_ASAP7_75t_L g12352 ( 
.A(n_10980),
.Y(n_12352)
);

BUFx2_ASAP7_75t_SL g12353 ( 
.A(n_10812),
.Y(n_12353)
);

AND2x2_ASAP7_75t_L g12354 ( 
.A(n_10923),
.B(n_9393),
.Y(n_12354)
);

OR2x2_ASAP7_75t_L g12355 ( 
.A(n_11435),
.B(n_10115),
.Y(n_12355)
);

AND2x2_ASAP7_75t_L g12356 ( 
.A(n_10923),
.B(n_9393),
.Y(n_12356)
);

AND2x2_ASAP7_75t_L g12357 ( 
.A(n_10923),
.B(n_10971),
.Y(n_12357)
);

INVx1_ASAP7_75t_L g12358 ( 
.A(n_10418),
.Y(n_12358)
);

BUFx3_ASAP7_75t_L g12359 ( 
.A(n_11615),
.Y(n_12359)
);

NAND2xp5_ASAP7_75t_L g12360 ( 
.A(n_11440),
.B(n_8261),
.Y(n_12360)
);

OAI22xp5_ASAP7_75t_L g12361 ( 
.A1(n_11444),
.A2(n_9681),
.B1(n_9444),
.B2(n_9647),
.Y(n_12361)
);

BUFx3_ASAP7_75t_L g12362 ( 
.A(n_11615),
.Y(n_12362)
);

OA21x2_ASAP7_75t_L g12363 ( 
.A1(n_11003),
.A2(n_10957),
.B(n_10953),
.Y(n_12363)
);

INVx2_ASAP7_75t_L g12364 ( 
.A(n_10980),
.Y(n_12364)
);

O2A1O1Ixp33_ASAP7_75t_L g12365 ( 
.A1(n_10504),
.A2(n_11395),
.B(n_11496),
.C(n_10764),
.Y(n_12365)
);

NAND2xp5_ASAP7_75t_L g12366 ( 
.A(n_11440),
.B(n_8270),
.Y(n_12366)
);

OA21x2_ASAP7_75t_L g12367 ( 
.A1(n_10953),
.A2(n_9006),
.B(n_9593),
.Y(n_12367)
);

INVx1_ASAP7_75t_L g12368 ( 
.A(n_10418),
.Y(n_12368)
);

OR2x2_ASAP7_75t_L g12369 ( 
.A(n_10450),
.B(n_10115),
.Y(n_12369)
);

HB1xp67_ASAP7_75t_L g12370 ( 
.A(n_11055),
.Y(n_12370)
);

INVx1_ASAP7_75t_SL g12371 ( 
.A(n_10948),
.Y(n_12371)
);

AOI21x1_ASAP7_75t_SL g12372 ( 
.A1(n_11413),
.A2(n_9826),
.B(n_9751),
.Y(n_12372)
);

BUFx3_ASAP7_75t_L g12373 ( 
.A(n_11615),
.Y(n_12373)
);

O2A1O1Ixp33_ASAP7_75t_L g12374 ( 
.A1(n_10504),
.A2(n_11496),
.B(n_10764),
.C(n_11385),
.Y(n_12374)
);

INVx2_ASAP7_75t_L g12375 ( 
.A(n_10980),
.Y(n_12375)
);

AOI21x1_ASAP7_75t_SL g12376 ( 
.A1(n_11413),
.A2(n_11420),
.B(n_11414),
.Y(n_12376)
);

INVx3_ASAP7_75t_L g12377 ( 
.A(n_10619),
.Y(n_12377)
);

A2O1A1Ixp33_ASAP7_75t_L g12378 ( 
.A1(n_11120),
.A2(n_9431),
.B(n_9743),
.C(n_9737),
.Y(n_12378)
);

AND2x2_ASAP7_75t_L g12379 ( 
.A(n_10971),
.B(n_9492),
.Y(n_12379)
);

INVx1_ASAP7_75t_L g12380 ( 
.A(n_10429),
.Y(n_12380)
);

AND2x2_ASAP7_75t_L g12381 ( 
.A(n_10971),
.B(n_9492),
.Y(n_12381)
);

A2O1A1Ixp33_ASAP7_75t_L g12382 ( 
.A1(n_11486),
.A2(n_9737),
.B(n_9760),
.C(n_9743),
.Y(n_12382)
);

OR2x2_ASAP7_75t_L g12383 ( 
.A(n_10450),
.B(n_10115),
.Y(n_12383)
);

AOI21xp5_ASAP7_75t_SL g12384 ( 
.A1(n_10535),
.A2(n_11486),
.B(n_11385),
.Y(n_12384)
);

NAND2xp5_ASAP7_75t_L g12385 ( 
.A(n_11350),
.B(n_8270),
.Y(n_12385)
);

AND2x2_ASAP7_75t_L g12386 ( 
.A(n_11333),
.B(n_9492),
.Y(n_12386)
);

OAI22xp5_ASAP7_75t_L g12387 ( 
.A1(n_11457),
.A2(n_9444),
.B1(n_9647),
.B2(n_9635),
.Y(n_12387)
);

INVx1_ASAP7_75t_L g12388 ( 
.A(n_10429),
.Y(n_12388)
);

NAND2xp5_ASAP7_75t_L g12389 ( 
.A(n_11350),
.B(n_8297),
.Y(n_12389)
);

AND2x2_ASAP7_75t_L g12390 ( 
.A(n_11333),
.B(n_9492),
.Y(n_12390)
);

A2O1A1Ixp33_ASAP7_75t_SL g12391 ( 
.A1(n_10285),
.A2(n_11100),
.B(n_11427),
.C(n_11194),
.Y(n_12391)
);

AND2x4_ASAP7_75t_L g12392 ( 
.A(n_10602),
.B(n_9869),
.Y(n_12392)
);

O2A1O1Ixp5_ASAP7_75t_L g12393 ( 
.A1(n_11166),
.A2(n_9823),
.B(n_9861),
.C(n_9635),
.Y(n_12393)
);

OAI22xp5_ASAP7_75t_L g12394 ( 
.A1(n_11457),
.A2(n_9444),
.B1(n_9647),
.B2(n_9635),
.Y(n_12394)
);

NAND2xp5_ASAP7_75t_L g12395 ( 
.A(n_11351),
.B(n_8297),
.Y(n_12395)
);

INVx1_ASAP7_75t_L g12396 ( 
.A(n_10436),
.Y(n_12396)
);

AOI21xp5_ASAP7_75t_L g12397 ( 
.A1(n_10488),
.A2(n_11010),
.B(n_11000),
.Y(n_12397)
);

AOI21x1_ASAP7_75t_SL g12398 ( 
.A1(n_11414),
.A2(n_11420),
.B(n_10671),
.Y(n_12398)
);

AOI21xp5_ASAP7_75t_SL g12399 ( 
.A1(n_10535),
.A2(n_10193),
.B(n_9402),
.Y(n_12399)
);

INVx4_ASAP7_75t_L g12400 ( 
.A(n_10514),
.Y(n_12400)
);

O2A1O1Ixp5_ASAP7_75t_L g12401 ( 
.A1(n_11166),
.A2(n_11010),
.B(n_11049),
.C(n_11000),
.Y(n_12401)
);

O2A1O1Ixp5_ASAP7_75t_L g12402 ( 
.A1(n_11049),
.A2(n_9861),
.B(n_9823),
.C(n_9735),
.Y(n_12402)
);

AND2x2_ASAP7_75t_L g12403 ( 
.A(n_11333),
.B(n_9492),
.Y(n_12403)
);

AOI21xp5_ASAP7_75t_SL g12404 ( 
.A1(n_10535),
.A2(n_10193),
.B(n_9402),
.Y(n_12404)
);

BUFx6f_ASAP7_75t_L g12405 ( 
.A(n_11123),
.Y(n_12405)
);

OAI22xp5_ASAP7_75t_L g12406 ( 
.A1(n_11510),
.A2(n_9444),
.B1(n_9647),
.B2(n_8934),
.Y(n_12406)
);

CKINVDCx16_ASAP7_75t_R g12407 ( 
.A(n_11593),
.Y(n_12407)
);

HB1xp67_ASAP7_75t_L g12408 ( 
.A(n_11055),
.Y(n_12408)
);

INVx1_ASAP7_75t_L g12409 ( 
.A(n_10436),
.Y(n_12409)
);

O2A1O1Ixp5_ASAP7_75t_L g12410 ( 
.A1(n_11154),
.A2(n_9735),
.B(n_9734),
.C(n_9051),
.Y(n_12410)
);

NAND2xp5_ASAP7_75t_L g12411 ( 
.A(n_11351),
.B(n_11355),
.Y(n_12411)
);

INVx3_ASAP7_75t_L g12412 ( 
.A(n_10619),
.Y(n_12412)
);

AND2x2_ASAP7_75t_L g12413 ( 
.A(n_11521),
.B(n_9499),
.Y(n_12413)
);

INVx1_ASAP7_75t_L g12414 ( 
.A(n_10501),
.Y(n_12414)
);

CKINVDCx16_ASAP7_75t_R g12415 ( 
.A(n_11593),
.Y(n_12415)
);

O2A1O1Ixp5_ASAP7_75t_L g12416 ( 
.A1(n_11154),
.A2(n_11391),
.B(n_11372),
.C(n_10844),
.Y(n_12416)
);

AND2x2_ASAP7_75t_L g12417 ( 
.A(n_11521),
.B(n_9499),
.Y(n_12417)
);

NOR2xp67_ASAP7_75t_L g12418 ( 
.A(n_11268),
.B(n_9669),
.Y(n_12418)
);

O2A1O1Ixp5_ASAP7_75t_L g12419 ( 
.A1(n_11372),
.A2(n_9735),
.B(n_9734),
.C(n_9051),
.Y(n_12419)
);

INVx4_ASAP7_75t_SL g12420 ( 
.A(n_10644),
.Y(n_12420)
);

OA21x2_ASAP7_75t_L g12421 ( 
.A1(n_10953),
.A2(n_9006),
.B(n_9593),
.Y(n_12421)
);

NAND2xp5_ASAP7_75t_L g12422 ( 
.A(n_11355),
.B(n_10430),
.Y(n_12422)
);

AOI21xp5_ASAP7_75t_L g12423 ( 
.A1(n_11263),
.A2(n_10111),
.B(n_9372),
.Y(n_12423)
);

O2A1O1Ixp33_ASAP7_75t_L g12424 ( 
.A1(n_10764),
.A2(n_9776),
.B(n_10111),
.C(n_10097),
.Y(n_12424)
);

AND2x2_ASAP7_75t_L g12425 ( 
.A(n_11521),
.B(n_9499),
.Y(n_12425)
);

INVx1_ASAP7_75t_L g12426 ( 
.A(n_10501),
.Y(n_12426)
);

AOI21xp5_ASAP7_75t_SL g12427 ( 
.A1(n_10602),
.A2(n_10193),
.B(n_9402),
.Y(n_12427)
);

INVx1_ASAP7_75t_L g12428 ( 
.A(n_10508),
.Y(n_12428)
);

AOI21xp5_ASAP7_75t_SL g12429 ( 
.A1(n_10604),
.A2(n_10193),
.B(n_9402),
.Y(n_12429)
);

AOI21xp5_ASAP7_75t_L g12430 ( 
.A1(n_11263),
.A2(n_10111),
.B(n_10097),
.Y(n_12430)
);

AOI21x1_ASAP7_75t_SL g12431 ( 
.A1(n_10587),
.A2(n_10693),
.B(n_10671),
.Y(n_12431)
);

AND2x2_ASAP7_75t_L g12432 ( 
.A(n_11536),
.B(n_9499),
.Y(n_12432)
);

INVx1_ASAP7_75t_L g12433 ( 
.A(n_10508),
.Y(n_12433)
);

INVx1_ASAP7_75t_L g12434 ( 
.A(n_10510),
.Y(n_12434)
);

AOI21xp5_ASAP7_75t_L g12435 ( 
.A1(n_10844),
.A2(n_10538),
.B(n_10517),
.Y(n_12435)
);

AOI31xp33_ASAP7_75t_L g12436 ( 
.A1(n_11427),
.A2(n_8650),
.A3(n_8671),
.B(n_8634),
.Y(n_12436)
);

BUFx3_ASAP7_75t_L g12437 ( 
.A(n_11615),
.Y(n_12437)
);

AND2x2_ASAP7_75t_L g12438 ( 
.A(n_11536),
.B(n_9499),
.Y(n_12438)
);

AND2x2_ASAP7_75t_L g12439 ( 
.A(n_11536),
.B(n_7771),
.Y(n_12439)
);

AND2x2_ASAP7_75t_L g12440 ( 
.A(n_11405),
.B(n_7771),
.Y(n_12440)
);

OAI22xp5_ASAP7_75t_L g12441 ( 
.A1(n_11510),
.A2(n_9444),
.B1(n_8934),
.B2(n_9774),
.Y(n_12441)
);

AOI21x1_ASAP7_75t_SL g12442 ( 
.A1(n_10587),
.A2(n_9826),
.B(n_9751),
.Y(n_12442)
);

HB1xp67_ASAP7_75t_L g12443 ( 
.A(n_10577),
.Y(n_12443)
);

AND2x4_ASAP7_75t_L g12444 ( 
.A(n_10604),
.B(n_9382),
.Y(n_12444)
);

BUFx4f_ASAP7_75t_SL g12445 ( 
.A(n_10696),
.Y(n_12445)
);

AOI21x1_ASAP7_75t_SL g12446 ( 
.A1(n_10693),
.A2(n_9826),
.B(n_9751),
.Y(n_12446)
);

AND2x2_ASAP7_75t_L g12447 ( 
.A(n_11405),
.B(n_7771),
.Y(n_12447)
);

AND2x2_ASAP7_75t_L g12448 ( 
.A(n_11405),
.B(n_7771),
.Y(n_12448)
);

INVx3_ASAP7_75t_L g12449 ( 
.A(n_10619),
.Y(n_12449)
);

NAND2xp5_ASAP7_75t_L g12450 ( 
.A(n_10430),
.B(n_8301),
.Y(n_12450)
);

OA21x2_ASAP7_75t_L g12451 ( 
.A1(n_10957),
.A2(n_9605),
.B(n_9604),
.Y(n_12451)
);

OR2x2_ASAP7_75t_L g12452 ( 
.A(n_10471),
.B(n_10115),
.Y(n_12452)
);

A2O1A1Ixp33_ASAP7_75t_L g12453 ( 
.A1(n_10517),
.A2(n_10538),
.B(n_11206),
.C(n_11004),
.Y(n_12453)
);

INVx5_ASAP7_75t_L g12454 ( 
.A(n_10734),
.Y(n_12454)
);

OR2x2_ASAP7_75t_L g12455 ( 
.A(n_10471),
.B(n_10115),
.Y(n_12455)
);

O2A1O1Ixp5_ASAP7_75t_L g12456 ( 
.A1(n_11372),
.A2(n_9734),
.B(n_9051),
.C(n_9240),
.Y(n_12456)
);

OAI22xp5_ASAP7_75t_L g12457 ( 
.A1(n_11608),
.A2(n_9444),
.B1(n_9780),
.B2(n_9774),
.Y(n_12457)
);

OAI22xp5_ASAP7_75t_L g12458 ( 
.A1(n_11608),
.A2(n_9444),
.B1(n_9780),
.B2(n_9774),
.Y(n_12458)
);

NAND2xp5_ASAP7_75t_L g12459 ( 
.A(n_10503),
.B(n_8301),
.Y(n_12459)
);

AND2x2_ASAP7_75t_L g12460 ( 
.A(n_11405),
.B(n_7771),
.Y(n_12460)
);

OA21x2_ASAP7_75t_L g12461 ( 
.A1(n_10973),
.A2(n_9605),
.B(n_9604),
.Y(n_12461)
);

NAND2xp5_ASAP7_75t_L g12462 ( 
.A(n_10503),
.B(n_8302),
.Y(n_12462)
);

INVx1_ASAP7_75t_L g12463 ( 
.A(n_10510),
.Y(n_12463)
);

AOI21xp5_ASAP7_75t_L g12464 ( 
.A1(n_11225),
.A2(n_10097),
.B(n_9760),
.Y(n_12464)
);

HB1xp67_ASAP7_75t_L g12465 ( 
.A(n_10577),
.Y(n_12465)
);

INVx1_ASAP7_75t_L g12466 ( 
.A(n_10515),
.Y(n_12466)
);

OR2x2_ASAP7_75t_L g12467 ( 
.A(n_10528),
.B(n_10115),
.Y(n_12467)
);

O2A1O1Ixp33_ASAP7_75t_L g12468 ( 
.A1(n_11194),
.A2(n_9776),
.B(n_10097),
.C(n_9597),
.Y(n_12468)
);

INVx1_ASAP7_75t_L g12469 ( 
.A(n_10515),
.Y(n_12469)
);

OAI22xp5_ASAP7_75t_L g12470 ( 
.A1(n_11004),
.A2(n_9444),
.B1(n_9780),
.B2(n_8542),
.Y(n_12470)
);

OA21x2_ASAP7_75t_L g12471 ( 
.A1(n_10973),
.A2(n_9605),
.B(n_9604),
.Y(n_12471)
);

NOR2xp33_ASAP7_75t_L g12472 ( 
.A(n_10434),
.B(n_9509),
.Y(n_12472)
);

INVx1_ASAP7_75t_L g12473 ( 
.A(n_10520),
.Y(n_12473)
);

AND2x4_ASAP7_75t_L g12474 ( 
.A(n_10604),
.B(n_9382),
.Y(n_12474)
);

OR2x2_ASAP7_75t_L g12475 ( 
.A(n_10528),
.B(n_10115),
.Y(n_12475)
);

INVx1_ASAP7_75t_L g12476 ( 
.A(n_10520),
.Y(n_12476)
);

AND2x2_ASAP7_75t_L g12477 ( 
.A(n_11447),
.B(n_7771),
.Y(n_12477)
);

AND2x2_ASAP7_75t_L g12478 ( 
.A(n_11447),
.B(n_7785),
.Y(n_12478)
);

INVx1_ASAP7_75t_L g12479 ( 
.A(n_10521),
.Y(n_12479)
);

AOI221xp5_ASAP7_75t_L g12480 ( 
.A1(n_11243),
.A2(n_9892),
.B1(n_9911),
.B2(n_9872),
.C(n_9838),
.Y(n_12480)
);

NOR2xp33_ASAP7_75t_R g12481 ( 
.A(n_10696),
.B(n_9669),
.Y(n_12481)
);

INVx1_ASAP7_75t_L g12482 ( 
.A(n_10521),
.Y(n_12482)
);

NAND2xp5_ASAP7_75t_L g12483 ( 
.A(n_11324),
.B(n_8302),
.Y(n_12483)
);

INVx1_ASAP7_75t_L g12484 ( 
.A(n_10523),
.Y(n_12484)
);

AND2x2_ASAP7_75t_L g12485 ( 
.A(n_11447),
.B(n_7785),
.Y(n_12485)
);

OR2x2_ASAP7_75t_L g12486 ( 
.A(n_10703),
.B(n_10115),
.Y(n_12486)
);

OAI22xp5_ASAP7_75t_L g12487 ( 
.A1(n_11365),
.A2(n_9444),
.B1(n_9016),
.B2(n_9098),
.Y(n_12487)
);

AND2x2_ASAP7_75t_L g12488 ( 
.A(n_11447),
.B(n_7785),
.Y(n_12488)
);

INVx1_ASAP7_75t_L g12489 ( 
.A(n_10523),
.Y(n_12489)
);

INVx1_ASAP7_75t_L g12490 ( 
.A(n_10524),
.Y(n_12490)
);

AND2x2_ASAP7_75t_L g12491 ( 
.A(n_11471),
.B(n_7785),
.Y(n_12491)
);

AND2x4_ASAP7_75t_L g12492 ( 
.A(n_10604),
.B(n_9382),
.Y(n_12492)
);

AND2x2_ASAP7_75t_L g12493 ( 
.A(n_11471),
.B(n_7785),
.Y(n_12493)
);

OAI22xp33_ASAP7_75t_L g12494 ( 
.A1(n_11206),
.A2(n_9010),
.B1(n_8458),
.B2(n_8197),
.Y(n_12494)
);

CKINVDCx20_ASAP7_75t_R g12495 ( 
.A(n_10948),
.Y(n_12495)
);

OA21x2_ASAP7_75t_L g12496 ( 
.A1(n_10973),
.A2(n_9605),
.B(n_9604),
.Y(n_12496)
);

HB1xp67_ASAP7_75t_L g12497 ( 
.A(n_10577),
.Y(n_12497)
);

AND2x4_ASAP7_75t_L g12498 ( 
.A(n_10665),
.B(n_9390),
.Y(n_12498)
);

AND2x2_ASAP7_75t_L g12499 ( 
.A(n_11471),
.B(n_7785),
.Y(n_12499)
);

BUFx8_ASAP7_75t_SL g12500 ( 
.A(n_10447),
.Y(n_12500)
);

NAND2xp5_ASAP7_75t_L g12501 ( 
.A(n_11324),
.B(n_8303),
.Y(n_12501)
);

OR2x6_ASAP7_75t_L g12502 ( 
.A(n_11280),
.B(n_9798),
.Y(n_12502)
);

NOR2xp33_ASAP7_75t_L g12503 ( 
.A(n_10512),
.B(n_10536),
.Y(n_12503)
);

AOI21xp5_ASAP7_75t_L g12504 ( 
.A1(n_11225),
.A2(n_10097),
.B(n_9760),
.Y(n_12504)
);

AND2x2_ASAP7_75t_L g12505 ( 
.A(n_11471),
.B(n_7915),
.Y(n_12505)
);

AND2x2_ASAP7_75t_L g12506 ( 
.A(n_11485),
.B(n_7915),
.Y(n_12506)
);

AOI21xp5_ASAP7_75t_L g12507 ( 
.A1(n_11225),
.A2(n_10097),
.B(n_9743),
.Y(n_12507)
);

OR2x2_ASAP7_75t_L g12508 ( 
.A(n_10703),
.B(n_10115),
.Y(n_12508)
);

O2A1O1Ixp33_ASAP7_75t_L g12509 ( 
.A1(n_10194),
.A2(n_9776),
.B(n_10097),
.C(n_9597),
.Y(n_12509)
);

A2O1A1Ixp33_ASAP7_75t_L g12510 ( 
.A1(n_11181),
.A2(n_9010),
.B(n_9665),
.C(n_9488),
.Y(n_12510)
);

CKINVDCx5p33_ASAP7_75t_R g12511 ( 
.A(n_10686),
.Y(n_12511)
);

INVx1_ASAP7_75t_L g12512 ( 
.A(n_10524),
.Y(n_12512)
);

AND2x2_ASAP7_75t_L g12513 ( 
.A(n_11485),
.B(n_7915),
.Y(n_12513)
);

AND2x4_ASAP7_75t_L g12514 ( 
.A(n_10665),
.B(n_9390),
.Y(n_12514)
);

AOI21xp5_ASAP7_75t_SL g12515 ( 
.A1(n_10665),
.A2(n_9910),
.B(n_9210),
.Y(n_12515)
);

AND2x2_ASAP7_75t_L g12516 ( 
.A(n_11485),
.B(n_7915),
.Y(n_12516)
);

AOI21x1_ASAP7_75t_SL g12517 ( 
.A1(n_10713),
.A2(n_11266),
.B(n_11254),
.Y(n_12517)
);

AOI21xp5_ASAP7_75t_L g12518 ( 
.A1(n_11225),
.A2(n_10097),
.B(n_9010),
.Y(n_12518)
);

OR2x2_ASAP7_75t_L g12519 ( 
.A(n_11599),
.B(n_10115),
.Y(n_12519)
);

OR2x2_ASAP7_75t_L g12520 ( 
.A(n_11599),
.B(n_10115),
.Y(n_12520)
);

INVxp67_ASAP7_75t_SL g12521 ( 
.A(n_10358),
.Y(n_12521)
);

NAND2xp5_ASAP7_75t_L g12522 ( 
.A(n_11254),
.B(n_8303),
.Y(n_12522)
);

INVx1_ASAP7_75t_L g12523 ( 
.A(n_10526),
.Y(n_12523)
);

A2O1A1Ixp33_ASAP7_75t_L g12524 ( 
.A1(n_11181),
.A2(n_11093),
.B(n_11079),
.C(n_11222),
.Y(n_12524)
);

NAND2xp5_ASAP7_75t_L g12525 ( 
.A(n_11266),
.B(n_8304),
.Y(n_12525)
);

AND2x2_ASAP7_75t_L g12526 ( 
.A(n_11485),
.B(n_7915),
.Y(n_12526)
);

INVx2_ASAP7_75t_L g12527 ( 
.A(n_10980),
.Y(n_12527)
);

AOI21x1_ASAP7_75t_SL g12528 ( 
.A1(n_10713),
.A2(n_9716),
.B(n_9702),
.Y(n_12528)
);

INVx1_ASAP7_75t_L g12529 ( 
.A(n_10526),
.Y(n_12529)
);

O2A1O1Ixp33_ASAP7_75t_L g12530 ( 
.A1(n_10194),
.A2(n_9597),
.B(n_9233),
.C(n_9116),
.Y(n_12530)
);

AOI211xp5_ASAP7_75t_L g12531 ( 
.A1(n_11360),
.A2(n_9007),
.B(n_9098),
.C(n_9016),
.Y(n_12531)
);

NAND2xp5_ASAP7_75t_L g12532 ( 
.A(n_11291),
.B(n_8304),
.Y(n_12532)
);

AND2x2_ASAP7_75t_L g12533 ( 
.A(n_11587),
.B(n_7915),
.Y(n_12533)
);

O2A1O1Ixp5_ASAP7_75t_L g12534 ( 
.A1(n_11391),
.A2(n_9210),
.B(n_9240),
.C(n_9051),
.Y(n_12534)
);

INVx1_ASAP7_75t_L g12535 ( 
.A(n_10537),
.Y(n_12535)
);

AND2x2_ASAP7_75t_L g12536 ( 
.A(n_11587),
.B(n_7952),
.Y(n_12536)
);

INVx1_ASAP7_75t_SL g12537 ( 
.A(n_11067),
.Y(n_12537)
);

INVx2_ASAP7_75t_L g12538 ( 
.A(n_10980),
.Y(n_12538)
);

INVx2_ASAP7_75t_L g12539 ( 
.A(n_10980),
.Y(n_12539)
);

AOI21x1_ASAP7_75t_SL g12540 ( 
.A1(n_11291),
.A2(n_9716),
.B(n_9702),
.Y(n_12540)
);

AND2x2_ASAP7_75t_L g12541 ( 
.A(n_11587),
.B(n_7952),
.Y(n_12541)
);

NAND2xp5_ASAP7_75t_L g12542 ( 
.A(n_11294),
.B(n_8311),
.Y(n_12542)
);

AND2x2_ASAP7_75t_L g12543 ( 
.A(n_11587),
.B(n_7952),
.Y(n_12543)
);

INVx1_ASAP7_75t_L g12544 ( 
.A(n_10537),
.Y(n_12544)
);

AND2x2_ASAP7_75t_SL g12545 ( 
.A(n_10734),
.B(n_9010),
.Y(n_12545)
);

NAND2xp5_ASAP7_75t_L g12546 ( 
.A(n_11294),
.B(n_8311),
.Y(n_12546)
);

OAI22xp5_ASAP7_75t_L g12547 ( 
.A1(n_11365),
.A2(n_9444),
.B1(n_9016),
.B2(n_9098),
.Y(n_12547)
);

NOR2xp33_ASAP7_75t_L g12548 ( 
.A(n_11067),
.B(n_9509),
.Y(n_12548)
);

NAND2xp5_ASAP7_75t_L g12549 ( 
.A(n_11581),
.B(n_8318),
.Y(n_12549)
);

BUFx6f_ASAP7_75t_L g12550 ( 
.A(n_11188),
.Y(n_12550)
);

AND2x4_ASAP7_75t_L g12551 ( 
.A(n_10665),
.B(n_10847),
.Y(n_12551)
);

OR2x2_ASAP7_75t_L g12552 ( 
.A(n_11568),
.B(n_10115),
.Y(n_12552)
);

OR2x2_ASAP7_75t_L g12553 ( 
.A(n_11568),
.B(n_7899),
.Y(n_12553)
);

AND2x2_ASAP7_75t_L g12554 ( 
.A(n_10318),
.B(n_7952),
.Y(n_12554)
);

AOI21xp5_ASAP7_75t_L g12555 ( 
.A1(n_11079),
.A2(n_9233),
.B(n_9937),
.Y(n_12555)
);

OA21x2_ASAP7_75t_L g12556 ( 
.A1(n_10677),
.A2(n_9605),
.B(n_9604),
.Y(n_12556)
);

HB1xp67_ASAP7_75t_L g12557 ( 
.A(n_10577),
.Y(n_12557)
);

AOI21xp5_ASAP7_75t_L g12558 ( 
.A1(n_11093),
.A2(n_9233),
.B(n_9937),
.Y(n_12558)
);

NAND2xp5_ASAP7_75t_L g12559 ( 
.A(n_11581),
.B(n_8318),
.Y(n_12559)
);

O2A1O1Ixp33_ASAP7_75t_L g12560 ( 
.A1(n_10194),
.A2(n_9597),
.B(n_9115),
.C(n_9116),
.Y(n_12560)
);

HB1xp67_ASAP7_75t_L g12561 ( 
.A(n_10577),
.Y(n_12561)
);

NAND2x1p5_ASAP7_75t_L g12562 ( 
.A(n_11100),
.B(n_9587),
.Y(n_12562)
);

BUFx3_ASAP7_75t_L g12563 ( 
.A(n_10696),
.Y(n_12563)
);

NAND2xp5_ASAP7_75t_L g12564 ( 
.A(n_11329),
.B(n_8331),
.Y(n_12564)
);

AOI221xp5_ASAP7_75t_L g12565 ( 
.A1(n_11360),
.A2(n_9892),
.B1(n_9911),
.B2(n_9872),
.C(n_9838),
.Y(n_12565)
);

AND2x2_ASAP7_75t_L g12566 ( 
.A(n_10318),
.B(n_7952),
.Y(n_12566)
);

INVx1_ASAP7_75t_L g12567 ( 
.A(n_10541),
.Y(n_12567)
);

NAND2xp5_ASAP7_75t_L g12568 ( 
.A(n_11329),
.B(n_8331),
.Y(n_12568)
);

BUFx3_ASAP7_75t_L g12569 ( 
.A(n_11453),
.Y(n_12569)
);

HB1xp67_ASAP7_75t_L g12570 ( 
.A(n_10439),
.Y(n_12570)
);

OAI22xp5_ASAP7_75t_L g12571 ( 
.A1(n_10236),
.A2(n_9444),
.B1(n_9016),
.B2(n_9098),
.Y(n_12571)
);

O2A1O1Ixp5_ASAP7_75t_L g12572 ( 
.A1(n_11391),
.A2(n_9051),
.B(n_9240),
.C(n_9210),
.Y(n_12572)
);

NAND2xp5_ASAP7_75t_L g12573 ( 
.A(n_11356),
.B(n_8587),
.Y(n_12573)
);

OAI22xp5_ASAP7_75t_L g12574 ( 
.A1(n_10236),
.A2(n_9016),
.B1(n_9098),
.B2(n_9051),
.Y(n_12574)
);

AOI221x1_ASAP7_75t_SL g12575 ( 
.A1(n_10676),
.A2(n_9796),
.B1(n_9843),
.B2(n_9809),
.C(n_9787),
.Y(n_12575)
);

HB1xp67_ASAP7_75t_L g12576 ( 
.A(n_10439),
.Y(n_12576)
);

INVx1_ASAP7_75t_L g12577 ( 
.A(n_10541),
.Y(n_12577)
);

INVx1_ASAP7_75t_L g12578 ( 
.A(n_10543),
.Y(n_12578)
);

O2A1O1Ixp33_ASAP7_75t_L g12579 ( 
.A1(n_11546),
.A2(n_9115),
.B(n_9116),
.C(n_9927),
.Y(n_12579)
);

OR2x2_ASAP7_75t_L g12580 ( 
.A(n_11601),
.B(n_8120),
.Y(n_12580)
);

AOI21xp5_ASAP7_75t_L g12581 ( 
.A1(n_11222),
.A2(n_9937),
.B(n_9385),
.Y(n_12581)
);

INVx3_ASAP7_75t_SL g12582 ( 
.A(n_11295),
.Y(n_12582)
);

AOI21xp5_ASAP7_75t_L g12583 ( 
.A1(n_11228),
.A2(n_9937),
.B(n_9385),
.Y(n_12583)
);

CKINVDCx5p33_ASAP7_75t_R g12584 ( 
.A(n_10772),
.Y(n_12584)
);

OA21x2_ASAP7_75t_L g12585 ( 
.A1(n_10677),
.A2(n_9605),
.B(n_9604),
.Y(n_12585)
);

INVx2_ASAP7_75t_L g12586 ( 
.A(n_11503),
.Y(n_12586)
);

AND2x2_ASAP7_75t_L g12587 ( 
.A(n_10318),
.B(n_7952),
.Y(n_12587)
);

INVx2_ASAP7_75t_L g12588 ( 
.A(n_11503),
.Y(n_12588)
);

HB1xp67_ASAP7_75t_L g12589 ( 
.A(n_10455),
.Y(n_12589)
);

INVx1_ASAP7_75t_L g12590 ( 
.A(n_10543),
.Y(n_12590)
);

AOI21x1_ASAP7_75t_SL g12591 ( 
.A1(n_11298),
.A2(n_9716),
.B(n_9702),
.Y(n_12591)
);

OAI22xp5_ASAP7_75t_L g12592 ( 
.A1(n_10721),
.A2(n_9051),
.B1(n_9240),
.B2(n_9210),
.Y(n_12592)
);

INVx6_ASAP7_75t_L g12593 ( 
.A(n_10271),
.Y(n_12593)
);

INVx2_ASAP7_75t_L g12594 ( 
.A(n_11503),
.Y(n_12594)
);

INVx1_ASAP7_75t_L g12595 ( 
.A(n_10565),
.Y(n_12595)
);

AOI21xp5_ASAP7_75t_SL g12596 ( 
.A1(n_10847),
.A2(n_9910),
.B(n_9210),
.Y(n_12596)
);

OR2x2_ASAP7_75t_L g12597 ( 
.A(n_11601),
.B(n_8120),
.Y(n_12597)
);

AOI21x1_ASAP7_75t_SL g12598 ( 
.A1(n_11298),
.A2(n_9721),
.B(n_9720),
.Y(n_12598)
);

AOI21x1_ASAP7_75t_SL g12599 ( 
.A1(n_11316),
.A2(n_9721),
.B(n_9720),
.Y(n_12599)
);

AND2x2_ASAP7_75t_L g12600 ( 
.A(n_10318),
.B(n_8038),
.Y(n_12600)
);

NAND2xp5_ASAP7_75t_L g12601 ( 
.A(n_11356),
.B(n_8587),
.Y(n_12601)
);

NOR2x1_ASAP7_75t_SL g12602 ( 
.A(n_10626),
.B(n_9574),
.Y(n_12602)
);

HB1xp67_ASAP7_75t_L g12603 ( 
.A(n_10455),
.Y(n_12603)
);

AOI21xp5_ASAP7_75t_SL g12604 ( 
.A1(n_10847),
.A2(n_9210),
.B(n_9051),
.Y(n_12604)
);

CKINVDCx5p33_ASAP7_75t_R g12605 ( 
.A(n_11453),
.Y(n_12605)
);

CKINVDCx11_ASAP7_75t_R g12606 ( 
.A(n_11188),
.Y(n_12606)
);

OAI22xp5_ASAP7_75t_L g12607 ( 
.A1(n_10721),
.A2(n_9210),
.B1(n_9243),
.B2(n_9240),
.Y(n_12607)
);

AND2x2_ASAP7_75t_L g12608 ( 
.A(n_10318),
.B(n_8038),
.Y(n_12608)
);

O2A1O1Ixp5_ASAP7_75t_L g12609 ( 
.A1(n_11584),
.A2(n_9210),
.B(n_9243),
.C(n_9240),
.Y(n_12609)
);

INVx2_ASAP7_75t_L g12610 ( 
.A(n_10540),
.Y(n_12610)
);

AND2x2_ASAP7_75t_L g12611 ( 
.A(n_10323),
.B(n_8038),
.Y(n_12611)
);

OAI22xp5_ASAP7_75t_L g12612 ( 
.A1(n_11466),
.A2(n_9240),
.B1(n_9354),
.B2(n_9243),
.Y(n_12612)
);

INVx2_ASAP7_75t_L g12613 ( 
.A(n_10540),
.Y(n_12613)
);

NAND2xp5_ASAP7_75t_L g12614 ( 
.A(n_11394),
.B(n_11403),
.Y(n_12614)
);

BUFx2_ASAP7_75t_L g12615 ( 
.A(n_10271),
.Y(n_12615)
);

AOI21xp5_ASAP7_75t_L g12616 ( 
.A1(n_11228),
.A2(n_9937),
.B(n_9385),
.Y(n_12616)
);

AND2x2_ASAP7_75t_L g12617 ( 
.A(n_10323),
.B(n_8038),
.Y(n_12617)
);

BUFx2_ASAP7_75t_R g12618 ( 
.A(n_10644),
.Y(n_12618)
);

BUFx10_ASAP7_75t_L g12619 ( 
.A(n_11334),
.Y(n_12619)
);

AND2x2_ASAP7_75t_L g12620 ( 
.A(n_10323),
.B(n_8038),
.Y(n_12620)
);

NAND2xp5_ASAP7_75t_L g12621 ( 
.A(n_11394),
.B(n_8127),
.Y(n_12621)
);

O2A1O1Ixp33_ASAP7_75t_L g12622 ( 
.A1(n_11546),
.A2(n_11584),
.B(n_10358),
.C(n_11526),
.Y(n_12622)
);

OAI22xp5_ASAP7_75t_L g12623 ( 
.A1(n_11466),
.A2(n_9240),
.B1(n_9354),
.B2(n_9243),
.Y(n_12623)
);

AOI21xp5_ASAP7_75t_SL g12624 ( 
.A1(n_10847),
.A2(n_9354),
.B(n_9243),
.Y(n_12624)
);

OAI22xp5_ASAP7_75t_L g12625 ( 
.A1(n_11540),
.A2(n_9243),
.B1(n_9583),
.B2(n_9354),
.Y(n_12625)
);

OA21x2_ASAP7_75t_L g12626 ( 
.A1(n_10677),
.A2(n_9649),
.B(n_10087),
.Y(n_12626)
);

AND2x2_ASAP7_75t_L g12627 ( 
.A(n_10323),
.B(n_8038),
.Y(n_12627)
);

AND2x2_ASAP7_75t_L g12628 ( 
.A(n_10323),
.B(n_8063),
.Y(n_12628)
);

O2A1O1Ixp33_ASAP7_75t_L g12629 ( 
.A1(n_11546),
.A2(n_9115),
.B(n_9927),
.C(n_9554),
.Y(n_12629)
);

A2O1A1Ixp33_ASAP7_75t_L g12630 ( 
.A1(n_10676),
.A2(n_9665),
.B(n_9488),
.C(n_9475),
.Y(n_12630)
);

O2A1O1Ixp33_ASAP7_75t_L g12631 ( 
.A1(n_10358),
.A2(n_9927),
.B(n_9554),
.C(n_9937),
.Y(n_12631)
);

INVx1_ASAP7_75t_L g12632 ( 
.A(n_10565),
.Y(n_12632)
);

AOI21xp5_ASAP7_75t_SL g12633 ( 
.A1(n_10854),
.A2(n_9354),
.B(n_9243),
.Y(n_12633)
);

CKINVDCx20_ASAP7_75t_R g12634 ( 
.A(n_11460),
.Y(n_12634)
);

A2O1A1Ixp33_ASAP7_75t_L g12635 ( 
.A1(n_10681),
.A2(n_10902),
.B(n_10724),
.C(n_11141),
.Y(n_12635)
);

AND2x2_ASAP7_75t_L g12636 ( 
.A(n_10333),
.B(n_8063),
.Y(n_12636)
);

AOI21xp5_ASAP7_75t_L g12637 ( 
.A1(n_10237),
.A2(n_9937),
.B(n_9385),
.Y(n_12637)
);

AOI21x1_ASAP7_75t_SL g12638 ( 
.A1(n_11316),
.A2(n_9721),
.B(n_9720),
.Y(n_12638)
);

AOI21xp5_ASAP7_75t_L g12639 ( 
.A1(n_10477),
.A2(n_9937),
.B(n_9385),
.Y(n_12639)
);

HB1xp67_ASAP7_75t_L g12640 ( 
.A(n_10456),
.Y(n_12640)
);

AND2x2_ASAP7_75t_L g12641 ( 
.A(n_10333),
.B(n_8063),
.Y(n_12641)
);

INVx3_ASAP7_75t_L g12642 ( 
.A(n_10619),
.Y(n_12642)
);

O2A1O1Ixp33_ASAP7_75t_L g12643 ( 
.A1(n_10358),
.A2(n_9927),
.B(n_9554),
.C(n_9905),
.Y(n_12643)
);

CKINVDCx11_ASAP7_75t_R g12644 ( 
.A(n_11203),
.Y(n_12644)
);

INVx2_ASAP7_75t_L g12645 ( 
.A(n_10540),
.Y(n_12645)
);

INVx1_ASAP7_75t_SL g12646 ( 
.A(n_11460),
.Y(n_12646)
);

AOI21x1_ASAP7_75t_SL g12647 ( 
.A1(n_11403),
.A2(n_9359),
.B(n_9341),
.Y(n_12647)
);

INVx3_ASAP7_75t_L g12648 ( 
.A(n_10619),
.Y(n_12648)
);

NOR2xp33_ASAP7_75t_L g12649 ( 
.A(n_10817),
.B(n_9660),
.Y(n_12649)
);

AOI21xp5_ASAP7_75t_SL g12650 ( 
.A1(n_10854),
.A2(n_11077),
.B(n_10992),
.Y(n_12650)
);

NOR2xp67_ASAP7_75t_L g12651 ( 
.A(n_11268),
.B(n_10333),
.Y(n_12651)
);

OR2x2_ASAP7_75t_L g12652 ( 
.A(n_11620),
.B(n_8120),
.Y(n_12652)
);

OR2x2_ASAP7_75t_L g12653 ( 
.A(n_11620),
.B(n_10021),
.Y(n_12653)
);

INVx2_ASAP7_75t_L g12654 ( 
.A(n_11565),
.Y(n_12654)
);

INVx5_ASAP7_75t_L g12655 ( 
.A(n_10734),
.Y(n_12655)
);

AND2x2_ASAP7_75t_L g12656 ( 
.A(n_10333),
.B(n_8063),
.Y(n_12656)
);

AOI21x1_ASAP7_75t_SL g12657 ( 
.A1(n_11241),
.A2(n_9359),
.B(n_9341),
.Y(n_12657)
);

AND2x2_ASAP7_75t_L g12658 ( 
.A(n_10333),
.B(n_10337),
.Y(n_12658)
);

OAI22xp5_ASAP7_75t_L g12659 ( 
.A1(n_11540),
.A2(n_9243),
.B1(n_9583),
.B2(n_9354),
.Y(n_12659)
);

AOI21xp5_ASAP7_75t_L g12660 ( 
.A1(n_10477),
.A2(n_9385),
.B(n_8225),
.Y(n_12660)
);

A2O1A1Ixp33_ASAP7_75t_L g12661 ( 
.A1(n_10681),
.A2(n_9665),
.B(n_9488),
.C(n_9475),
.Y(n_12661)
);

AOI21x1_ASAP7_75t_SL g12662 ( 
.A1(n_11241),
.A2(n_9359),
.B(n_9341),
.Y(n_12662)
);

BUFx2_ASAP7_75t_L g12663 ( 
.A(n_10271),
.Y(n_12663)
);

HB1xp67_ASAP7_75t_L g12664 ( 
.A(n_10456),
.Y(n_12664)
);

INVx2_ASAP7_75t_L g12665 ( 
.A(n_11565),
.Y(n_12665)
);

A2O1A1Ixp33_ASAP7_75t_SL g12666 ( 
.A1(n_10285),
.A2(n_8611),
.B(n_8151),
.C(n_8191),
.Y(n_12666)
);

NOR2xp67_ASAP7_75t_L g12667 ( 
.A(n_10337),
.B(n_10373),
.Y(n_12667)
);

OAI22xp5_ASAP7_75t_L g12668 ( 
.A1(n_11557),
.A2(n_9354),
.B1(n_9592),
.B2(n_9583),
.Y(n_12668)
);

INVx1_ASAP7_75t_L g12669 ( 
.A(n_10584),
.Y(n_12669)
);

NOR2x1_ASAP7_75t_SL g12670 ( 
.A(n_10626),
.B(n_9574),
.Y(n_12670)
);

INVx3_ASAP7_75t_L g12671 ( 
.A(n_10619),
.Y(n_12671)
);

AOI21xp5_ASAP7_75t_L g12672 ( 
.A1(n_10582),
.A2(n_9385),
.B(n_8225),
.Y(n_12672)
);

INVx1_ASAP7_75t_L g12673 ( 
.A(n_10584),
.Y(n_12673)
);

AOI21xp5_ASAP7_75t_SL g12674 ( 
.A1(n_10854),
.A2(n_9583),
.B(n_9354),
.Y(n_12674)
);

OAI22xp5_ASAP7_75t_L g12675 ( 
.A1(n_11557),
.A2(n_9583),
.B1(n_9614),
.B2(n_9592),
.Y(n_12675)
);

INVx2_ASAP7_75t_L g12676 ( 
.A(n_11565),
.Y(n_12676)
);

INVx1_ASAP7_75t_L g12677 ( 
.A(n_10594),
.Y(n_12677)
);

OAI22xp5_ASAP7_75t_L g12678 ( 
.A1(n_11430),
.A2(n_9583),
.B1(n_9614),
.B2(n_9592),
.Y(n_12678)
);

AOI21x1_ASAP7_75t_SL g12679 ( 
.A1(n_11250),
.A2(n_9418),
.B(n_9394),
.Y(n_12679)
);

OAI22xp5_ASAP7_75t_L g12680 ( 
.A1(n_11430),
.A2(n_9583),
.B1(n_9614),
.B2(n_9592),
.Y(n_12680)
);

AND2x2_ASAP7_75t_L g12681 ( 
.A(n_10337),
.B(n_8063),
.Y(n_12681)
);

INVx2_ASAP7_75t_L g12682 ( 
.A(n_11565),
.Y(n_12682)
);

OA21x2_ASAP7_75t_L g12683 ( 
.A1(n_10630),
.A2(n_9649),
.B(n_10087),
.Y(n_12683)
);

AND2x2_ASAP7_75t_SL g12684 ( 
.A(n_10734),
.B(n_9775),
.Y(n_12684)
);

O2A1O1Ixp33_ASAP7_75t_L g12685 ( 
.A1(n_11526),
.A2(n_10715),
.B(n_10698),
.C(n_10890),
.Y(n_12685)
);

INVxp67_ASAP7_75t_SL g12686 ( 
.A(n_11258),
.Y(n_12686)
);

AOI21x1_ASAP7_75t_SL g12687 ( 
.A1(n_11250),
.A2(n_9418),
.B(n_9394),
.Y(n_12687)
);

BUFx12f_ASAP7_75t_L g12688 ( 
.A(n_11203),
.Y(n_12688)
);

AND2x2_ASAP7_75t_L g12689 ( 
.A(n_10337),
.B(n_8063),
.Y(n_12689)
);

AOI21xp5_ASAP7_75t_L g12690 ( 
.A1(n_10582),
.A2(n_10344),
.B(n_11141),
.Y(n_12690)
);

HB1xp67_ASAP7_75t_L g12691 ( 
.A(n_11588),
.Y(n_12691)
);

OAI22xp5_ASAP7_75t_L g12692 ( 
.A1(n_11376),
.A2(n_9583),
.B1(n_9614),
.B2(n_9592),
.Y(n_12692)
);

NAND2xp5_ASAP7_75t_L g12693 ( 
.A(n_11472),
.B(n_8127),
.Y(n_12693)
);

AOI21x1_ASAP7_75t_SL g12694 ( 
.A1(n_11628),
.A2(n_9418),
.B(n_9394),
.Y(n_12694)
);

BUFx12f_ASAP7_75t_L g12695 ( 
.A(n_11235),
.Y(n_12695)
);

AND2x2_ASAP7_75t_L g12696 ( 
.A(n_10337),
.B(n_8694),
.Y(n_12696)
);

NAND2xp5_ASAP7_75t_L g12697 ( 
.A(n_11472),
.B(n_8136),
.Y(n_12697)
);

INVx4_ASAP7_75t_L g12698 ( 
.A(n_11280),
.Y(n_12698)
);

AOI21xp5_ASAP7_75t_L g12699 ( 
.A1(n_10344),
.A2(n_10332),
.B(n_10298),
.Y(n_12699)
);

O2A1O1Ixp33_ASAP7_75t_L g12700 ( 
.A1(n_10698),
.A2(n_9927),
.B(n_9905),
.C(n_9923),
.Y(n_12700)
);

NAND2xp5_ASAP7_75t_L g12701 ( 
.A(n_11512),
.B(n_8136),
.Y(n_12701)
);

AND2x2_ASAP7_75t_L g12702 ( 
.A(n_10373),
.B(n_10387),
.Y(n_12702)
);

AND2x2_ASAP7_75t_L g12703 ( 
.A(n_10373),
.B(n_8694),
.Y(n_12703)
);

NAND2xp5_ASAP7_75t_L g12704 ( 
.A(n_11512),
.B(n_8646),
.Y(n_12704)
);

O2A1O1Ixp33_ASAP7_75t_L g12705 ( 
.A1(n_10698),
.A2(n_9927),
.B(n_9905),
.C(n_9923),
.Y(n_12705)
);

AOI21xp5_ASAP7_75t_SL g12706 ( 
.A1(n_10854),
.A2(n_9614),
.B(n_9592),
.Y(n_12706)
);

OA21x2_ASAP7_75t_L g12707 ( 
.A1(n_10630),
.A2(n_9649),
.B(n_10087),
.Y(n_12707)
);

INVx1_ASAP7_75t_L g12708 ( 
.A(n_10594),
.Y(n_12708)
);

A2O1A1Ixp33_ASAP7_75t_L g12709 ( 
.A1(n_10724),
.A2(n_9475),
.B(n_9531),
.C(n_9031),
.Y(n_12709)
);

O2A1O1Ixp5_ASAP7_75t_L g12710 ( 
.A1(n_11613),
.A2(n_9592),
.B(n_9670),
.C(n_9614),
.Y(n_12710)
);

O2A1O1Ixp33_ASAP7_75t_L g12711 ( 
.A1(n_10698),
.A2(n_9927),
.B(n_9923),
.C(n_9856),
.Y(n_12711)
);

AOI21xp5_ASAP7_75t_SL g12712 ( 
.A1(n_10992),
.A2(n_9614),
.B(n_9592),
.Y(n_12712)
);

INVx2_ASAP7_75t_L g12713 ( 
.A(n_11565),
.Y(n_12713)
);

OAI22xp5_ASAP7_75t_L g12714 ( 
.A1(n_11376),
.A2(n_9670),
.B1(n_9683),
.B2(n_9614),
.Y(n_12714)
);

AOI21xp5_ASAP7_75t_L g12715 ( 
.A1(n_10344),
.A2(n_10332),
.B(n_10298),
.Y(n_12715)
);

O2A1O1Ixp33_ASAP7_75t_L g12716 ( 
.A1(n_10715),
.A2(n_10891),
.B(n_10890),
.C(n_11428),
.Y(n_12716)
);

AND2x2_ASAP7_75t_L g12717 ( 
.A(n_10373),
.B(n_8694),
.Y(n_12717)
);

INVx2_ASAP7_75t_SL g12718 ( 
.A(n_11246),
.Y(n_12718)
);

NOR2x1_ASAP7_75t_SL g12719 ( 
.A(n_10626),
.B(n_9574),
.Y(n_12719)
);

NAND2xp5_ASAP7_75t_L g12720 ( 
.A(n_11567),
.B(n_8646),
.Y(n_12720)
);

AND2x2_ASAP7_75t_L g12721 ( 
.A(n_10373),
.B(n_8694),
.Y(n_12721)
);

CKINVDCx5p33_ASAP7_75t_R g12722 ( 
.A(n_10884),
.Y(n_12722)
);

OAI22xp5_ASAP7_75t_L g12723 ( 
.A1(n_10902),
.A2(n_9683),
.B1(n_9724),
.B2(n_9670),
.Y(n_12723)
);

INVx1_ASAP7_75t_L g12724 ( 
.A(n_10595),
.Y(n_12724)
);

OA21x2_ASAP7_75t_L g12725 ( 
.A1(n_10630),
.A2(n_9649),
.B(n_10087),
.Y(n_12725)
);

OAI22xp5_ASAP7_75t_L g12726 ( 
.A1(n_11334),
.A2(n_9683),
.B1(n_9724),
.B2(n_9670),
.Y(n_12726)
);

AND2x2_ASAP7_75t_L g12727 ( 
.A(n_10387),
.B(n_8880),
.Y(n_12727)
);

AND2x2_ASAP7_75t_L g12728 ( 
.A(n_10387),
.B(n_8880),
.Y(n_12728)
);

AND2x2_ASAP7_75t_L g12729 ( 
.A(n_10387),
.B(n_10442),
.Y(n_12729)
);

OA21x2_ASAP7_75t_L g12730 ( 
.A1(n_10645),
.A2(n_9649),
.B(n_10087),
.Y(n_12730)
);

INVx1_ASAP7_75t_L g12731 ( 
.A(n_10595),
.Y(n_12731)
);

OAI22xp5_ASAP7_75t_L g12732 ( 
.A1(n_10715),
.A2(n_9683),
.B1(n_9724),
.B2(n_9670),
.Y(n_12732)
);

INVx1_ASAP7_75t_L g12733 ( 
.A(n_10601),
.Y(n_12733)
);

CKINVDCx5p33_ASAP7_75t_R g12734 ( 
.A(n_11229),
.Y(n_12734)
);

NAND2xp5_ASAP7_75t_L g12735 ( 
.A(n_11567),
.B(n_8667),
.Y(n_12735)
);

NAND2xp5_ASAP7_75t_L g12736 ( 
.A(n_11428),
.B(n_8667),
.Y(n_12736)
);

NOR2xp33_ASAP7_75t_L g12737 ( 
.A(n_11437),
.B(n_9660),
.Y(n_12737)
);

AND2x2_ASAP7_75t_L g12738 ( 
.A(n_10387),
.B(n_8880),
.Y(n_12738)
);

AND2x2_ASAP7_75t_L g12739 ( 
.A(n_10442),
.B(n_8880),
.Y(n_12739)
);

AND2x2_ASAP7_75t_L g12740 ( 
.A(n_10442),
.B(n_10482),
.Y(n_12740)
);

AND2x2_ASAP7_75t_L g12741 ( 
.A(n_10442),
.B(n_9390),
.Y(n_12741)
);

OR2x2_ASAP7_75t_L g12742 ( 
.A(n_10404),
.B(n_10021),
.Y(n_12742)
);

AOI21xp5_ASAP7_75t_L g12743 ( 
.A1(n_10344),
.A2(n_9385),
.B(n_9007),
.Y(n_12743)
);

CKINVDCx6p67_ASAP7_75t_R g12744 ( 
.A(n_10600),
.Y(n_12744)
);

OAI22xp5_ASAP7_75t_L g12745 ( 
.A1(n_10715),
.A2(n_9683),
.B1(n_9724),
.B2(n_9670),
.Y(n_12745)
);

O2A1O1Ixp33_ASAP7_75t_L g12746 ( 
.A1(n_10890),
.A2(n_9927),
.B(n_9856),
.C(n_9230),
.Y(n_12746)
);

INVx2_ASAP7_75t_L g12747 ( 
.A(n_11586),
.Y(n_12747)
);

OAI22xp5_ASAP7_75t_SL g12748 ( 
.A1(n_10728),
.A2(n_9782),
.B1(n_9669),
.B2(n_9660),
.Y(n_12748)
);

AND2x2_ASAP7_75t_L g12749 ( 
.A(n_10442),
.B(n_9390),
.Y(n_12749)
);

INVx1_ASAP7_75t_SL g12750 ( 
.A(n_11529),
.Y(n_12750)
);

AND2x2_ASAP7_75t_L g12751 ( 
.A(n_10482),
.B(n_9390),
.Y(n_12751)
);

NAND2xp5_ASAP7_75t_L g12752 ( 
.A(n_11473),
.B(n_8676),
.Y(n_12752)
);

O2A1O1Ixp5_ASAP7_75t_L g12753 ( 
.A1(n_11613),
.A2(n_9670),
.B(n_9724),
.C(n_9683),
.Y(n_12753)
);

A2O1A1Ixp33_ASAP7_75t_L g12754 ( 
.A1(n_11189),
.A2(n_9531),
.B(n_9031),
.C(n_9049),
.Y(n_12754)
);

HB1xp67_ASAP7_75t_L g12755 ( 
.A(n_11588),
.Y(n_12755)
);

INVx1_ASAP7_75t_L g12756 ( 
.A(n_10601),
.Y(n_12756)
);

HB1xp67_ASAP7_75t_L g12757 ( 
.A(n_11588),
.Y(n_12757)
);

OAI22xp5_ASAP7_75t_L g12758 ( 
.A1(n_11295),
.A2(n_11348),
.B1(n_10460),
.B2(n_10862),
.Y(n_12758)
);

NOR2xp67_ASAP7_75t_L g12759 ( 
.A(n_10482),
.B(n_9669),
.Y(n_12759)
);

OA21x2_ASAP7_75t_L g12760 ( 
.A1(n_10645),
.A2(n_9649),
.B(n_9757),
.Y(n_12760)
);

BUFx3_ASAP7_75t_L g12761 ( 
.A(n_10271),
.Y(n_12761)
);

NAND2xp5_ASAP7_75t_L g12762 ( 
.A(n_11473),
.B(n_8676),
.Y(n_12762)
);

OAI22xp5_ASAP7_75t_SL g12763 ( 
.A1(n_10644),
.A2(n_9669),
.B1(n_9782),
.B2(n_10116),
.Y(n_12763)
);

NAND2xp5_ASAP7_75t_L g12764 ( 
.A(n_11174),
.B(n_8682),
.Y(n_12764)
);

AND2x4_ASAP7_75t_L g12765 ( 
.A(n_10992),
.B(n_9390),
.Y(n_12765)
);

HB1xp67_ASAP7_75t_L g12766 ( 
.A(n_11625),
.Y(n_12766)
);

INVx1_ASAP7_75t_L g12767 ( 
.A(n_10608),
.Y(n_12767)
);

NAND2xp5_ASAP7_75t_L g12768 ( 
.A(n_11174),
.B(n_8682),
.Y(n_12768)
);

INVx2_ASAP7_75t_L g12769 ( 
.A(n_11586),
.Y(n_12769)
);

AND2x4_ASAP7_75t_L g12770 ( 
.A(n_10992),
.B(n_9396),
.Y(n_12770)
);

OA21x2_ASAP7_75t_L g12771 ( 
.A1(n_10645),
.A2(n_10653),
.B(n_11155),
.Y(n_12771)
);

OA21x2_ASAP7_75t_L g12772 ( 
.A1(n_10653),
.A2(n_9772),
.B(n_9757),
.Y(n_12772)
);

OAI22xp5_ASAP7_75t_L g12773 ( 
.A1(n_11295),
.A2(n_9683),
.B1(n_9724),
.B2(n_9670),
.Y(n_12773)
);

AND2x2_ASAP7_75t_L g12774 ( 
.A(n_10482),
.B(n_9396),
.Y(n_12774)
);

NAND2xp5_ASAP7_75t_L g12775 ( 
.A(n_11240),
.B(n_8062),
.Y(n_12775)
);

AOI21xp5_ASAP7_75t_L g12776 ( 
.A1(n_10344),
.A2(n_9007),
.B(n_9029),
.Y(n_12776)
);

INVx2_ASAP7_75t_L g12777 ( 
.A(n_11586),
.Y(n_12777)
);

OAI22xp5_ASAP7_75t_L g12778 ( 
.A1(n_11348),
.A2(n_9724),
.B1(n_9855),
.B2(n_9683),
.Y(n_12778)
);

OAI22xp5_ASAP7_75t_L g12779 ( 
.A1(n_11348),
.A2(n_9855),
.B1(n_9873),
.B2(n_9724),
.Y(n_12779)
);

OAI22xp5_ASAP7_75t_L g12780 ( 
.A1(n_10219),
.A2(n_9873),
.B1(n_9874),
.B2(n_9855),
.Y(n_12780)
);

AOI21xp5_ASAP7_75t_L g12781 ( 
.A1(n_10332),
.A2(n_10298),
.B(n_10306),
.Y(n_12781)
);

AOI21xp5_ASAP7_75t_L g12782 ( 
.A1(n_10332),
.A2(n_9031),
.B(n_9029),
.Y(n_12782)
);

INVx1_ASAP7_75t_L g12783 ( 
.A(n_10608),
.Y(n_12783)
);

OAI22xp5_ASAP7_75t_L g12784 ( 
.A1(n_10219),
.A2(n_9873),
.B1(n_9874),
.B2(n_9855),
.Y(n_12784)
);

BUFx12f_ASAP7_75t_L g12785 ( 
.A(n_11235),
.Y(n_12785)
);

AOI21x1_ASAP7_75t_SL g12786 ( 
.A1(n_11628),
.A2(n_9426),
.B(n_10021),
.Y(n_12786)
);

OR2x2_ASAP7_75t_L g12787 ( 
.A(n_10404),
.B(n_10037),
.Y(n_12787)
);

OR2x2_ASAP7_75t_L g12788 ( 
.A(n_10404),
.B(n_10037),
.Y(n_12788)
);

O2A1O1Ixp33_ASAP7_75t_L g12789 ( 
.A1(n_10891),
.A2(n_9856),
.B(n_9230),
.C(n_9244),
.Y(n_12789)
);

AND2x2_ASAP7_75t_L g12790 ( 
.A(n_10482),
.B(n_9396),
.Y(n_12790)
);

O2A1O1Ixp5_ASAP7_75t_L g12791 ( 
.A1(n_11613),
.A2(n_9873),
.B(n_9874),
.C(n_9855),
.Y(n_12791)
);

OAI22xp5_ASAP7_75t_SL g12792 ( 
.A1(n_10644),
.A2(n_9782),
.B1(n_10116),
.B2(n_8154),
.Y(n_12792)
);

AND2x2_ASAP7_75t_L g12793 ( 
.A(n_10500),
.B(n_9396),
.Y(n_12793)
);

AOI21xp5_ASAP7_75t_L g12794 ( 
.A1(n_10332),
.A2(n_9049),
.B(n_9029),
.Y(n_12794)
);

AOI21xp5_ASAP7_75t_L g12795 ( 
.A1(n_10298),
.A2(n_9049),
.B(n_9603),
.Y(n_12795)
);

OR2x2_ASAP7_75t_L g12796 ( 
.A(n_10404),
.B(n_10037),
.Y(n_12796)
);

CKINVDCx5p33_ASAP7_75t_R g12797 ( 
.A(n_11518),
.Y(n_12797)
);

AND2x4_ASAP7_75t_L g12798 ( 
.A(n_11077),
.B(n_9869),
.Y(n_12798)
);

AOI21xp5_ASAP7_75t_L g12799 ( 
.A1(n_10298),
.A2(n_10306),
.B(n_11280),
.Y(n_12799)
);

AND2x2_ASAP7_75t_L g12800 ( 
.A(n_10500),
.B(n_9396),
.Y(n_12800)
);

AO21x2_ASAP7_75t_L g12801 ( 
.A1(n_11598),
.A2(n_9976),
.B(n_9952),
.Y(n_12801)
);

BUFx4f_ASAP7_75t_SL g12802 ( 
.A(n_10435),
.Y(n_12802)
);

INVx2_ASAP7_75t_L g12803 ( 
.A(n_11586),
.Y(n_12803)
);

OAI22xp5_ASAP7_75t_L g12804 ( 
.A1(n_10219),
.A2(n_9873),
.B1(n_9874),
.B2(n_9855),
.Y(n_12804)
);

AOI21x1_ASAP7_75t_SL g12805 ( 
.A1(n_11628),
.A2(n_9426),
.B(n_9842),
.Y(n_12805)
);

AND2x2_ASAP7_75t_L g12806 ( 
.A(n_10500),
.B(n_9396),
.Y(n_12806)
);

OR2x2_ASAP7_75t_L g12807 ( 
.A(n_10404),
.B(n_8306),
.Y(n_12807)
);

BUFx6f_ASAP7_75t_L g12808 ( 
.A(n_11518),
.Y(n_12808)
);

NOR2xp67_ASAP7_75t_L g12809 ( 
.A(n_10500),
.B(n_10516),
.Y(n_12809)
);

AOI21xp5_ASAP7_75t_SL g12810 ( 
.A1(n_11077),
.A2(n_9873),
.B(n_9855),
.Y(n_12810)
);

AOI21x1_ASAP7_75t_SL g12811 ( 
.A1(n_11628),
.A2(n_9426),
.B(n_9842),
.Y(n_12811)
);

INVx1_ASAP7_75t_L g12812 ( 
.A(n_10609),
.Y(n_12812)
);

O2A1O1Ixp5_ASAP7_75t_L g12813 ( 
.A1(n_11258),
.A2(n_9855),
.B(n_9874),
.C(n_9873),
.Y(n_12813)
);

INVx2_ASAP7_75t_L g12814 ( 
.A(n_11586),
.Y(n_12814)
);

NAND2xp5_ASAP7_75t_L g12815 ( 
.A(n_11240),
.B(n_8062),
.Y(n_12815)
);

OA21x2_ASAP7_75t_L g12816 ( 
.A1(n_10653),
.A2(n_9772),
.B(n_9757),
.Y(n_12816)
);

AOI221x1_ASAP7_75t_SL g12817 ( 
.A1(n_11397),
.A2(n_9796),
.B1(n_9843),
.B2(n_9809),
.C(n_9787),
.Y(n_12817)
);

AND2x4_ASAP7_75t_L g12818 ( 
.A(n_11077),
.B(n_9869),
.Y(n_12818)
);

NOR2xp67_ASAP7_75t_L g12819 ( 
.A(n_10500),
.B(n_9782),
.Y(n_12819)
);

OAI22xp5_ASAP7_75t_L g12820 ( 
.A1(n_10219),
.A2(n_9874),
.B1(n_9989),
.B2(n_9873),
.Y(n_12820)
);

INVxp67_ASAP7_75t_L g12821 ( 
.A(n_11625),
.Y(n_12821)
);

CKINVDCx14_ASAP7_75t_R g12822 ( 
.A(n_10219),
.Y(n_12822)
);

O2A1O1Ixp33_ASAP7_75t_L g12823 ( 
.A1(n_10891),
.A2(n_11230),
.B(n_11159),
.C(n_11115),
.Y(n_12823)
);

AND2x2_ASAP7_75t_L g12824 ( 
.A(n_10516),
.B(n_9453),
.Y(n_12824)
);

INVx1_ASAP7_75t_L g12825 ( 
.A(n_10609),
.Y(n_12825)
);

INVx3_ASAP7_75t_L g12826 ( 
.A(n_10711),
.Y(n_12826)
);

BUFx6f_ASAP7_75t_L g12827 ( 
.A(n_11175),
.Y(n_12827)
);

AOI21x1_ASAP7_75t_SL g12828 ( 
.A1(n_11628),
.A2(n_9842),
.B(n_7723),
.Y(n_12828)
);

AOI21xp5_ASAP7_75t_L g12829 ( 
.A1(n_10306),
.A2(n_9611),
.B(n_9603),
.Y(n_12829)
);

BUFx2_ASAP7_75t_R g12830 ( 
.A(n_11175),
.Y(n_12830)
);

AND2x2_ASAP7_75t_L g12831 ( 
.A(n_10516),
.B(n_9453),
.Y(n_12831)
);

BUFx2_ASAP7_75t_L g12832 ( 
.A(n_10435),
.Y(n_12832)
);

OA21x2_ASAP7_75t_L g12833 ( 
.A1(n_11155),
.A2(n_9772),
.B(n_9757),
.Y(n_12833)
);

NAND2xp5_ASAP7_75t_L g12834 ( 
.A(n_11345),
.B(n_8068),
.Y(n_12834)
);

AND2x2_ASAP7_75t_L g12835 ( 
.A(n_10516),
.B(n_10689),
.Y(n_12835)
);

OA21x2_ASAP7_75t_L g12836 ( 
.A1(n_11155),
.A2(n_9778),
.B(n_9772),
.Y(n_12836)
);

INVx1_ASAP7_75t_L g12837 ( 
.A(n_10615),
.Y(n_12837)
);

OR2x2_ASAP7_75t_L g12838 ( 
.A(n_10404),
.B(n_8306),
.Y(n_12838)
);

AOI21x1_ASAP7_75t_SL g12839 ( 
.A1(n_11577),
.A2(n_7723),
.B(n_7722),
.Y(n_12839)
);

NAND2xp5_ASAP7_75t_L g12840 ( 
.A(n_11345),
.B(n_8068),
.Y(n_12840)
);

INVx2_ASAP7_75t_L g12841 ( 
.A(n_11625),
.Y(n_12841)
);

INVx1_ASAP7_75t_SL g12842 ( 
.A(n_11175),
.Y(n_12842)
);

AOI21xp5_ASAP7_75t_SL g12843 ( 
.A1(n_11273),
.A2(n_9989),
.B(n_9874),
.Y(n_12843)
);

AND2x2_ASAP7_75t_L g12844 ( 
.A(n_10516),
.B(n_9453),
.Y(n_12844)
);

NAND2xp5_ASAP7_75t_L g12845 ( 
.A(n_11401),
.B(n_7970),
.Y(n_12845)
);

AND2x4_ASAP7_75t_L g12846 ( 
.A(n_11273),
.B(n_9453),
.Y(n_12846)
);

NAND2xp5_ASAP7_75t_L g12847 ( 
.A(n_11401),
.B(n_7970),
.Y(n_12847)
);

INVx1_ASAP7_75t_L g12848 ( 
.A(n_10615),
.Y(n_12848)
);

INVx2_ASAP7_75t_L g12849 ( 
.A(n_10622),
.Y(n_12849)
);

AOI21xp5_ASAP7_75t_SL g12850 ( 
.A1(n_11273),
.A2(n_9989),
.B(n_9874),
.Y(n_12850)
);

O2A1O1Ixp5_ASAP7_75t_L g12851 ( 
.A1(n_11258),
.A2(n_10285),
.B(n_11161),
.C(n_10685),
.Y(n_12851)
);

AND2x2_ASAP7_75t_L g12852 ( 
.A(n_10689),
.B(n_9453),
.Y(n_12852)
);

INVx1_ASAP7_75t_SL g12853 ( 
.A(n_11175),
.Y(n_12853)
);

AND2x2_ASAP7_75t_L g12854 ( 
.A(n_10689),
.B(n_9453),
.Y(n_12854)
);

INVx1_ASAP7_75t_L g12855 ( 
.A(n_10622),
.Y(n_12855)
);

AND2x2_ASAP7_75t_L g12856 ( 
.A(n_10689),
.B(n_9460),
.Y(n_12856)
);

HB1xp67_ASAP7_75t_L g12857 ( 
.A(n_10464),
.Y(n_12857)
);

AOI21xp5_ASAP7_75t_L g12858 ( 
.A1(n_10306),
.A2(n_9611),
.B(n_9603),
.Y(n_12858)
);

NAND2xp5_ASAP7_75t_L g12859 ( 
.A(n_11412),
.B(n_7976),
.Y(n_12859)
);

AOI21xp5_ASAP7_75t_SL g12860 ( 
.A1(n_11273),
.A2(n_10012),
.B(n_9989),
.Y(n_12860)
);

NAND2xp5_ASAP7_75t_L g12861 ( 
.A(n_11412),
.B(n_7976),
.Y(n_12861)
);

A2O1A1Ixp33_ASAP7_75t_L g12862 ( 
.A1(n_11189),
.A2(n_11197),
.B(n_11278),
.C(n_11272),
.Y(n_12862)
);

AOI21xp5_ASAP7_75t_L g12863 ( 
.A1(n_10306),
.A2(n_9611),
.B(n_9756),
.Y(n_12863)
);

AND2x2_ASAP7_75t_L g12864 ( 
.A(n_10689),
.B(n_9460),
.Y(n_12864)
);

O2A1O1Ixp33_ASAP7_75t_L g12865 ( 
.A1(n_11230),
.A2(n_9230),
.B(n_9244),
.C(n_9231),
.Y(n_12865)
);

O2A1O1Ixp33_ASAP7_75t_L g12866 ( 
.A1(n_11230),
.A2(n_9230),
.B(n_9244),
.C(n_9231),
.Y(n_12866)
);

NAND2xp5_ASAP7_75t_L g12867 ( 
.A(n_10227),
.B(n_7980),
.Y(n_12867)
);

INVx1_ASAP7_75t_L g12868 ( 
.A(n_10640),
.Y(n_12868)
);

AND2x4_ASAP7_75t_L g12869 ( 
.A(n_11576),
.B(n_9460),
.Y(n_12869)
);

AND2x2_ASAP7_75t_L g12870 ( 
.A(n_10725),
.B(n_10779),
.Y(n_12870)
);

O2A1O1Ixp33_ASAP7_75t_L g12871 ( 
.A1(n_11115),
.A2(n_11159),
.B(n_10278),
.C(n_10364),
.Y(n_12871)
);

AOI21xp5_ASAP7_75t_SL g12872 ( 
.A1(n_10734),
.A2(n_10012),
.B(n_9989),
.Y(n_12872)
);

O2A1O1Ixp33_ASAP7_75t_L g12873 ( 
.A1(n_11115),
.A2(n_9230),
.B(n_9244),
.C(n_9231),
.Y(n_12873)
);

AOI21xp5_ASAP7_75t_L g12874 ( 
.A1(n_11280),
.A2(n_10027),
.B(n_9756),
.Y(n_12874)
);

AND2x2_ASAP7_75t_L g12875 ( 
.A(n_10725),
.B(n_9460),
.Y(n_12875)
);

BUFx12f_ASAP7_75t_L g12876 ( 
.A(n_10435),
.Y(n_12876)
);

AND2x4_ASAP7_75t_L g12877 ( 
.A(n_11576),
.B(n_9460),
.Y(n_12877)
);

OR2x2_ASAP7_75t_L g12878 ( 
.A(n_10404),
.B(n_8306),
.Y(n_12878)
);

INVx2_ASAP7_75t_L g12879 ( 
.A(n_10640),
.Y(n_12879)
);

A2O1A1Ixp33_ASAP7_75t_L g12880 ( 
.A1(n_11197),
.A2(n_11278),
.B(n_11272),
.C(n_11285),
.Y(n_12880)
);

OAI22xp5_ASAP7_75t_L g12881 ( 
.A1(n_10219),
.A2(n_10012),
.B1(n_10049),
.B2(n_9989),
.Y(n_12881)
);

AND2x2_ASAP7_75t_SL g12882 ( 
.A(n_10867),
.B(n_9775),
.Y(n_12882)
);

AOI211xp5_ASAP7_75t_L g12883 ( 
.A1(n_11491),
.A2(n_9231),
.B(n_9308),
.C(n_9244),
.Y(n_12883)
);

INVx4_ASAP7_75t_L g12884 ( 
.A(n_11280),
.Y(n_12884)
);

AND2x2_ASAP7_75t_L g12885 ( 
.A(n_10725),
.B(n_9460),
.Y(n_12885)
);

INVx2_ASAP7_75t_L g12886 ( 
.A(n_10649),
.Y(n_12886)
);

OA21x2_ASAP7_75t_L g12887 ( 
.A1(n_11155),
.A2(n_9779),
.B(n_9778),
.Y(n_12887)
);

AND2x2_ASAP7_75t_L g12888 ( 
.A(n_10725),
.B(n_9461),
.Y(n_12888)
);

NAND2xp5_ASAP7_75t_L g12889 ( 
.A(n_10227),
.B(n_7980),
.Y(n_12889)
);

OAI22xp5_ASAP7_75t_L g12890 ( 
.A1(n_10460),
.A2(n_10012),
.B1(n_10049),
.B2(n_9989),
.Y(n_12890)
);

CKINVDCx5p33_ASAP7_75t_R g12891 ( 
.A(n_10435),
.Y(n_12891)
);

AOI21xp5_ASAP7_75t_L g12892 ( 
.A1(n_11285),
.A2(n_11292),
.B(n_11491),
.Y(n_12892)
);

INVx2_ASAP7_75t_L g12893 ( 
.A(n_10649),
.Y(n_12893)
);

AOI22xp5_ASAP7_75t_L g12894 ( 
.A1(n_11005),
.A2(n_8513),
.B1(n_9349),
.B2(n_8454),
.Y(n_12894)
);

AND2x2_ASAP7_75t_L g12895 ( 
.A(n_10725),
.B(n_9461),
.Y(n_12895)
);

NAND2xp5_ASAP7_75t_L g12896 ( 
.A(n_10227),
.B(n_7981),
.Y(n_12896)
);

AOI21x1_ASAP7_75t_SL g12897 ( 
.A1(n_11577),
.A2(n_7731),
.B(n_7722),
.Y(n_12897)
);

INVxp67_ASAP7_75t_L g12898 ( 
.A(n_10808),
.Y(n_12898)
);

INVx1_ASAP7_75t_L g12899 ( 
.A(n_10656),
.Y(n_12899)
);

INVxp67_ASAP7_75t_L g12900 ( 
.A(n_10808),
.Y(n_12900)
);

AND2x2_ASAP7_75t_L g12901 ( 
.A(n_10779),
.B(n_9461),
.Y(n_12901)
);

OR2x2_ASAP7_75t_L g12902 ( 
.A(n_10404),
.B(n_9512),
.Y(n_12902)
);

INVx1_ASAP7_75t_L g12903 ( 
.A(n_10656),
.Y(n_12903)
);

AOI21xp5_ASAP7_75t_SL g12904 ( 
.A1(n_10867),
.A2(n_10012),
.B(n_9989),
.Y(n_12904)
);

OR2x2_ASAP7_75t_L g12905 ( 
.A(n_10965),
.B(n_9512),
.Y(n_12905)
);

INVx1_ASAP7_75t_L g12906 ( 
.A(n_10662),
.Y(n_12906)
);

INVx2_ASAP7_75t_L g12907 ( 
.A(n_10662),
.Y(n_12907)
);

AO21x2_ASAP7_75t_L g12908 ( 
.A1(n_12384),
.A2(n_11161),
.B(n_10685),
.Y(n_12908)
);

OAI21xp5_ASAP7_75t_L g12909 ( 
.A1(n_11642),
.A2(n_11600),
.B(n_11558),
.Y(n_12909)
);

OR2x2_ASAP7_75t_L g12910 ( 
.A(n_11987),
.B(n_9512),
.Y(n_12910)
);

INVx2_ASAP7_75t_L g12911 ( 
.A(n_11794),
.Y(n_12911)
);

INVx1_ASAP7_75t_L g12912 ( 
.A(n_11657),
.Y(n_12912)
);

OR2x2_ASAP7_75t_L g12913 ( 
.A(n_11771),
.B(n_9512),
.Y(n_12913)
);

INVx1_ASAP7_75t_L g12914 ( 
.A(n_11657),
.Y(n_12914)
);

INVx1_ASAP7_75t_L g12915 ( 
.A(n_11658),
.Y(n_12915)
);

INVx3_ASAP7_75t_L g12916 ( 
.A(n_11954),
.Y(n_12916)
);

AOI21x1_ASAP7_75t_L g12917 ( 
.A1(n_12155),
.A2(n_11100),
.B(n_10666),
.Y(n_12917)
);

INVx3_ASAP7_75t_L g12918 ( 
.A(n_11954),
.Y(n_12918)
);

OA21x2_ASAP7_75t_L g12919 ( 
.A1(n_11865),
.A2(n_11191),
.B(n_11156),
.Y(n_12919)
);

INVx1_ASAP7_75t_L g12920 ( 
.A(n_11658),
.Y(n_12920)
);

HB1xp67_ASAP7_75t_L g12921 ( 
.A(n_11746),
.Y(n_12921)
);

INVx2_ASAP7_75t_L g12922 ( 
.A(n_11794),
.Y(n_12922)
);

AND2x2_ASAP7_75t_L g12923 ( 
.A(n_12284),
.B(n_10867),
.Y(n_12923)
);

INVx3_ASAP7_75t_L g12924 ( 
.A(n_11975),
.Y(n_12924)
);

INVx1_ASAP7_75t_L g12925 ( 
.A(n_11667),
.Y(n_12925)
);

INVx1_ASAP7_75t_L g12926 ( 
.A(n_11667),
.Y(n_12926)
);

AOI22xp33_ASAP7_75t_L g12927 ( 
.A1(n_12206),
.A2(n_11005),
.B1(n_10388),
.B2(n_10383),
.Y(n_12927)
);

OR2x6_ASAP7_75t_L g12928 ( 
.A(n_12650),
.B(n_10867),
.Y(n_12928)
);

INVx2_ASAP7_75t_L g12929 ( 
.A(n_11967),
.Y(n_12929)
);

INVx2_ASAP7_75t_L g12930 ( 
.A(n_11967),
.Y(n_12930)
);

INVx2_ASAP7_75t_L g12931 ( 
.A(n_12002),
.Y(n_12931)
);

AOI21x1_ASAP7_75t_L g12932 ( 
.A1(n_12155),
.A2(n_10666),
.B(n_10637),
.Y(n_12932)
);

OA21x2_ASAP7_75t_L g12933 ( 
.A1(n_11865),
.A2(n_11191),
.B(n_11156),
.Y(n_12933)
);

HB1xp67_ASAP7_75t_L g12934 ( 
.A(n_11746),
.Y(n_12934)
);

INVx2_ASAP7_75t_L g12935 ( 
.A(n_12002),
.Y(n_12935)
);

INVx3_ASAP7_75t_L g12936 ( 
.A(n_11975),
.Y(n_12936)
);

HB1xp67_ASAP7_75t_L g12937 ( 
.A(n_11746),
.Y(n_12937)
);

INVx5_ASAP7_75t_SL g12938 ( 
.A(n_11887),
.Y(n_12938)
);

INVx2_ASAP7_75t_SL g12939 ( 
.A(n_11933),
.Y(n_12939)
);

BUFx6f_ASAP7_75t_L g12940 ( 
.A(n_12149),
.Y(n_12940)
);

BUFx3_ASAP7_75t_L g12941 ( 
.A(n_12500),
.Y(n_12941)
);

INVx2_ASAP7_75t_SL g12942 ( 
.A(n_11933),
.Y(n_12942)
);

AND2x2_ASAP7_75t_L g12943 ( 
.A(n_12120),
.B(n_10867),
.Y(n_12943)
);

INVx1_ASAP7_75t_L g12944 ( 
.A(n_11675),
.Y(n_12944)
);

OA21x2_ASAP7_75t_L g12945 ( 
.A1(n_12074),
.A2(n_12686),
.B(n_12416),
.Y(n_12945)
);

BUFx2_ASAP7_75t_L g12946 ( 
.A(n_12196),
.Y(n_12946)
);

NAND2xp5_ASAP7_75t_SL g12947 ( 
.A(n_12407),
.B(n_10970),
.Y(n_12947)
);

INVx2_ASAP7_75t_L g12948 ( 
.A(n_12008),
.Y(n_12948)
);

OAI21x1_ASAP7_75t_SL g12949 ( 
.A1(n_11724),
.A2(n_12328),
.B(n_12622),
.Y(n_12949)
);

HB1xp67_ASAP7_75t_L g12950 ( 
.A(n_12691),
.Y(n_12950)
);

INVx1_ASAP7_75t_L g12951 ( 
.A(n_11675),
.Y(n_12951)
);

AO21x2_ASAP7_75t_L g12952 ( 
.A1(n_12686),
.A2(n_11598),
.B(n_10999),
.Y(n_12952)
);

INVx1_ASAP7_75t_L g12953 ( 
.A(n_11709),
.Y(n_12953)
);

INVx1_ASAP7_75t_L g12954 ( 
.A(n_11709),
.Y(n_12954)
);

OA21x2_ASAP7_75t_L g12955 ( 
.A1(n_12074),
.A2(n_11191),
.B(n_11156),
.Y(n_12955)
);

NOR2x1_ASAP7_75t_R g12956 ( 
.A(n_11799),
.B(n_9782),
.Y(n_12956)
);

INVx1_ASAP7_75t_L g12957 ( 
.A(n_11716),
.Y(n_12957)
);

HB1xp67_ASAP7_75t_L g12958 ( 
.A(n_12691),
.Y(n_12958)
);

INVx1_ASAP7_75t_L g12959 ( 
.A(n_11716),
.Y(n_12959)
);

AND2x2_ASAP7_75t_L g12960 ( 
.A(n_12121),
.B(n_10970),
.Y(n_12960)
);

AO21x1_ASAP7_75t_SL g12961 ( 
.A1(n_12243),
.A2(n_10355),
.B(n_10278),
.Y(n_12961)
);

BUFx3_ASAP7_75t_L g12962 ( 
.A(n_12500),
.Y(n_12962)
);

OR2x2_ASAP7_75t_L g12963 ( 
.A(n_11772),
.B(n_9512),
.Y(n_12963)
);

INVx1_ASAP7_75t_SL g12964 ( 
.A(n_12078),
.Y(n_12964)
);

HB1xp67_ASAP7_75t_L g12965 ( 
.A(n_12755),
.Y(n_12965)
);

BUFx4f_ASAP7_75t_SL g12966 ( 
.A(n_12196),
.Y(n_12966)
);

BUFx2_ASAP7_75t_L g12967 ( 
.A(n_12688),
.Y(n_12967)
);

INVx1_ASAP7_75t_L g12968 ( 
.A(n_11753),
.Y(n_12968)
);

NAND2xp5_ASAP7_75t_L g12969 ( 
.A(n_11683),
.B(n_9641),
.Y(n_12969)
);

HB1xp67_ASAP7_75t_L g12970 ( 
.A(n_12755),
.Y(n_12970)
);

INVx1_ASAP7_75t_L g12971 ( 
.A(n_11753),
.Y(n_12971)
);

INVxp67_ASAP7_75t_L g12972 ( 
.A(n_11818),
.Y(n_12972)
);

INVx1_ASAP7_75t_L g12973 ( 
.A(n_11790),
.Y(n_12973)
);

NAND2xp5_ASAP7_75t_L g12974 ( 
.A(n_12199),
.B(n_9641),
.Y(n_12974)
);

INVx1_ASAP7_75t_L g12975 ( 
.A(n_11790),
.Y(n_12975)
);

HB1xp67_ASAP7_75t_L g12976 ( 
.A(n_12757),
.Y(n_12976)
);

BUFx6f_ASAP7_75t_L g12977 ( 
.A(n_12149),
.Y(n_12977)
);

BUFx3_ASAP7_75t_L g12978 ( 
.A(n_12688),
.Y(n_12978)
);

AND2x2_ASAP7_75t_L g12979 ( 
.A(n_11804),
.B(n_10970),
.Y(n_12979)
);

AND2x4_ASAP7_75t_L g12980 ( 
.A(n_12273),
.B(n_10970),
.Y(n_12980)
);

OAI21x1_ASAP7_75t_L g12981 ( 
.A1(n_12416),
.A2(n_10419),
.B(n_11159),
.Y(n_12981)
);

OR2x2_ASAP7_75t_L g12982 ( 
.A(n_12004),
.B(n_9512),
.Y(n_12982)
);

OR2x2_ASAP7_75t_L g12983 ( 
.A(n_11935),
.B(n_9512),
.Y(n_12983)
);

OAI21x1_ASAP7_75t_L g12984 ( 
.A1(n_12189),
.A2(n_10419),
.B(n_10417),
.Y(n_12984)
);

BUFx2_ASAP7_75t_L g12985 ( 
.A(n_12695),
.Y(n_12985)
);

AND2x4_ASAP7_75t_L g12986 ( 
.A(n_12420),
.B(n_10970),
.Y(n_12986)
);

BUFx3_ASAP7_75t_L g12987 ( 
.A(n_11713),
.Y(n_12987)
);

OAI21x1_ASAP7_75t_L g12988 ( 
.A1(n_12189),
.A2(n_10419),
.B(n_10417),
.Y(n_12988)
);

INVx2_ASAP7_75t_L g12989 ( 
.A(n_12008),
.Y(n_12989)
);

INVx2_ASAP7_75t_L g12990 ( 
.A(n_12065),
.Y(n_12990)
);

INVx1_ASAP7_75t_L g12991 ( 
.A(n_11815),
.Y(n_12991)
);

AND2x2_ASAP7_75t_L g12992 ( 
.A(n_12551),
.B(n_11135),
.Y(n_12992)
);

AO21x2_ASAP7_75t_L g12993 ( 
.A1(n_12095),
.A2(n_11598),
.B(n_10999),
.Y(n_12993)
);

INVx2_ASAP7_75t_L g12994 ( 
.A(n_12065),
.Y(n_12994)
);

AND2x4_ASAP7_75t_L g12995 ( 
.A(n_12420),
.B(n_11135),
.Y(n_12995)
);

HB1xp67_ASAP7_75t_L g12996 ( 
.A(n_12757),
.Y(n_12996)
);

INVx1_ASAP7_75t_L g12997 ( 
.A(n_11815),
.Y(n_12997)
);

INVx2_ASAP7_75t_L g12998 ( 
.A(n_12569),
.Y(n_12998)
);

INVx1_ASAP7_75t_L g12999 ( 
.A(n_11637),
.Y(n_12999)
);

INVx2_ASAP7_75t_L g13000 ( 
.A(n_12569),
.Y(n_13000)
);

HB1xp67_ASAP7_75t_L g13001 ( 
.A(n_12766),
.Y(n_13001)
);

INVx2_ASAP7_75t_L g13002 ( 
.A(n_11788),
.Y(n_13002)
);

AO31x2_ASAP7_75t_L g13003 ( 
.A1(n_11858),
.A2(n_11443),
.A3(n_11234),
.B(n_11393),
.Y(n_13003)
);

INVx1_ASAP7_75t_L g13004 ( 
.A(n_11637),
.Y(n_13004)
);

OAI21x1_ASAP7_75t_L g13005 ( 
.A1(n_12306),
.A2(n_10417),
.B(n_11164),
.Y(n_13005)
);

INVx1_ASAP7_75t_L g13006 ( 
.A(n_12570),
.Y(n_13006)
);

BUFx2_ASAP7_75t_L g13007 ( 
.A(n_12695),
.Y(n_13007)
);

HB1xp67_ASAP7_75t_L g13008 ( 
.A(n_12766),
.Y(n_13008)
);

INVx2_ASAP7_75t_L g13009 ( 
.A(n_11973),
.Y(n_13009)
);

INVx1_ASAP7_75t_L g13010 ( 
.A(n_12570),
.Y(n_13010)
);

INVx2_ASAP7_75t_L g13011 ( 
.A(n_11982),
.Y(n_13011)
);

NAND2xp5_ASAP7_75t_SL g13012 ( 
.A(n_12415),
.B(n_11135),
.Y(n_13012)
);

INVx2_ASAP7_75t_SL g13013 ( 
.A(n_11650),
.Y(n_13013)
);

AND2x2_ASAP7_75t_L g13014 ( 
.A(n_12551),
.B(n_11991),
.Y(n_13014)
);

HB1xp67_ASAP7_75t_L g13015 ( 
.A(n_12092),
.Y(n_13015)
);

OR2x2_ASAP7_75t_L g13016 ( 
.A(n_11937),
.B(n_9512),
.Y(n_13016)
);

AND2x2_ASAP7_75t_L g13017 ( 
.A(n_11991),
.B(n_12028),
.Y(n_13017)
);

HB1xp67_ASAP7_75t_L g13018 ( 
.A(n_12092),
.Y(n_13018)
);

OA21x2_ASAP7_75t_L g13019 ( 
.A1(n_12401),
.A2(n_11191),
.B(n_11156),
.Y(n_13019)
);

INVx1_ASAP7_75t_L g13020 ( 
.A(n_12576),
.Y(n_13020)
);

INVx1_ASAP7_75t_L g13021 ( 
.A(n_12576),
.Y(n_13021)
);

INVx1_ASAP7_75t_L g13022 ( 
.A(n_12589),
.Y(n_13022)
);

BUFx3_ASAP7_75t_L g13023 ( 
.A(n_12785),
.Y(n_13023)
);

BUFx3_ASAP7_75t_L g13024 ( 
.A(n_12785),
.Y(n_13024)
);

INVx2_ASAP7_75t_L g13025 ( 
.A(n_12841),
.Y(n_13025)
);

INVx2_ASAP7_75t_SL g13026 ( 
.A(n_11650),
.Y(n_13026)
);

INVx1_ASAP7_75t_L g13027 ( 
.A(n_12589),
.Y(n_13027)
);

OAI21x1_ASAP7_75t_L g13028 ( 
.A1(n_12306),
.A2(n_11164),
.B(n_10245),
.Y(n_13028)
);

NAND2xp5_ASAP7_75t_L g13029 ( 
.A(n_12234),
.B(n_9641),
.Y(n_13029)
);

INVx1_ASAP7_75t_L g13030 ( 
.A(n_12603),
.Y(n_13030)
);

AND2x2_ASAP7_75t_L g13031 ( 
.A(n_12028),
.B(n_11135),
.Y(n_13031)
);

INVx1_ASAP7_75t_L g13032 ( 
.A(n_12603),
.Y(n_13032)
);

INVx2_ASAP7_75t_L g13033 ( 
.A(n_12841),
.Y(n_13033)
);

INVx1_ASAP7_75t_L g13034 ( 
.A(n_12640),
.Y(n_13034)
);

INVx1_ASAP7_75t_L g13035 ( 
.A(n_12640),
.Y(n_13035)
);

INVxp67_ASAP7_75t_SL g13036 ( 
.A(n_12443),
.Y(n_13036)
);

NOR2xp33_ASAP7_75t_L g13037 ( 
.A(n_11906),
.B(n_10116),
.Y(n_13037)
);

CKINVDCx20_ASAP7_75t_R g13038 ( 
.A(n_11713),
.Y(n_13038)
);

INVx2_ASAP7_75t_L g13039 ( 
.A(n_11672),
.Y(n_13039)
);

INVx3_ASAP7_75t_L g13040 ( 
.A(n_12149),
.Y(n_13040)
);

AND2x4_ASAP7_75t_L g13041 ( 
.A(n_12420),
.B(n_11135),
.Y(n_13041)
);

AND2x2_ASAP7_75t_L g13042 ( 
.A(n_12073),
.B(n_11234),
.Y(n_13042)
);

INVx3_ASAP7_75t_L g13043 ( 
.A(n_12149),
.Y(n_13043)
);

INVx1_ASAP7_75t_L g13044 ( 
.A(n_12664),
.Y(n_13044)
);

INVx3_ASAP7_75t_L g13045 ( 
.A(n_11665),
.Y(n_13045)
);

INVx2_ASAP7_75t_L g13046 ( 
.A(n_11699),
.Y(n_13046)
);

INVx1_ASAP7_75t_L g13047 ( 
.A(n_12664),
.Y(n_13047)
);

INVx2_ASAP7_75t_L g13048 ( 
.A(n_11732),
.Y(n_13048)
);

NAND2xp5_ASAP7_75t_L g13049 ( 
.A(n_12411),
.B(n_9641),
.Y(n_13049)
);

OA21x2_ASAP7_75t_L g13050 ( 
.A1(n_12401),
.A2(n_11207),
.B(n_11192),
.Y(n_13050)
);

INVx1_ASAP7_75t_L g13051 ( 
.A(n_12097),
.Y(n_13051)
);

INVx1_ASAP7_75t_L g13052 ( 
.A(n_12097),
.Y(n_13052)
);

OR2x6_ASAP7_75t_L g13053 ( 
.A(n_12047),
.B(n_11234),
.Y(n_13053)
);

INVxp67_ASAP7_75t_L g13054 ( 
.A(n_12170),
.Y(n_13054)
);

INVx1_ASAP7_75t_L g13055 ( 
.A(n_12143),
.Y(n_13055)
);

NAND2xp5_ASAP7_75t_SL g13056 ( 
.A(n_11635),
.B(n_11234),
.Y(n_13056)
);

INVx2_ASAP7_75t_SL g13057 ( 
.A(n_11839),
.Y(n_13057)
);

INVx1_ASAP7_75t_L g13058 ( 
.A(n_12143),
.Y(n_13058)
);

OAI22xp33_ASAP7_75t_SL g13059 ( 
.A1(n_12333),
.A2(n_10319),
.B1(n_10499),
.B2(n_10268),
.Y(n_13059)
);

HB1xp67_ASAP7_75t_L g13060 ( 
.A(n_12170),
.Y(n_13060)
);

BUFx3_ASAP7_75t_L g13061 ( 
.A(n_11877),
.Y(n_13061)
);

INVxp33_ASAP7_75t_L g13062 ( 
.A(n_11799),
.Y(n_13062)
);

INVx2_ASAP7_75t_L g13063 ( 
.A(n_12214),
.Y(n_13063)
);

INVx1_ASAP7_75t_L g13064 ( 
.A(n_12204),
.Y(n_13064)
);

AO21x2_ASAP7_75t_L g13065 ( 
.A1(n_12326),
.A2(n_10999),
.B(n_10954),
.Y(n_13065)
);

INVx1_ASAP7_75t_L g13066 ( 
.A(n_12204),
.Y(n_13066)
);

INVx2_ASAP7_75t_SL g13067 ( 
.A(n_11839),
.Y(n_13067)
);

INVx3_ASAP7_75t_L g13068 ( 
.A(n_11665),
.Y(n_13068)
);

INVx2_ASAP7_75t_L g13069 ( 
.A(n_12228),
.Y(n_13069)
);

AND2x2_ASAP7_75t_L g13070 ( 
.A(n_12073),
.B(n_11234),
.Y(n_13070)
);

BUFx3_ASAP7_75t_L g13071 ( 
.A(n_11828),
.Y(n_13071)
);

INVx2_ASAP7_75t_L g13072 ( 
.A(n_11633),
.Y(n_13072)
);

INVx1_ASAP7_75t_L g13073 ( 
.A(n_12209),
.Y(n_13073)
);

BUFx3_ASAP7_75t_L g13074 ( 
.A(n_11828),
.Y(n_13074)
);

HB1xp67_ASAP7_75t_L g13075 ( 
.A(n_12209),
.Y(n_13075)
);

OA21x2_ASAP7_75t_L g13076 ( 
.A1(n_12851),
.A2(n_11207),
.B(n_11192),
.Y(n_13076)
);

INVxp33_ASAP7_75t_L g13077 ( 
.A(n_12259),
.Y(n_13077)
);

INVx2_ASAP7_75t_L g13078 ( 
.A(n_11639),
.Y(n_13078)
);

OA21x2_ASAP7_75t_L g13079 ( 
.A1(n_12851),
.A2(n_11207),
.B(n_11192),
.Y(n_13079)
);

AND2x2_ASAP7_75t_L g13080 ( 
.A(n_12084),
.B(n_11393),
.Y(n_13080)
);

INVx2_ASAP7_75t_L g13081 ( 
.A(n_11644),
.Y(n_13081)
);

AND2x2_ASAP7_75t_L g13082 ( 
.A(n_12084),
.B(n_11393),
.Y(n_13082)
);

HB1xp67_ASAP7_75t_L g13083 ( 
.A(n_12211),
.Y(n_13083)
);

INVx1_ASAP7_75t_L g13084 ( 
.A(n_12211),
.Y(n_13084)
);

INVx2_ASAP7_75t_L g13085 ( 
.A(n_11670),
.Y(n_13085)
);

INVx1_ASAP7_75t_L g13086 ( 
.A(n_12222),
.Y(n_13086)
);

INVx3_ASAP7_75t_L g13087 ( 
.A(n_11669),
.Y(n_13087)
);

INVx2_ASAP7_75t_L g13088 ( 
.A(n_12117),
.Y(n_13088)
);

AND2x4_ASAP7_75t_L g13089 ( 
.A(n_12418),
.B(n_11393),
.Y(n_13089)
);

INVxp67_ASAP7_75t_SL g13090 ( 
.A(n_12443),
.Y(n_13090)
);

HB1xp67_ASAP7_75t_L g13091 ( 
.A(n_12222),
.Y(n_13091)
);

INVx2_ASAP7_75t_L g13092 ( 
.A(n_12118),
.Y(n_13092)
);

NOR2x1_ASAP7_75t_L g13093 ( 
.A(n_12045),
.B(n_11393),
.Y(n_13093)
);

OAI21x1_ASAP7_75t_L g13094 ( 
.A1(n_12534),
.A2(n_11164),
.B(n_10245),
.Y(n_13094)
);

BUFx3_ASAP7_75t_L g13095 ( 
.A(n_11877),
.Y(n_13095)
);

BUFx2_ASAP7_75t_L g13096 ( 
.A(n_12481),
.Y(n_13096)
);

INVx3_ASAP7_75t_L g13097 ( 
.A(n_11669),
.Y(n_13097)
);

INVx1_ASAP7_75t_L g13098 ( 
.A(n_12227),
.Y(n_13098)
);

OAI21xp5_ASAP7_75t_L g13099 ( 
.A1(n_12333),
.A2(n_11600),
.B(n_11558),
.Y(n_13099)
);

BUFx3_ASAP7_75t_L g13100 ( 
.A(n_11730),
.Y(n_13100)
);

BUFx2_ASAP7_75t_SL g13101 ( 
.A(n_12103),
.Y(n_13101)
);

AND2x2_ASAP7_75t_L g13102 ( 
.A(n_12096),
.B(n_11576),
.Y(n_13102)
);

INVx1_ASAP7_75t_L g13103 ( 
.A(n_12227),
.Y(n_13103)
);

OR2x2_ASAP7_75t_L g13104 ( 
.A(n_12030),
.B(n_9518),
.Y(n_13104)
);

NOR2xp33_ASAP7_75t_L g13105 ( 
.A(n_11906),
.B(n_9782),
.Y(n_13105)
);

INVx1_ASAP7_75t_L g13106 ( 
.A(n_12236),
.Y(n_13106)
);

INVx1_ASAP7_75t_L g13107 ( 
.A(n_12236),
.Y(n_13107)
);

INVx2_ASAP7_75t_L g13108 ( 
.A(n_12130),
.Y(n_13108)
);

HB1xp67_ASAP7_75t_L g13109 ( 
.A(n_12240),
.Y(n_13109)
);

INVx2_ASAP7_75t_L g13110 ( 
.A(n_12141),
.Y(n_13110)
);

INVx1_ASAP7_75t_L g13111 ( 
.A(n_12240),
.Y(n_13111)
);

BUFx3_ASAP7_75t_L g13112 ( 
.A(n_11730),
.Y(n_13112)
);

INVx2_ASAP7_75t_L g13113 ( 
.A(n_12827),
.Y(n_13113)
);

INVx1_ASAP7_75t_L g13114 ( 
.A(n_12250),
.Y(n_13114)
);

BUFx2_ASAP7_75t_L g13115 ( 
.A(n_12481),
.Y(n_13115)
);

HB1xp67_ASAP7_75t_L g13116 ( 
.A(n_12250),
.Y(n_13116)
);

BUFx3_ASAP7_75t_L g13117 ( 
.A(n_12103),
.Y(n_13117)
);

INVx1_ASAP7_75t_SL g13118 ( 
.A(n_11825),
.Y(n_13118)
);

INVx1_ASAP7_75t_L g13119 ( 
.A(n_12255),
.Y(n_13119)
);

AOI21xp33_ASAP7_75t_L g13120 ( 
.A1(n_12206),
.A2(n_10773),
.B(n_10614),
.Y(n_13120)
);

OA21x2_ASAP7_75t_L g13121 ( 
.A1(n_12068),
.A2(n_11207),
.B(n_11192),
.Y(n_13121)
);

AND2x2_ASAP7_75t_L g13122 ( 
.A(n_12096),
.B(n_11576),
.Y(n_13122)
);

AO21x2_ASAP7_75t_L g13123 ( 
.A1(n_11893),
.A2(n_11006),
.B(n_10954),
.Y(n_13123)
);

AND2x2_ASAP7_75t_L g13124 ( 
.A(n_12107),
.B(n_11576),
.Y(n_13124)
);

INVx1_ASAP7_75t_L g13125 ( 
.A(n_12255),
.Y(n_13125)
);

INVx1_ASAP7_75t_L g13126 ( 
.A(n_12272),
.Y(n_13126)
);

BUFx4f_ASAP7_75t_SL g13127 ( 
.A(n_11959),
.Y(n_13127)
);

AND2x2_ASAP7_75t_L g13128 ( 
.A(n_12107),
.B(n_11399),
.Y(n_13128)
);

NAND2xp5_ASAP7_75t_L g13129 ( 
.A(n_12063),
.B(n_9641),
.Y(n_13129)
);

NAND2x1p5_ASAP7_75t_L g13130 ( 
.A(n_11641),
.B(n_11621),
.Y(n_13130)
);

INVx1_ASAP7_75t_L g13131 ( 
.A(n_12272),
.Y(n_13131)
);

AND2x2_ASAP7_75t_L g13132 ( 
.A(n_12167),
.B(n_11399),
.Y(n_13132)
);

HB1xp67_ASAP7_75t_L g13133 ( 
.A(n_12275),
.Y(n_13133)
);

INVxp67_ASAP7_75t_SL g13134 ( 
.A(n_12465),
.Y(n_13134)
);

INVx1_ASAP7_75t_L g13135 ( 
.A(n_12275),
.Y(n_13135)
);

AND2x2_ASAP7_75t_L g13136 ( 
.A(n_12167),
.B(n_11399),
.Y(n_13136)
);

OR2x6_ASAP7_75t_L g13137 ( 
.A(n_11929),
.B(n_9798),
.Y(n_13137)
);

INVx2_ASAP7_75t_L g13138 ( 
.A(n_12827),
.Y(n_13138)
);

INVx1_ASAP7_75t_L g13139 ( 
.A(n_12313),
.Y(n_13139)
);

OAI21x1_ASAP7_75t_L g13140 ( 
.A1(n_12534),
.A2(n_10245),
.B(n_10933),
.Y(n_13140)
);

OR2x2_ASAP7_75t_L g13141 ( 
.A(n_12483),
.B(n_9518),
.Y(n_13141)
);

INVx2_ASAP7_75t_L g13142 ( 
.A(n_12827),
.Y(n_13142)
);

INVx1_ASAP7_75t_L g13143 ( 
.A(n_12313),
.Y(n_13143)
);

INVx1_ASAP7_75t_L g13144 ( 
.A(n_12370),
.Y(n_13144)
);

INVx1_ASAP7_75t_L g13145 ( 
.A(n_12370),
.Y(n_13145)
);

BUFx6f_ASAP7_75t_L g13146 ( 
.A(n_12347),
.Y(n_13146)
);

INVx2_ASAP7_75t_L g13147 ( 
.A(n_12827),
.Y(n_13147)
);

INVx1_ASAP7_75t_L g13148 ( 
.A(n_12408),
.Y(n_13148)
);

INVx1_ASAP7_75t_L g13149 ( 
.A(n_12408),
.Y(n_13149)
);

INVx1_ASAP7_75t_L g13150 ( 
.A(n_11629),
.Y(n_13150)
);

INVx2_ASAP7_75t_L g13151 ( 
.A(n_12741),
.Y(n_13151)
);

INVx2_ASAP7_75t_SL g13152 ( 
.A(n_12347),
.Y(n_13152)
);

HB1xp67_ASAP7_75t_L g13153 ( 
.A(n_12821),
.Y(n_13153)
);

HB1xp67_ASAP7_75t_L g13154 ( 
.A(n_12821),
.Y(n_13154)
);

INVx2_ASAP7_75t_L g13155 ( 
.A(n_12749),
.Y(n_13155)
);

OAI21x1_ASAP7_75t_L g13156 ( 
.A1(n_12572),
.A2(n_10933),
.B(n_11187),
.Y(n_13156)
);

INVx2_ASAP7_75t_SL g13157 ( 
.A(n_12347),
.Y(n_13157)
);

INVx2_ASAP7_75t_L g13158 ( 
.A(n_12751),
.Y(n_13158)
);

INVx2_ASAP7_75t_L g13159 ( 
.A(n_12774),
.Y(n_13159)
);

OR2x2_ASAP7_75t_L g13160 ( 
.A(n_12501),
.B(n_9518),
.Y(n_13160)
);

INVx1_ASAP7_75t_L g13161 ( 
.A(n_11643),
.Y(n_13161)
);

OR2x2_ASAP7_75t_L g13162 ( 
.A(n_12764),
.B(n_9518),
.Y(n_13162)
);

INVx2_ASAP7_75t_L g13163 ( 
.A(n_12790),
.Y(n_13163)
);

AND2x2_ASAP7_75t_L g13164 ( 
.A(n_12188),
.B(n_11399),
.Y(n_13164)
);

AOI21xp5_ASAP7_75t_L g13165 ( 
.A1(n_12391),
.A2(n_11611),
.B(n_11602),
.Y(n_13165)
);

INVx1_ASAP7_75t_L g13166 ( 
.A(n_11652),
.Y(n_13166)
);

INVx1_ASAP7_75t_L g13167 ( 
.A(n_11653),
.Y(n_13167)
);

INVx2_ASAP7_75t_L g13168 ( 
.A(n_12793),
.Y(n_13168)
);

OAI21x1_ASAP7_75t_L g13169 ( 
.A1(n_12572),
.A2(n_10933),
.B(n_11187),
.Y(n_13169)
);

INVx2_ASAP7_75t_L g13170 ( 
.A(n_12800),
.Y(n_13170)
);

INVx1_ASAP7_75t_L g13171 ( 
.A(n_11664),
.Y(n_13171)
);

AO21x2_ASAP7_75t_L g13172 ( 
.A1(n_11893),
.A2(n_11006),
.B(n_10954),
.Y(n_13172)
);

INVx1_ASAP7_75t_L g13173 ( 
.A(n_11673),
.Y(n_13173)
);

INVx2_ASAP7_75t_L g13174 ( 
.A(n_12806),
.Y(n_13174)
);

AND2x2_ASAP7_75t_L g13175 ( 
.A(n_12188),
.B(n_12229),
.Y(n_13175)
);

INVx1_ASAP7_75t_L g13176 ( 
.A(n_11702),
.Y(n_13176)
);

NOR2x1_ASAP7_75t_SL g13177 ( 
.A(n_11742),
.B(n_10626),
.Y(n_13177)
);

INVx2_ASAP7_75t_L g13178 ( 
.A(n_12824),
.Y(n_13178)
);

INVx2_ASAP7_75t_L g13179 ( 
.A(n_12831),
.Y(n_13179)
);

INVx1_ASAP7_75t_L g13180 ( 
.A(n_11705),
.Y(n_13180)
);

INVx2_ASAP7_75t_L g13181 ( 
.A(n_12844),
.Y(n_13181)
);

INVx2_ASAP7_75t_L g13182 ( 
.A(n_12852),
.Y(n_13182)
);

AND2x2_ASAP7_75t_L g13183 ( 
.A(n_12229),
.B(n_11399),
.Y(n_13183)
);

AND2x4_ASAP7_75t_L g13184 ( 
.A(n_12042),
.B(n_11541),
.Y(n_13184)
);

HB1xp67_ASAP7_75t_L g13185 ( 
.A(n_12465),
.Y(n_13185)
);

HB1xp67_ASAP7_75t_L g13186 ( 
.A(n_12497),
.Y(n_13186)
);

HB1xp67_ASAP7_75t_L g13187 ( 
.A(n_12497),
.Y(n_13187)
);

INVx4_ASAP7_75t_L g13188 ( 
.A(n_11959),
.Y(n_13188)
);

BUFx3_ASAP7_75t_L g13189 ( 
.A(n_12606),
.Y(n_13189)
);

OA21x2_ASAP7_75t_L g13190 ( 
.A1(n_12068),
.A2(n_11220),
.B(n_11216),
.Y(n_13190)
);

AND2x2_ASAP7_75t_L g13191 ( 
.A(n_12444),
.B(n_11399),
.Y(n_13191)
);

INVx1_ASAP7_75t_L g13192 ( 
.A(n_11736),
.Y(n_13192)
);

AND2x2_ASAP7_75t_L g13193 ( 
.A(n_12444),
.B(n_11410),
.Y(n_13193)
);

INVx1_ASAP7_75t_L g13194 ( 
.A(n_11740),
.Y(n_13194)
);

HB1xp67_ASAP7_75t_L g13195 ( 
.A(n_12557),
.Y(n_13195)
);

INVx1_ASAP7_75t_L g13196 ( 
.A(n_11747),
.Y(n_13196)
);

INVx2_ASAP7_75t_L g13197 ( 
.A(n_12854),
.Y(n_13197)
);

OR2x2_ASAP7_75t_L g13198 ( 
.A(n_12768),
.B(n_9518),
.Y(n_13198)
);

INVx1_ASAP7_75t_L g13199 ( 
.A(n_11760),
.Y(n_13199)
);

AND2x2_ASAP7_75t_L g13200 ( 
.A(n_12474),
.B(n_11410),
.Y(n_13200)
);

AOI22xp33_ASAP7_75t_L g13201 ( 
.A1(n_11745),
.A2(n_11005),
.B1(n_10388),
.B2(n_10383),
.Y(n_13201)
);

INVx1_ASAP7_75t_L g13202 ( 
.A(n_11764),
.Y(n_13202)
);

INVx1_ASAP7_75t_L g13203 ( 
.A(n_11773),
.Y(n_13203)
);

AND2x4_ASAP7_75t_L g13204 ( 
.A(n_12042),
.B(n_11541),
.Y(n_13204)
);

INVx1_ASAP7_75t_L g13205 ( 
.A(n_11774),
.Y(n_13205)
);

OA21x2_ASAP7_75t_L g13206 ( 
.A1(n_12345),
.A2(n_11220),
.B(n_11216),
.Y(n_13206)
);

INVx1_ASAP7_75t_L g13207 ( 
.A(n_11777),
.Y(n_13207)
);

INVx1_ASAP7_75t_L g13208 ( 
.A(n_11779),
.Y(n_13208)
);

INVx1_ASAP7_75t_L g13209 ( 
.A(n_11789),
.Y(n_13209)
);

INVxp67_ASAP7_75t_SL g13210 ( 
.A(n_12557),
.Y(n_13210)
);

CKINVDCx5p33_ASAP7_75t_R g13211 ( 
.A(n_11978),
.Y(n_13211)
);

OA21x2_ASAP7_75t_L g13212 ( 
.A1(n_12345),
.A2(n_11220),
.B(n_11216),
.Y(n_13212)
);

INVx1_ASAP7_75t_L g13213 ( 
.A(n_11808),
.Y(n_13213)
);

INVx1_ASAP7_75t_L g13214 ( 
.A(n_11811),
.Y(n_13214)
);

AND2x2_ASAP7_75t_L g13215 ( 
.A(n_12474),
.B(n_11410),
.Y(n_13215)
);

INVx1_ASAP7_75t_L g13216 ( 
.A(n_11836),
.Y(n_13216)
);

INVx1_ASAP7_75t_L g13217 ( 
.A(n_11848),
.Y(n_13217)
);

BUFx2_ASAP7_75t_L g13218 ( 
.A(n_12876),
.Y(n_13218)
);

INVx2_ASAP7_75t_L g13219 ( 
.A(n_12856),
.Y(n_13219)
);

INVx1_ASAP7_75t_L g13220 ( 
.A(n_11852),
.Y(n_13220)
);

BUFx6f_ASAP7_75t_L g13221 ( 
.A(n_12347),
.Y(n_13221)
);

CKINVDCx6p67_ASAP7_75t_R g13222 ( 
.A(n_11986),
.Y(n_13222)
);

AND2x2_ASAP7_75t_L g13223 ( 
.A(n_12492),
.B(n_11410),
.Y(n_13223)
);

INVx2_ASAP7_75t_SL g13224 ( 
.A(n_12405),
.Y(n_13224)
);

OR2x2_ASAP7_75t_L g13225 ( 
.A(n_11787),
.B(n_9518),
.Y(n_13225)
);

INVx2_ASAP7_75t_L g13226 ( 
.A(n_12864),
.Y(n_13226)
);

INVx2_ASAP7_75t_L g13227 ( 
.A(n_12875),
.Y(n_13227)
);

AND2x4_ASAP7_75t_L g13228 ( 
.A(n_12055),
.B(n_11443),
.Y(n_13228)
);

INVx1_ASAP7_75t_L g13229 ( 
.A(n_11854),
.Y(n_13229)
);

HB1xp67_ASAP7_75t_L g13230 ( 
.A(n_12561),
.Y(n_13230)
);

INVx1_ASAP7_75t_L g13231 ( 
.A(n_11861),
.Y(n_13231)
);

OA21x2_ASAP7_75t_L g13232 ( 
.A1(n_12266),
.A2(n_11220),
.B(n_11216),
.Y(n_13232)
);

INVx1_ASAP7_75t_L g13233 ( 
.A(n_11888),
.Y(n_13233)
);

OAI21x1_ASAP7_75t_L g13234 ( 
.A1(n_12813),
.A2(n_11187),
.B(n_10319),
.Y(n_13234)
);

NAND2xp5_ASAP7_75t_L g13235 ( 
.A(n_11645),
.B(n_9648),
.Y(n_13235)
);

HB1xp67_ASAP7_75t_L g13236 ( 
.A(n_12561),
.Y(n_13236)
);

OAI21xp5_ASAP7_75t_L g13237 ( 
.A1(n_12293),
.A2(n_11868),
.B(n_11735),
.Y(n_13237)
);

NAND2xp5_ASAP7_75t_L g13238 ( 
.A(n_11703),
.B(n_9648),
.Y(n_13238)
);

INVx1_ASAP7_75t_L g13239 ( 
.A(n_11900),
.Y(n_13239)
);

INVx1_ASAP7_75t_L g13240 ( 
.A(n_11916),
.Y(n_13240)
);

INVx1_ASAP7_75t_L g13241 ( 
.A(n_11940),
.Y(n_13241)
);

BUFx3_ASAP7_75t_L g13242 ( 
.A(n_12606),
.Y(n_13242)
);

INVx2_ASAP7_75t_L g13243 ( 
.A(n_12885),
.Y(n_13243)
);

OAI21x1_ASAP7_75t_L g13244 ( 
.A1(n_12813),
.A2(n_12753),
.B(n_12710),
.Y(n_13244)
);

INVx2_ASAP7_75t_L g13245 ( 
.A(n_12888),
.Y(n_13245)
);

INVx2_ASAP7_75t_SL g13246 ( 
.A(n_12405),
.Y(n_13246)
);

INVx1_ASAP7_75t_L g13247 ( 
.A(n_11942),
.Y(n_13247)
);

INVx1_ASAP7_75t_L g13248 ( 
.A(n_11945),
.Y(n_13248)
);

OR2x2_ASAP7_75t_L g13249 ( 
.A(n_11951),
.B(n_9518),
.Y(n_13249)
);

OAI21x1_ASAP7_75t_L g13250 ( 
.A1(n_12710),
.A2(n_12791),
.B(n_12753),
.Y(n_13250)
);

INVx2_ASAP7_75t_L g13251 ( 
.A(n_12895),
.Y(n_13251)
);

HB1xp67_ASAP7_75t_L g13252 ( 
.A(n_12022),
.Y(n_13252)
);

OAI21x1_ASAP7_75t_L g13253 ( 
.A1(n_12791),
.A2(n_10319),
.B(n_10268),
.Y(n_13253)
);

CKINVDCx6p67_ASAP7_75t_R g13254 ( 
.A(n_12644),
.Y(n_13254)
);

INVx2_ASAP7_75t_L g13255 ( 
.A(n_12901),
.Y(n_13255)
);

INVxp67_ASAP7_75t_L g13256 ( 
.A(n_12353),
.Y(n_13256)
);

INVx1_ASAP7_75t_L g13257 ( 
.A(n_11966),
.Y(n_13257)
);

INVx2_ASAP7_75t_SL g13258 ( 
.A(n_12405),
.Y(n_13258)
);

NAND2x1_ASAP7_75t_L g13259 ( 
.A(n_12604),
.B(n_9976),
.Y(n_13259)
);

AOI21x1_ASAP7_75t_L g13260 ( 
.A1(n_11868),
.A2(n_10637),
.B(n_10242),
.Y(n_13260)
);

INVx2_ASAP7_75t_L g13261 ( 
.A(n_12658),
.Y(n_13261)
);

INVx1_ASAP7_75t_L g13262 ( 
.A(n_11992),
.Y(n_13262)
);

INVx1_ASAP7_75t_L g13263 ( 
.A(n_11997),
.Y(n_13263)
);

INVx1_ASAP7_75t_L g13264 ( 
.A(n_12023),
.Y(n_13264)
);

AND2x2_ASAP7_75t_L g13265 ( 
.A(n_12492),
.B(n_11410),
.Y(n_13265)
);

INVx1_ASAP7_75t_L g13266 ( 
.A(n_12027),
.Y(n_13266)
);

OAI21x1_ASAP7_75t_L g13267 ( 
.A1(n_12456),
.A2(n_12164),
.B(n_12041),
.Y(n_13267)
);

INVx2_ASAP7_75t_L g13268 ( 
.A(n_12702),
.Y(n_13268)
);

OR2x2_ASAP7_75t_L g13269 ( 
.A(n_11957),
.B(n_11958),
.Y(n_13269)
);

INVx1_ASAP7_75t_L g13270 ( 
.A(n_12036),
.Y(n_13270)
);

AND2x2_ASAP7_75t_L g13271 ( 
.A(n_12498),
.B(n_11410),
.Y(n_13271)
);

INVx3_ASAP7_75t_L g13272 ( 
.A(n_11681),
.Y(n_13272)
);

AO21x2_ASAP7_75t_L g13273 ( 
.A1(n_12524),
.A2(n_11041),
.B(n_11006),
.Y(n_13273)
);

INVx1_ASAP7_75t_SL g13274 ( 
.A(n_12244),
.Y(n_13274)
);

INVx1_ASAP7_75t_L g13275 ( 
.A(n_12039),
.Y(n_13275)
);

AO21x2_ASAP7_75t_L g13276 ( 
.A1(n_12524),
.A2(n_11041),
.B(n_10242),
.Y(n_13276)
);

INVx1_ASAP7_75t_L g13277 ( 
.A(n_12046),
.Y(n_13277)
);

AO21x2_ASAP7_75t_L g13278 ( 
.A1(n_12346),
.A2(n_11041),
.B(n_10201),
.Y(n_13278)
);

INVx2_ASAP7_75t_L g13279 ( 
.A(n_12729),
.Y(n_13279)
);

INVx1_ASAP7_75t_L g13280 ( 
.A(n_12058),
.Y(n_13280)
);

INVx2_ASAP7_75t_L g13281 ( 
.A(n_12740),
.Y(n_13281)
);

OA21x2_ASAP7_75t_L g13282 ( 
.A1(n_12266),
.A2(n_11436),
.B(n_11432),
.Y(n_13282)
);

NOR2xp33_ASAP7_75t_L g13283 ( 
.A(n_12040),
.B(n_8154),
.Y(n_13283)
);

HB1xp67_ASAP7_75t_L g13284 ( 
.A(n_11990),
.Y(n_13284)
);

INVx1_ASAP7_75t_L g13285 ( 
.A(n_12069),
.Y(n_13285)
);

INVx1_ASAP7_75t_L g13286 ( 
.A(n_12080),
.Y(n_13286)
);

INVx1_ASAP7_75t_L g13287 ( 
.A(n_12081),
.Y(n_13287)
);

OR2x6_ASAP7_75t_L g13288 ( 
.A(n_11989),
.B(n_9847),
.Y(n_13288)
);

INVx1_ASAP7_75t_L g13289 ( 
.A(n_12105),
.Y(n_13289)
);

INVx1_ASAP7_75t_L g13290 ( 
.A(n_12116),
.Y(n_13290)
);

INVx1_ASAP7_75t_L g13291 ( 
.A(n_12129),
.Y(n_13291)
);

INVx1_ASAP7_75t_L g13292 ( 
.A(n_12138),
.Y(n_13292)
);

INVx11_ASAP7_75t_L g13293 ( 
.A(n_12876),
.Y(n_13293)
);

NAND2x1_ASAP7_75t_L g13294 ( 
.A(n_12624),
.B(n_9976),
.Y(n_13294)
);

INVx1_ASAP7_75t_L g13295 ( 
.A(n_12142),
.Y(n_13295)
);

AOI21xp33_ASAP7_75t_L g13296 ( 
.A1(n_11791),
.A2(n_10773),
.B(n_10614),
.Y(n_13296)
);

INVx2_ASAP7_75t_L g13297 ( 
.A(n_12835),
.Y(n_13297)
);

INVx2_ASAP7_75t_L g13298 ( 
.A(n_12870),
.Y(n_13298)
);

HB1xp67_ASAP7_75t_L g13299 ( 
.A(n_12022),
.Y(n_13299)
);

INVx1_ASAP7_75t_L g13300 ( 
.A(n_12146),
.Y(n_13300)
);

BUFx2_ASAP7_75t_L g13301 ( 
.A(n_12797),
.Y(n_13301)
);

INVx2_ASAP7_75t_L g13302 ( 
.A(n_12289),
.Y(n_13302)
);

AO21x1_ASAP7_75t_L g13303 ( 
.A1(n_12365),
.A2(n_12374),
.B(n_12397),
.Y(n_13303)
);

BUFx4f_ASAP7_75t_L g13304 ( 
.A(n_12405),
.Y(n_13304)
);

INVx1_ASAP7_75t_L g13305 ( 
.A(n_12150),
.Y(n_13305)
);

INVx1_ASAP7_75t_L g13306 ( 
.A(n_12151),
.Y(n_13306)
);

BUFx3_ASAP7_75t_L g13307 ( 
.A(n_12644),
.Y(n_13307)
);

AO21x2_ASAP7_75t_L g13308 ( 
.A1(n_12346),
.A2(n_12635),
.B(n_11648),
.Y(n_13308)
);

BUFx3_ASAP7_75t_L g13309 ( 
.A(n_12179),
.Y(n_13309)
);

HB1xp67_ASAP7_75t_L g13310 ( 
.A(n_11990),
.Y(n_13310)
);

INVx1_ASAP7_75t_L g13311 ( 
.A(n_12152),
.Y(n_13311)
);

INVx3_ASAP7_75t_L g13312 ( 
.A(n_11681),
.Y(n_13312)
);

INVx1_ASAP7_75t_L g13313 ( 
.A(n_12154),
.Y(n_13313)
);

INVx2_ASAP7_75t_L g13314 ( 
.A(n_12289),
.Y(n_13314)
);

INVx2_ASAP7_75t_L g13315 ( 
.A(n_12312),
.Y(n_13315)
);

INVx2_ASAP7_75t_L g13316 ( 
.A(n_12312),
.Y(n_13316)
);

INVx3_ASAP7_75t_L g13317 ( 
.A(n_11682),
.Y(n_13317)
);

INVx2_ASAP7_75t_L g13318 ( 
.A(n_12377),
.Y(n_13318)
);

INVx3_ASAP7_75t_L g13319 ( 
.A(n_11682),
.Y(n_13319)
);

INVx1_ASAP7_75t_L g13320 ( 
.A(n_12212),
.Y(n_13320)
);

AND2x2_ASAP7_75t_L g13321 ( 
.A(n_12498),
.B(n_10231),
.Y(n_13321)
);

INVx2_ASAP7_75t_L g13322 ( 
.A(n_12377),
.Y(n_13322)
);

INVx1_ASAP7_75t_L g13323 ( 
.A(n_12221),
.Y(n_13323)
);

INVx1_ASAP7_75t_L g13324 ( 
.A(n_12251),
.Y(n_13324)
);

HB1xp67_ASAP7_75t_L g13325 ( 
.A(n_12000),
.Y(n_13325)
);

OA21x2_ASAP7_75t_L g13326 ( 
.A1(n_12393),
.A2(n_11436),
.B(n_11432),
.Y(n_13326)
);

INVx2_ASAP7_75t_SL g13327 ( 
.A(n_12550),
.Y(n_13327)
);

AO21x2_ASAP7_75t_L g13328 ( 
.A1(n_12635),
.A2(n_10201),
.B(n_11219),
.Y(n_13328)
);

INVx1_ASAP7_75t_L g13329 ( 
.A(n_12262),
.Y(n_13329)
);

HB1xp67_ASAP7_75t_L g13330 ( 
.A(n_12000),
.Y(n_13330)
);

INVx1_ASAP7_75t_L g13331 ( 
.A(n_12267),
.Y(n_13331)
);

INVx2_ASAP7_75t_L g13332 ( 
.A(n_12412),
.Y(n_13332)
);

INVx1_ASAP7_75t_L g13333 ( 
.A(n_12270),
.Y(n_13333)
);

AND2x2_ASAP7_75t_L g13334 ( 
.A(n_12514),
.B(n_10231),
.Y(n_13334)
);

AO21x2_ASAP7_75t_L g13335 ( 
.A1(n_11648),
.A2(n_11396),
.B(n_11219),
.Y(n_13335)
);

OA21x2_ASAP7_75t_L g13336 ( 
.A1(n_12393),
.A2(n_11436),
.B(n_11432),
.Y(n_13336)
);

OR2x2_ASAP7_75t_L g13337 ( 
.A(n_12136),
.B(n_9518),
.Y(n_13337)
);

INVx1_ASAP7_75t_L g13338 ( 
.A(n_12271),
.Y(n_13338)
);

OAI21x1_ASAP7_75t_L g13339 ( 
.A1(n_12456),
.A2(n_10319),
.B(n_10268),
.Y(n_13339)
);

INVx2_ASAP7_75t_L g13340 ( 
.A(n_12412),
.Y(n_13340)
);

INVx2_ASAP7_75t_L g13341 ( 
.A(n_12449),
.Y(n_13341)
);

AND2x2_ASAP7_75t_L g13342 ( 
.A(n_12514),
.B(n_12765),
.Y(n_13342)
);

INVx2_ASAP7_75t_L g13343 ( 
.A(n_12449),
.Y(n_13343)
);

INVx1_ASAP7_75t_L g13344 ( 
.A(n_12300),
.Y(n_13344)
);

INVx1_ASAP7_75t_L g13345 ( 
.A(n_12307),
.Y(n_13345)
);

INVx2_ASAP7_75t_L g13346 ( 
.A(n_12642),
.Y(n_13346)
);

INVx2_ASAP7_75t_L g13347 ( 
.A(n_12642),
.Y(n_13347)
);

INVx2_ASAP7_75t_L g13348 ( 
.A(n_12648),
.Y(n_13348)
);

AOI22xp33_ASAP7_75t_L g13349 ( 
.A1(n_11964),
.A2(n_11005),
.B1(n_10388),
.B2(n_10383),
.Y(n_13349)
);

INVx3_ASAP7_75t_L g13350 ( 
.A(n_11647),
.Y(n_13350)
);

INVx1_ASAP7_75t_L g13351 ( 
.A(n_12320),
.Y(n_13351)
);

BUFx10_ASAP7_75t_L g13352 ( 
.A(n_12550),
.Y(n_13352)
);

INVx2_ASAP7_75t_L g13353 ( 
.A(n_12648),
.Y(n_13353)
);

INVx4_ASAP7_75t_L g13354 ( 
.A(n_12550),
.Y(n_13354)
);

BUFx2_ASAP7_75t_L g13355 ( 
.A(n_12797),
.Y(n_13355)
);

AND2x2_ASAP7_75t_L g13356 ( 
.A(n_12765),
.B(n_10231),
.Y(n_13356)
);

NAND2xp5_ASAP7_75t_L g13357 ( 
.A(n_11686),
.B(n_9648),
.Y(n_13357)
);

INVxp67_ASAP7_75t_L g13358 ( 
.A(n_12618),
.Y(n_13358)
);

INVx1_ASAP7_75t_L g13359 ( 
.A(n_12327),
.Y(n_13359)
);

OR2x2_ASAP7_75t_L g13360 ( 
.A(n_12340),
.B(n_10227),
.Y(n_13360)
);

BUFx3_ASAP7_75t_L g13361 ( 
.A(n_12550),
.Y(n_13361)
);

BUFx2_ASAP7_75t_SL g13362 ( 
.A(n_12179),
.Y(n_13362)
);

BUFx2_ASAP7_75t_L g13363 ( 
.A(n_12055),
.Y(n_13363)
);

AND2x2_ASAP7_75t_L g13364 ( 
.A(n_12770),
.B(n_10283),
.Y(n_13364)
);

NOR2xp33_ASAP7_75t_L g13365 ( 
.A(n_12040),
.B(n_12064),
.Y(n_13365)
);

INVx3_ASAP7_75t_L g13366 ( 
.A(n_11647),
.Y(n_13366)
);

AND2x2_ASAP7_75t_L g13367 ( 
.A(n_12770),
.B(n_10283),
.Y(n_13367)
);

OR2x2_ASAP7_75t_L g13368 ( 
.A(n_12342),
.B(n_10227),
.Y(n_13368)
);

INVx1_ASAP7_75t_L g13369 ( 
.A(n_12331),
.Y(n_13369)
);

OA21x2_ASAP7_75t_L g13370 ( 
.A1(n_12086),
.A2(n_11436),
.B(n_11432),
.Y(n_13370)
);

INVx2_ASAP7_75t_L g13371 ( 
.A(n_12671),
.Y(n_13371)
);

NAND2xp5_ASAP7_75t_L g13372 ( 
.A(n_12614),
.B(n_9648),
.Y(n_13372)
);

OR2x2_ASAP7_75t_L g13373 ( 
.A(n_12332),
.B(n_10227),
.Y(n_13373)
);

INVx1_ASAP7_75t_L g13374 ( 
.A(n_12335),
.Y(n_13374)
);

INVx1_ASAP7_75t_L g13375 ( 
.A(n_12358),
.Y(n_13375)
);

INVx2_ASAP7_75t_L g13376 ( 
.A(n_12671),
.Y(n_13376)
);

INVx3_ASAP7_75t_L g13377 ( 
.A(n_11647),
.Y(n_13377)
);

AND2x4_ASAP7_75t_SL g13378 ( 
.A(n_11981),
.B(n_8183),
.Y(n_13378)
);

INVx3_ASAP7_75t_L g13379 ( 
.A(n_11678),
.Y(n_13379)
);

AO21x2_ASAP7_75t_L g13380 ( 
.A1(n_12100),
.A2(n_11481),
.B(n_11396),
.Y(n_13380)
);

INVx2_ASAP7_75t_L g13381 ( 
.A(n_12826),
.Y(n_13381)
);

AOI22xp33_ASAP7_75t_L g13382 ( 
.A1(n_11939),
.A2(n_11005),
.B1(n_10388),
.B2(n_10383),
.Y(n_13382)
);

BUFx2_ASAP7_75t_L g13383 ( 
.A(n_12162),
.Y(n_13383)
);

AND2x4_ASAP7_75t_L g13384 ( 
.A(n_12162),
.B(n_10283),
.Y(n_13384)
);

AOI21xp33_ASAP7_75t_SL g13385 ( 
.A1(n_11978),
.A2(n_8685),
.B(n_8671),
.Y(n_13385)
);

INVx2_ASAP7_75t_L g13386 ( 
.A(n_12826),
.Y(n_13386)
);

INVx3_ASAP7_75t_L g13387 ( 
.A(n_11678),
.Y(n_13387)
);

INVx2_ASAP7_75t_L g13388 ( 
.A(n_11793),
.Y(n_13388)
);

INVx2_ASAP7_75t_L g13389 ( 
.A(n_11796),
.Y(n_13389)
);

AND2x4_ASAP7_75t_L g13390 ( 
.A(n_12213),
.B(n_10286),
.Y(n_13390)
);

INVx2_ASAP7_75t_L g13391 ( 
.A(n_11800),
.Y(n_13391)
);

BUFx2_ASAP7_75t_L g13392 ( 
.A(n_12213),
.Y(n_13392)
);

BUFx2_ASAP7_75t_L g13393 ( 
.A(n_12808),
.Y(n_13393)
);

INVx1_ASAP7_75t_L g13394 ( 
.A(n_12368),
.Y(n_13394)
);

INVx1_ASAP7_75t_L g13395 ( 
.A(n_12380),
.Y(n_13395)
);

INVxp67_ASAP7_75t_L g13396 ( 
.A(n_12830),
.Y(n_13396)
);

INVx2_ASAP7_75t_L g13397 ( 
.A(n_11995),
.Y(n_13397)
);

INVx2_ASAP7_75t_L g13398 ( 
.A(n_12144),
.Y(n_13398)
);

INVx1_ASAP7_75t_L g13399 ( 
.A(n_12388),
.Y(n_13399)
);

NAND2xp5_ASAP7_75t_L g13400 ( 
.A(n_12134),
.B(n_9648),
.Y(n_13400)
);

OAI22xp5_ASAP7_75t_L g13401 ( 
.A1(n_12453),
.A2(n_11418),
.B1(n_11419),
.B2(n_11397),
.Y(n_13401)
);

BUFx2_ASAP7_75t_L g13402 ( 
.A(n_12808),
.Y(n_13402)
);

INVx1_ASAP7_75t_L g13403 ( 
.A(n_12396),
.Y(n_13403)
);

INVxp67_ASAP7_75t_SL g13404 ( 
.A(n_12011),
.Y(n_13404)
);

BUFx2_ASAP7_75t_L g13405 ( 
.A(n_12808),
.Y(n_13405)
);

AO21x1_ASAP7_75t_SL g13406 ( 
.A1(n_11688),
.A2(n_10364),
.B(n_10355),
.Y(n_13406)
);

INVx2_ASAP7_75t_SL g13407 ( 
.A(n_12808),
.Y(n_13407)
);

OR2x2_ASAP7_75t_L g13408 ( 
.A(n_12140),
.B(n_10227),
.Y(n_13408)
);

AND2x2_ASAP7_75t_L g13409 ( 
.A(n_12846),
.B(n_10286),
.Y(n_13409)
);

BUFx2_ASAP7_75t_L g13410 ( 
.A(n_12006),
.Y(n_13410)
);

INVx1_ASAP7_75t_L g13411 ( 
.A(n_12409),
.Y(n_13411)
);

INVx1_ASAP7_75t_L g13412 ( 
.A(n_12414),
.Y(n_13412)
);

OR2x6_ASAP7_75t_L g13413 ( 
.A(n_11742),
.B(n_12515),
.Y(n_13413)
);

HB1xp67_ASAP7_75t_L g13414 ( 
.A(n_12011),
.Y(n_13414)
);

INVx2_ASAP7_75t_L g13415 ( 
.A(n_12148),
.Y(n_13415)
);

INVx2_ASAP7_75t_L g13416 ( 
.A(n_12153),
.Y(n_13416)
);

OA21x2_ASAP7_75t_L g13417 ( 
.A1(n_12086),
.A2(n_11253),
.B(n_11223),
.Y(n_13417)
);

OR2x2_ASAP7_75t_L g13418 ( 
.A(n_12174),
.B(n_10227),
.Y(n_13418)
);

INVx2_ASAP7_75t_L g13419 ( 
.A(n_12156),
.Y(n_13419)
);

AOI21x1_ASAP7_75t_L g13420 ( 
.A1(n_11802),
.A2(n_10295),
.B(n_10286),
.Y(n_13420)
);

INVx2_ASAP7_75t_L g13421 ( 
.A(n_12157),
.Y(n_13421)
);

OR2x2_ASAP7_75t_L g13422 ( 
.A(n_12185),
.B(n_10457),
.Y(n_13422)
);

INVx1_ASAP7_75t_L g13423 ( 
.A(n_12426),
.Y(n_13423)
);

INVx2_ASAP7_75t_L g13424 ( 
.A(n_12160),
.Y(n_13424)
);

INVx2_ASAP7_75t_L g13425 ( 
.A(n_12177),
.Y(n_13425)
);

INVx1_ASAP7_75t_L g13426 ( 
.A(n_12428),
.Y(n_13426)
);

CKINVDCx5p33_ASAP7_75t_R g13427 ( 
.A(n_12088),
.Y(n_13427)
);

INVx1_ASAP7_75t_L g13428 ( 
.A(n_12433),
.Y(n_13428)
);

INVx1_ASAP7_75t_L g13429 ( 
.A(n_12434),
.Y(n_13429)
);

AND2x2_ASAP7_75t_L g13430 ( 
.A(n_12846),
.B(n_12066),
.Y(n_13430)
);

INVx1_ASAP7_75t_L g13431 ( 
.A(n_12463),
.Y(n_13431)
);

INVx2_ASAP7_75t_L g13432 ( 
.A(n_12181),
.Y(n_13432)
);

OR2x2_ASAP7_75t_L g13433 ( 
.A(n_12459),
.B(n_10457),
.Y(n_13433)
);

INVx2_ASAP7_75t_L g13434 ( 
.A(n_12182),
.Y(n_13434)
);

BUFx2_ASAP7_75t_L g13435 ( 
.A(n_12006),
.Y(n_13435)
);

HB1xp67_ASAP7_75t_L g13436 ( 
.A(n_12012),
.Y(n_13436)
);

INVx1_ASAP7_75t_L g13437 ( 
.A(n_12466),
.Y(n_13437)
);

AOI21xp5_ASAP7_75t_L g13438 ( 
.A1(n_12391),
.A2(n_11611),
.B(n_11602),
.Y(n_13438)
);

INVx2_ASAP7_75t_L g13439 ( 
.A(n_12192),
.Y(n_13439)
);

INVx1_ASAP7_75t_L g13440 ( 
.A(n_12469),
.Y(n_13440)
);

NAND2xp5_ASAP7_75t_L g13441 ( 
.A(n_12422),
.B(n_9650),
.Y(n_13441)
);

OAI21xp5_ASAP7_75t_L g13442 ( 
.A1(n_12453),
.A2(n_11476),
.B(n_10499),
.Y(n_13442)
);

INVx2_ASAP7_75t_L g13443 ( 
.A(n_12195),
.Y(n_13443)
);

INVx1_ASAP7_75t_L g13444 ( 
.A(n_12473),
.Y(n_13444)
);

OA21x2_ASAP7_75t_L g13445 ( 
.A1(n_12419),
.A2(n_11253),
.B(n_11223),
.Y(n_13445)
);

INVx2_ASAP7_75t_L g13446 ( 
.A(n_12224),
.Y(n_13446)
);

AND2x2_ASAP7_75t_L g13447 ( 
.A(n_12615),
.B(n_10295),
.Y(n_13447)
);

AND2x2_ASAP7_75t_L g13448 ( 
.A(n_12663),
.B(n_10295),
.Y(n_13448)
);

OR2x2_ASAP7_75t_L g13449 ( 
.A(n_12462),
.B(n_10457),
.Y(n_13449)
);

OR2x2_ASAP7_75t_L g13450 ( 
.A(n_11899),
.B(n_10457),
.Y(n_13450)
);

AND2x2_ASAP7_75t_L g13451 ( 
.A(n_12832),
.B(n_10310),
.Y(n_13451)
);

HB1xp67_ASAP7_75t_L g13452 ( 
.A(n_12012),
.Y(n_13452)
);

INVx2_ASAP7_75t_L g13453 ( 
.A(n_12239),
.Y(n_13453)
);

INVx2_ASAP7_75t_L g13454 ( 
.A(n_12246),
.Y(n_13454)
);

INVx2_ASAP7_75t_L g13455 ( 
.A(n_11685),
.Y(n_13455)
);

INVx2_ASAP7_75t_L g13456 ( 
.A(n_11711),
.Y(n_13456)
);

OR2x2_ASAP7_75t_L g13457 ( 
.A(n_11905),
.B(n_10457),
.Y(n_13457)
);

BUFx3_ASAP7_75t_L g13458 ( 
.A(n_12088),
.Y(n_13458)
);

BUFx3_ASAP7_75t_L g13459 ( 
.A(n_12172),
.Y(n_13459)
);

AND2x4_ASAP7_75t_L g13460 ( 
.A(n_12563),
.B(n_10310),
.Y(n_13460)
);

INVx1_ASAP7_75t_L g13461 ( 
.A(n_12476),
.Y(n_13461)
);

BUFx2_ASAP7_75t_L g13462 ( 
.A(n_12064),
.Y(n_13462)
);

INVxp33_ASAP7_75t_L g13463 ( 
.A(n_12748),
.Y(n_13463)
);

OAI21x1_ASAP7_75t_L g13464 ( 
.A1(n_12041),
.A2(n_10499),
.B(n_10268),
.Y(n_13464)
);

INVx2_ASAP7_75t_L g13465 ( 
.A(n_11722),
.Y(n_13465)
);

INVx2_ASAP7_75t_SL g13466 ( 
.A(n_12172),
.Y(n_13466)
);

AND2x4_ASAP7_75t_L g13467 ( 
.A(n_12563),
.B(n_10310),
.Y(n_13467)
);

OA21x2_ASAP7_75t_L g13468 ( 
.A1(n_12419),
.A2(n_11253),
.B(n_11223),
.Y(n_13468)
);

INVx2_ASAP7_75t_L g13469 ( 
.A(n_11728),
.Y(n_13469)
);

BUFx3_ASAP7_75t_L g13470 ( 
.A(n_12297),
.Y(n_13470)
);

INVx2_ASAP7_75t_SL g13471 ( 
.A(n_12254),
.Y(n_13471)
);

HB1xp67_ASAP7_75t_L g13472 ( 
.A(n_12071),
.Y(n_13472)
);

INVx1_ASAP7_75t_L g13473 ( 
.A(n_12479),
.Y(n_13473)
);

INVx2_ASAP7_75t_SL g13474 ( 
.A(n_12254),
.Y(n_13474)
);

INVx1_ASAP7_75t_L g13475 ( 
.A(n_12482),
.Y(n_13475)
);

BUFx6f_ASAP7_75t_L g13476 ( 
.A(n_12013),
.Y(n_13476)
);

INVx1_ASAP7_75t_L g13477 ( 
.A(n_12484),
.Y(n_13477)
);

INVx1_ASAP7_75t_L g13478 ( 
.A(n_12489),
.Y(n_13478)
);

INVx2_ASAP7_75t_L g13479 ( 
.A(n_11729),
.Y(n_13479)
);

INVx2_ASAP7_75t_L g13480 ( 
.A(n_11752),
.Y(n_13480)
);

CKINVDCx6p67_ASAP7_75t_R g13481 ( 
.A(n_12744),
.Y(n_13481)
);

OAI21x1_ASAP7_75t_L g13482 ( 
.A1(n_12164),
.A2(n_10527),
.B(n_10499),
.Y(n_13482)
);

NAND2x1_ASAP7_75t_L g13483 ( 
.A(n_12633),
.B(n_10009),
.Y(n_13483)
);

AND2x2_ASAP7_75t_L g13484 ( 
.A(n_12822),
.B(n_10327),
.Y(n_13484)
);

AO21x2_ASAP7_75t_L g13485 ( 
.A1(n_12435),
.A2(n_11481),
.B(n_10466),
.Y(n_13485)
);

AO21x2_ASAP7_75t_L g13486 ( 
.A1(n_12690),
.A2(n_10466),
.B(n_10464),
.Y(n_13486)
);

INVx3_ASAP7_75t_L g13487 ( 
.A(n_11816),
.Y(n_13487)
);

AO21x2_ASAP7_75t_L g13488 ( 
.A1(n_12180),
.A2(n_10466),
.B(n_10464),
.Y(n_13488)
);

INVx2_ASAP7_75t_L g13489 ( 
.A(n_11754),
.Y(n_13489)
);

INVx2_ASAP7_75t_L g13490 ( 
.A(n_11758),
.Y(n_13490)
);

INVx1_ASAP7_75t_L g13491 ( 
.A(n_12490),
.Y(n_13491)
);

AND2x2_ASAP7_75t_L g13492 ( 
.A(n_12822),
.B(n_10327),
.Y(n_13492)
);

INVx1_ASAP7_75t_L g13493 ( 
.A(n_12512),
.Y(n_13493)
);

AND2x2_ASAP7_75t_L g13494 ( 
.A(n_12869),
.B(n_10327),
.Y(n_13494)
);

INVx3_ASAP7_75t_L g13495 ( 
.A(n_11816),
.Y(n_13495)
);

AND2x4_ASAP7_75t_L g13496 ( 
.A(n_12013),
.B(n_10431),
.Y(n_13496)
);

INVx1_ASAP7_75t_L g13497 ( 
.A(n_12523),
.Y(n_13497)
);

INVx1_ASAP7_75t_L g13498 ( 
.A(n_12529),
.Y(n_13498)
);

AND2x2_ASAP7_75t_L g13499 ( 
.A(n_12869),
.B(n_10431),
.Y(n_13499)
);

INVx1_ASAP7_75t_L g13500 ( 
.A(n_12535),
.Y(n_13500)
);

INVx1_ASAP7_75t_L g13501 ( 
.A(n_12544),
.Y(n_13501)
);

OA21x2_ASAP7_75t_L g13502 ( 
.A1(n_12071),
.A2(n_11411),
.B(n_11260),
.Y(n_13502)
);

NOR2xp33_ASAP7_75t_L g13503 ( 
.A(n_11859),
.B(n_8685),
.Y(n_13503)
);

INVx1_ASAP7_75t_L g13504 ( 
.A(n_12567),
.Y(n_13504)
);

INVx3_ASAP7_75t_L g13505 ( 
.A(n_11816),
.Y(n_13505)
);

OAI21x1_ASAP7_75t_L g13506 ( 
.A1(n_12609),
.A2(n_10545),
.B(n_10527),
.Y(n_13506)
);

INVx1_ASAP7_75t_L g13507 ( 
.A(n_12577),
.Y(n_13507)
);

AND2x2_ASAP7_75t_L g13508 ( 
.A(n_12877),
.B(n_10431),
.Y(n_13508)
);

INVx1_ASAP7_75t_L g13509 ( 
.A(n_12578),
.Y(n_13509)
);

NOR2xp33_ASAP7_75t_L g13510 ( 
.A(n_11859),
.B(n_8725),
.Y(n_13510)
);

AOI21x1_ASAP7_75t_L g13511 ( 
.A1(n_11952),
.A2(n_10574),
.B(n_10446),
.Y(n_13511)
);

INVx1_ASAP7_75t_L g13512 ( 
.A(n_12590),
.Y(n_13512)
);

INVx2_ASAP7_75t_L g13513 ( 
.A(n_11769),
.Y(n_13513)
);

AO21x2_ASAP7_75t_L g13514 ( 
.A1(n_12252),
.A2(n_10466),
.B(n_10464),
.Y(n_13514)
);

INVx2_ASAP7_75t_L g13515 ( 
.A(n_11776),
.Y(n_13515)
);

AND2x4_ASAP7_75t_L g13516 ( 
.A(n_12761),
.B(n_10446),
.Y(n_13516)
);

INVx1_ASAP7_75t_L g13517 ( 
.A(n_12595),
.Y(n_13517)
);

CKINVDCx10_ASAP7_75t_R g13518 ( 
.A(n_11742),
.Y(n_13518)
);

INVx3_ASAP7_75t_L g13519 ( 
.A(n_11816),
.Y(n_13519)
);

INVxp67_ASAP7_75t_L g13520 ( 
.A(n_12619),
.Y(n_13520)
);

INVx1_ASAP7_75t_L g13521 ( 
.A(n_12632),
.Y(n_13521)
);

INVx3_ASAP7_75t_L g13522 ( 
.A(n_11816),
.Y(n_13522)
);

OAI21x1_ASAP7_75t_L g13523 ( 
.A1(n_12609),
.A2(n_10545),
.B(n_10527),
.Y(n_13523)
);

AND2x2_ASAP7_75t_L g13524 ( 
.A(n_12877),
.B(n_10446),
.Y(n_13524)
);

OR2x2_ASAP7_75t_L g13525 ( 
.A(n_11908),
.B(n_10457),
.Y(n_13525)
);

BUFx2_ASAP7_75t_L g13526 ( 
.A(n_12891),
.Y(n_13526)
);

OR2x2_ASAP7_75t_L g13527 ( 
.A(n_11870),
.B(n_10457),
.Y(n_13527)
);

INVx2_ASAP7_75t_L g13528 ( 
.A(n_11782),
.Y(n_13528)
);

INVx3_ASAP7_75t_L g13529 ( 
.A(n_11662),
.Y(n_13529)
);

OAI21x1_ASAP7_75t_L g13530 ( 
.A1(n_12562),
.A2(n_10545),
.B(n_10527),
.Y(n_13530)
);

INVx1_ASAP7_75t_L g13531 ( 
.A(n_12669),
.Y(n_13531)
);

BUFx6f_ASAP7_75t_L g13532 ( 
.A(n_12582),
.Y(n_13532)
);

AND2x2_ASAP7_75t_L g13533 ( 
.A(n_12287),
.B(n_10574),
.Y(n_13533)
);

INVx2_ASAP7_75t_L g13534 ( 
.A(n_11783),
.Y(n_13534)
);

INVx2_ASAP7_75t_L g13535 ( 
.A(n_11784),
.Y(n_13535)
);

INVx1_ASAP7_75t_L g13536 ( 
.A(n_12673),
.Y(n_13536)
);

AOI22xp33_ASAP7_75t_L g13537 ( 
.A1(n_11931),
.A2(n_10388),
.B1(n_10383),
.B2(n_10749),
.Y(n_13537)
);

BUFx6f_ASAP7_75t_L g13538 ( 
.A(n_12582),
.Y(n_13538)
);

AO21x2_ASAP7_75t_L g13539 ( 
.A1(n_12104),
.A2(n_10466),
.B(n_10464),
.Y(n_13539)
);

OR2x2_ASAP7_75t_L g13540 ( 
.A(n_11873),
.B(n_10457),
.Y(n_13540)
);

OR2x6_ASAP7_75t_L g13541 ( 
.A(n_12596),
.B(n_9847),
.Y(n_13541)
);

AND2x4_ASAP7_75t_L g13542 ( 
.A(n_12761),
.B(n_10574),
.Y(n_13542)
);

OAI21x1_ASAP7_75t_L g13543 ( 
.A1(n_12562),
.A2(n_10550),
.B(n_10545),
.Y(n_13543)
);

AOI21xp33_ASAP7_75t_L g13544 ( 
.A1(n_11921),
.A2(n_12190),
.B(n_11830),
.Y(n_13544)
);

AND2x2_ASAP7_75t_L g13545 ( 
.A(n_12292),
.B(n_10779),
.Y(n_13545)
);

AND2x2_ASAP7_75t_L g13546 ( 
.A(n_12619),
.B(n_10779),
.Y(n_13546)
);

INVx2_ASAP7_75t_L g13547 ( 
.A(n_12357),
.Y(n_13547)
);

INVx1_ASAP7_75t_L g13548 ( 
.A(n_12677),
.Y(n_13548)
);

CKINVDCx11_ASAP7_75t_R g13549 ( 
.A(n_12297),
.Y(n_13549)
);

INVx1_ASAP7_75t_L g13550 ( 
.A(n_12708),
.Y(n_13550)
);

INVx3_ASAP7_75t_L g13551 ( 
.A(n_11662),
.Y(n_13551)
);

AOI22xp33_ASAP7_75t_L g13552 ( 
.A1(n_11756),
.A2(n_10749),
.B1(n_10614),
.B2(n_10746),
.Y(n_13552)
);

HB1xp67_ASAP7_75t_L g13553 ( 
.A(n_11801),
.Y(n_13553)
);

NAND2xp5_ASAP7_75t_L g13554 ( 
.A(n_12009),
.B(n_9650),
.Y(n_13554)
);

AO21x2_ASAP7_75t_L g13555 ( 
.A1(n_12163),
.A2(n_10472),
.B(n_10610),
.Y(n_13555)
);

INVx2_ASAP7_75t_SL g13556 ( 
.A(n_12290),
.Y(n_13556)
);

AND2x2_ASAP7_75t_L g13557 ( 
.A(n_12545),
.B(n_10779),
.Y(n_13557)
);

INVx2_ASAP7_75t_L g13558 ( 
.A(n_11956),
.Y(n_13558)
);

INVx1_ASAP7_75t_L g13559 ( 
.A(n_12724),
.Y(n_13559)
);

OR2x2_ASAP7_75t_L g13560 ( 
.A(n_11874),
.B(n_11621),
.Y(n_13560)
);

INVx1_ASAP7_75t_L g13561 ( 
.A(n_12731),
.Y(n_13561)
);

INVx1_ASAP7_75t_L g13562 ( 
.A(n_12733),
.Y(n_13562)
);

INVx1_ASAP7_75t_L g13563 ( 
.A(n_12756),
.Y(n_13563)
);

INVx2_ASAP7_75t_L g13564 ( 
.A(n_12005),
.Y(n_13564)
);

OR2x2_ASAP7_75t_L g13565 ( 
.A(n_12450),
.B(n_11418),
.Y(n_13565)
);

INVx1_ASAP7_75t_L g13566 ( 
.A(n_12767),
.Y(n_13566)
);

INVx2_ASAP7_75t_L g13567 ( 
.A(n_12007),
.Y(n_13567)
);

INVx2_ASAP7_75t_L g13568 ( 
.A(n_11846),
.Y(n_13568)
);

INVx2_ASAP7_75t_L g13569 ( 
.A(n_11849),
.Y(n_13569)
);

INVx1_ASAP7_75t_L g13570 ( 
.A(n_12783),
.Y(n_13570)
);

INVx2_ASAP7_75t_SL g13571 ( 
.A(n_12290),
.Y(n_13571)
);

NAND2xp5_ASAP7_75t_L g13572 ( 
.A(n_12010),
.B(n_9650),
.Y(n_13572)
);

CKINVDCx20_ASAP7_75t_R g13573 ( 
.A(n_12495),
.Y(n_13573)
);

INVx3_ASAP7_75t_L g13574 ( 
.A(n_11662),
.Y(n_13574)
);

AND2x2_ASAP7_75t_L g13575 ( 
.A(n_12545),
.B(n_10899),
.Y(n_13575)
);

BUFx2_ASAP7_75t_L g13576 ( 
.A(n_12891),
.Y(n_13576)
);

INVx1_ASAP7_75t_L g13577 ( 
.A(n_12812),
.Y(n_13577)
);

INVx1_ASAP7_75t_L g13578 ( 
.A(n_12825),
.Y(n_13578)
);

NAND2x1_ASAP7_75t_L g13579 ( 
.A(n_12674),
.B(n_10009),
.Y(n_13579)
);

AND2x2_ASAP7_75t_L g13580 ( 
.A(n_12698),
.B(n_10899),
.Y(n_13580)
);

AND2x4_ASAP7_75t_L g13581 ( 
.A(n_12454),
.B(n_10420),
.Y(n_13581)
);

AO21x1_ASAP7_75t_SL g13582 ( 
.A1(n_11814),
.A2(n_10452),
.B(n_10441),
.Y(n_13582)
);

INVx2_ASAP7_75t_L g13583 ( 
.A(n_11864),
.Y(n_13583)
);

INVxp67_ASAP7_75t_SL g13584 ( 
.A(n_11856),
.Y(n_13584)
);

INVx1_ASAP7_75t_L g13585 ( 
.A(n_12837),
.Y(n_13585)
);

OAI222xp33_ASAP7_75t_L g13586 ( 
.A1(n_11631),
.A2(n_10550),
.B1(n_11419),
.B2(n_10626),
.C1(n_10583),
.C2(n_11292),
.Y(n_13586)
);

INVx1_ASAP7_75t_L g13587 ( 
.A(n_12848),
.Y(n_13587)
);

BUFx3_ASAP7_75t_L g13588 ( 
.A(n_12495),
.Y(n_13588)
);

AOI21x1_ASAP7_75t_L g13589 ( 
.A1(n_12651),
.A2(n_10674),
.B(n_10673),
.Y(n_13589)
);

INVx1_ASAP7_75t_L g13590 ( 
.A(n_12855),
.Y(n_13590)
);

INVx1_ASAP7_75t_L g13591 ( 
.A(n_12868),
.Y(n_13591)
);

AND2x2_ASAP7_75t_L g13592 ( 
.A(n_12698),
.B(n_10899),
.Y(n_13592)
);

INVx1_ASAP7_75t_L g13593 ( 
.A(n_12899),
.Y(n_13593)
);

OA21x2_ASAP7_75t_L g13594 ( 
.A1(n_12898),
.A2(n_11411),
.B(n_11260),
.Y(n_13594)
);

INVx1_ASAP7_75t_L g13595 ( 
.A(n_12903),
.Y(n_13595)
);

INVxp67_ASAP7_75t_L g13596 ( 
.A(n_11891),
.Y(n_13596)
);

INVx1_ASAP7_75t_L g13597 ( 
.A(n_12906),
.Y(n_13597)
);

OAI21x1_ASAP7_75t_L g13598 ( 
.A1(n_12723),
.A2(n_10550),
.B(n_10009),
.Y(n_13598)
);

INVx1_ASAP7_75t_L g13599 ( 
.A(n_12849),
.Y(n_13599)
);

INVx1_ASAP7_75t_L g13600 ( 
.A(n_12849),
.Y(n_13600)
);

INVx1_ASAP7_75t_L g13601 ( 
.A(n_12879),
.Y(n_13601)
);

HB1xp67_ASAP7_75t_L g13602 ( 
.A(n_11801),
.Y(n_13602)
);

AND2x2_ASAP7_75t_L g13603 ( 
.A(n_12884),
.B(n_10899),
.Y(n_13603)
);

INVx1_ASAP7_75t_L g13604 ( 
.A(n_12879),
.Y(n_13604)
);

INVx1_ASAP7_75t_L g13605 ( 
.A(n_12886),
.Y(n_13605)
);

INVx1_ASAP7_75t_L g13606 ( 
.A(n_12886),
.Y(n_13606)
);

HB1xp67_ASAP7_75t_SL g13607 ( 
.A(n_11891),
.Y(n_13607)
);

INVx2_ASAP7_75t_SL g13608 ( 
.A(n_12511),
.Y(n_13608)
);

INVx2_ASAP7_75t_SL g13609 ( 
.A(n_12511),
.Y(n_13609)
);

INVx1_ASAP7_75t_L g13610 ( 
.A(n_12893),
.Y(n_13610)
);

BUFx3_ASAP7_75t_L g13611 ( 
.A(n_12634),
.Y(n_13611)
);

INVx1_ASAP7_75t_L g13612 ( 
.A(n_12893),
.Y(n_13612)
);

INVx1_ASAP7_75t_L g13613 ( 
.A(n_12907),
.Y(n_13613)
);

AO21x2_ASAP7_75t_L g13614 ( 
.A1(n_12166),
.A2(n_10472),
.B(n_10610),
.Y(n_13614)
);

INVx1_ASAP7_75t_L g13615 ( 
.A(n_12907),
.Y(n_13615)
);

OAI21x1_ASAP7_75t_SL g13616 ( 
.A1(n_12304),
.A2(n_10605),
.B(n_10420),
.Y(n_13616)
);

BUFx3_ASAP7_75t_L g13617 ( 
.A(n_12634),
.Y(n_13617)
);

INVx3_ASAP7_75t_L g13618 ( 
.A(n_11714),
.Y(n_13618)
);

INVx2_ASAP7_75t_L g13619 ( 
.A(n_11875),
.Y(n_13619)
);

INVx2_ASAP7_75t_L g13620 ( 
.A(n_11882),
.Y(n_13620)
);

AO21x2_ASAP7_75t_L g13621 ( 
.A1(n_12169),
.A2(n_10472),
.B(n_10610),
.Y(n_13621)
);

NAND2xp5_ASAP7_75t_L g13622 ( 
.A(n_12083),
.B(n_12385),
.Y(n_13622)
);

INVx1_ASAP7_75t_L g13623 ( 
.A(n_12586),
.Y(n_13623)
);

INVx2_ASAP7_75t_L g13624 ( 
.A(n_11884),
.Y(n_13624)
);

HB1xp67_ASAP7_75t_L g13625 ( 
.A(n_11834),
.Y(n_13625)
);

NAND2xp5_ASAP7_75t_L g13626 ( 
.A(n_12389),
.B(n_9650),
.Y(n_13626)
);

HB1xp67_ASAP7_75t_L g13627 ( 
.A(n_11834),
.Y(n_13627)
);

INVx1_ASAP7_75t_L g13628 ( 
.A(n_12586),
.Y(n_13628)
);

INVx1_ASAP7_75t_L g13629 ( 
.A(n_12588),
.Y(n_13629)
);

INVx3_ASAP7_75t_L g13630 ( 
.A(n_11714),
.Y(n_13630)
);

INVx2_ASAP7_75t_L g13631 ( 
.A(n_11886),
.Y(n_13631)
);

INVx2_ASAP7_75t_L g13632 ( 
.A(n_11894),
.Y(n_13632)
);

INVx1_ASAP7_75t_L g13633 ( 
.A(n_12588),
.Y(n_13633)
);

INVx2_ASAP7_75t_L g13634 ( 
.A(n_11896),
.Y(n_13634)
);

INVx1_ASAP7_75t_L g13635 ( 
.A(n_12594),
.Y(n_13635)
);

INVx1_ASAP7_75t_L g13636 ( 
.A(n_12594),
.Y(n_13636)
);

INVx1_ASAP7_75t_L g13637 ( 
.A(n_12736),
.Y(n_13637)
);

INVx2_ASAP7_75t_L g13638 ( 
.A(n_11903),
.Y(n_13638)
);

INVx1_ASAP7_75t_L g13639 ( 
.A(n_12395),
.Y(n_13639)
);

OA21x2_ASAP7_75t_L g13640 ( 
.A1(n_12898),
.A2(n_11411),
.B(n_11260),
.Y(n_13640)
);

INVx2_ASAP7_75t_L g13641 ( 
.A(n_11909),
.Y(n_13641)
);

OR2x6_ASAP7_75t_L g13642 ( 
.A(n_12034),
.B(n_9847),
.Y(n_13642)
);

INVx1_ASAP7_75t_L g13643 ( 
.A(n_12186),
.Y(n_13643)
);

INVxp67_ASAP7_75t_L g13644 ( 
.A(n_12085),
.Y(n_13644)
);

AO21x2_ASAP7_75t_L g13645 ( 
.A1(n_12277),
.A2(n_10472),
.B(n_10610),
.Y(n_13645)
);

AO21x2_ASAP7_75t_L g13646 ( 
.A1(n_12862),
.A2(n_10472),
.B(n_10610),
.Y(n_13646)
);

OAI21x1_ASAP7_75t_L g13647 ( 
.A1(n_11826),
.A2(n_10550),
.B(n_10009),
.Y(n_13647)
);

INVx1_ASAP7_75t_L g13648 ( 
.A(n_12210),
.Y(n_13648)
);

INVx2_ASAP7_75t_L g13649 ( 
.A(n_11915),
.Y(n_13649)
);

HB1xp67_ASAP7_75t_L g13650 ( 
.A(n_11856),
.Y(n_13650)
);

OR2x6_ASAP7_75t_L g13651 ( 
.A(n_11879),
.B(n_9847),
.Y(n_13651)
);

INVx3_ASAP7_75t_L g13652 ( 
.A(n_11737),
.Y(n_13652)
);

OA21x2_ASAP7_75t_L g13653 ( 
.A1(n_12900),
.A2(n_11446),
.B(n_11416),
.Y(n_13653)
);

INVx2_ASAP7_75t_L g13654 ( 
.A(n_11919),
.Y(n_13654)
);

AND2x2_ASAP7_75t_L g13655 ( 
.A(n_12884),
.B(n_10899),
.Y(n_13655)
);

INVx1_ASAP7_75t_L g13656 ( 
.A(n_12219),
.Y(n_13656)
);

INVx1_ASAP7_75t_L g13657 ( 
.A(n_12237),
.Y(n_13657)
);

INVx1_ASAP7_75t_L g13658 ( 
.A(n_11820),
.Y(n_13658)
);

AOI21x1_ASAP7_75t_L g13659 ( 
.A1(n_11700),
.A2(n_10674),
.B(n_10673),
.Y(n_13659)
);

AO21x2_ASAP7_75t_L g13660 ( 
.A1(n_12862),
.A2(n_10695),
.B(n_10682),
.Y(n_13660)
);

INVx1_ASAP7_75t_L g13661 ( 
.A(n_12019),
.Y(n_13661)
);

INVx1_ASAP7_75t_L g13662 ( 
.A(n_12021),
.Y(n_13662)
);

AND2x2_ASAP7_75t_L g13663 ( 
.A(n_11925),
.B(n_10908),
.Y(n_13663)
);

INVx2_ASAP7_75t_SL g13664 ( 
.A(n_12584),
.Y(n_13664)
);

OR2x2_ASAP7_75t_L g13665 ( 
.A(n_12031),
.B(n_10750),
.Y(n_13665)
);

INVx1_ASAP7_75t_L g13666 ( 
.A(n_12048),
.Y(n_13666)
);

AND2x2_ASAP7_75t_L g13667 ( 
.A(n_11925),
.B(n_10908),
.Y(n_13667)
);

INVx1_ASAP7_75t_L g13668 ( 
.A(n_12051),
.Y(n_13668)
);

INVx1_ASAP7_75t_L g13669 ( 
.A(n_12059),
.Y(n_13669)
);

INVx1_ASAP7_75t_L g13670 ( 
.A(n_12072),
.Y(n_13670)
);

NOR2xp33_ASAP7_75t_L g13671 ( 
.A(n_12029),
.B(n_8725),
.Y(n_13671)
);

HB1xp67_ASAP7_75t_L g13672 ( 
.A(n_11872),
.Y(n_13672)
);

NAND2xp5_ASAP7_75t_L g13673 ( 
.A(n_12247),
.B(n_9650),
.Y(n_13673)
);

AND2x2_ASAP7_75t_L g13674 ( 
.A(n_11925),
.B(n_10908),
.Y(n_13674)
);

INVx2_ASAP7_75t_L g13675 ( 
.A(n_11928),
.Y(n_13675)
);

INVx3_ASAP7_75t_L g13676 ( 
.A(n_11737),
.Y(n_13676)
);

OR2x6_ASAP7_75t_L g13677 ( 
.A(n_11955),
.B(n_9847),
.Y(n_13677)
);

INVx1_ASAP7_75t_L g13678 ( 
.A(n_12090),
.Y(n_13678)
);

INVx2_ASAP7_75t_L g13679 ( 
.A(n_11941),
.Y(n_13679)
);

INVx1_ASAP7_75t_L g13680 ( 
.A(n_12094),
.Y(n_13680)
);

INVx2_ASAP7_75t_L g13681 ( 
.A(n_11953),
.Y(n_13681)
);

AO21x2_ASAP7_75t_L g13682 ( 
.A1(n_12223),
.A2(n_10695),
.B(n_10682),
.Y(n_13682)
);

INVxp67_ASAP7_75t_L g13683 ( 
.A(n_12165),
.Y(n_13683)
);

INVx1_ASAP7_75t_L g13684 ( 
.A(n_12123),
.Y(n_13684)
);

OR2x6_ASAP7_75t_L g13685 ( 
.A(n_11955),
.B(n_9847),
.Y(n_13685)
);

INVx2_ASAP7_75t_L g13686 ( 
.A(n_11962),
.Y(n_13686)
);

INVx1_ASAP7_75t_L g13687 ( 
.A(n_12135),
.Y(n_13687)
);

INVxp67_ASAP7_75t_L g13688 ( 
.A(n_11666),
.Y(n_13688)
);

INVx2_ASAP7_75t_L g13689 ( 
.A(n_11972),
.Y(n_13689)
);

HB1xp67_ASAP7_75t_L g13690 ( 
.A(n_11872),
.Y(n_13690)
);

OAI21xp5_ASAP7_75t_L g13691 ( 
.A1(n_12201),
.A2(n_11476),
.B(n_11424),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_12349),
.Y(n_13692)
);

INVx1_ASAP7_75t_L g13693 ( 
.A(n_12360),
.Y(n_13693)
);

INVx1_ASAP7_75t_L g13694 ( 
.A(n_12366),
.Y(n_13694)
);

AND2x4_ASAP7_75t_L g13695 ( 
.A(n_12454),
.B(n_10605),
.Y(n_13695)
);

AND2x2_ASAP7_75t_L g13696 ( 
.A(n_12268),
.B(n_12279),
.Y(n_13696)
);

AND2x2_ASAP7_75t_L g13697 ( 
.A(n_12268),
.B(n_10908),
.Y(n_13697)
);

AO21x2_ASAP7_75t_L g13698 ( 
.A1(n_11706),
.A2(n_10706),
.B(n_10701),
.Y(n_13698)
);

INVx1_ASAP7_75t_L g13699 ( 
.A(n_12549),
.Y(n_13699)
);

INVx1_ASAP7_75t_L g13700 ( 
.A(n_12559),
.Y(n_13700)
);

INVx3_ASAP7_75t_L g13701 ( 
.A(n_11781),
.Y(n_13701)
);

INVx1_ASAP7_75t_L g13702 ( 
.A(n_12249),
.Y(n_13702)
);

AND2x4_ASAP7_75t_L g13703 ( 
.A(n_12454),
.B(n_10832),
.Y(n_13703)
);

INVx2_ASAP7_75t_L g13704 ( 
.A(n_11979),
.Y(n_13704)
);

INVx2_ASAP7_75t_L g13705 ( 
.A(n_11988),
.Y(n_13705)
);

INVx1_ASAP7_75t_L g13706 ( 
.A(n_12299),
.Y(n_13706)
);

INVx1_ASAP7_75t_L g13707 ( 
.A(n_12316),
.Y(n_13707)
);

INVx3_ASAP7_75t_L g13708 ( 
.A(n_11781),
.Y(n_13708)
);

INVx1_ASAP7_75t_L g13709 ( 
.A(n_11706),
.Y(n_13709)
);

INVx1_ASAP7_75t_L g13710 ( 
.A(n_12178),
.Y(n_13710)
);

HB1xp67_ASAP7_75t_L g13711 ( 
.A(n_11889),
.Y(n_13711)
);

AO21x2_ASAP7_75t_L g13712 ( 
.A1(n_12178),
.A2(n_10706),
.B(n_10701),
.Y(n_13712)
);

INVx2_ASAP7_75t_L g13713 ( 
.A(n_11993),
.Y(n_13713)
);

AO31x2_ASAP7_75t_L g13714 ( 
.A1(n_12758),
.A2(n_10832),
.A3(n_10735),
.B(n_10738),
.Y(n_13714)
);

INVx1_ASAP7_75t_L g13715 ( 
.A(n_12522),
.Y(n_13715)
);

INVx1_ASAP7_75t_L g13716 ( 
.A(n_12532),
.Y(n_13716)
);

INVx2_ASAP7_75t_L g13717 ( 
.A(n_12440),
.Y(n_13717)
);

INVx2_ASAP7_75t_SL g13718 ( 
.A(n_12584),
.Y(n_13718)
);

AO21x2_ASAP7_75t_L g13719 ( 
.A1(n_12242),
.A2(n_10735),
.B(n_10719),
.Y(n_13719)
);

OAI21x1_ASAP7_75t_L g13720 ( 
.A1(n_11826),
.A2(n_10826),
.B(n_10820),
.Y(n_13720)
);

INVxp67_ASAP7_75t_L g13721 ( 
.A(n_11666),
.Y(n_13721)
);

INVx3_ASAP7_75t_L g13722 ( 
.A(n_11851),
.Y(n_13722)
);

INVx2_ASAP7_75t_L g13723 ( 
.A(n_12447),
.Y(n_13723)
);

INVx3_ASAP7_75t_L g13724 ( 
.A(n_11851),
.Y(n_13724)
);

INVx1_ASAP7_75t_L g13725 ( 
.A(n_12525),
.Y(n_13725)
);

INVx2_ASAP7_75t_L g13726 ( 
.A(n_12448),
.Y(n_13726)
);

AO21x2_ASAP7_75t_L g13727 ( 
.A1(n_12245),
.A2(n_10738),
.B(n_10719),
.Y(n_13727)
);

INVx1_ASAP7_75t_L g13728 ( 
.A(n_12546),
.Y(n_13728)
);

BUFx2_ASAP7_75t_L g13729 ( 
.A(n_12445),
.Y(n_13729)
);

INVx2_ASAP7_75t_L g13730 ( 
.A(n_12460),
.Y(n_13730)
);

INVx1_ASAP7_75t_L g13731 ( 
.A(n_12542),
.Y(n_13731)
);

INVx2_ASAP7_75t_L g13732 ( 
.A(n_12477),
.Y(n_13732)
);

INVx1_ASAP7_75t_L g13733 ( 
.A(n_12573),
.Y(n_13733)
);

INVx1_ASAP7_75t_L g13734 ( 
.A(n_12601),
.Y(n_13734)
);

BUFx4f_ASAP7_75t_SL g13735 ( 
.A(n_12371),
.Y(n_13735)
);

INVx2_ASAP7_75t_L g13736 ( 
.A(n_12478),
.Y(n_13736)
);

OR2x2_ASAP7_75t_L g13737 ( 
.A(n_11938),
.B(n_10750),
.Y(n_13737)
);

HB1xp67_ASAP7_75t_L g13738 ( 
.A(n_11889),
.Y(n_13738)
);

INVx1_ASAP7_75t_L g13739 ( 
.A(n_12564),
.Y(n_13739)
);

BUFx2_ASAP7_75t_L g13740 ( 
.A(n_12445),
.Y(n_13740)
);

AO21x2_ASAP7_75t_L g13741 ( 
.A1(n_12230),
.A2(n_10747),
.B(n_10744),
.Y(n_13741)
);

AOI21x1_ASAP7_75t_L g13742 ( 
.A1(n_11719),
.A2(n_10747),
.B(n_10744),
.Y(n_13742)
);

AO21x2_ASAP7_75t_L g13743 ( 
.A1(n_12190),
.A2(n_11963),
.B(n_11890),
.Y(n_13743)
);

HB1xp67_ASAP7_75t_L g13744 ( 
.A(n_11890),
.Y(n_13744)
);

OAI21x1_ASAP7_75t_L g13745 ( 
.A1(n_12285),
.A2(n_10826),
.B(n_10820),
.Y(n_13745)
);

INVx1_ASAP7_75t_L g13746 ( 
.A(n_12568),
.Y(n_13746)
);

INVx1_ASAP7_75t_L g13747 ( 
.A(n_12621),
.Y(n_13747)
);

OR2x2_ASAP7_75t_L g13748 ( 
.A(n_11943),
.B(n_10750),
.Y(n_13748)
);

AND2x2_ASAP7_75t_L g13749 ( 
.A(n_12268),
.B(n_10908),
.Y(n_13749)
);

AO31x2_ASAP7_75t_L g13750 ( 
.A1(n_11744),
.A2(n_10786),
.A3(n_10789),
.B(n_10776),
.Y(n_13750)
);

INVx1_ASAP7_75t_L g13751 ( 
.A(n_11983),
.Y(n_13751)
);

INVx3_ASAP7_75t_L g13752 ( 
.A(n_11803),
.Y(n_13752)
);

HB1xp67_ASAP7_75t_L g13753 ( 
.A(n_11963),
.Y(n_13753)
);

BUFx10_ASAP7_75t_L g13754 ( 
.A(n_12503),
.Y(n_13754)
);

INVx2_ASAP7_75t_L g13755 ( 
.A(n_12485),
.Y(n_13755)
);

CKINVDCx20_ASAP7_75t_R g13756 ( 
.A(n_12605),
.Y(n_13756)
);

INVx1_ASAP7_75t_L g13757 ( 
.A(n_11983),
.Y(n_13757)
);

INVx1_ASAP7_75t_L g13758 ( 
.A(n_11996),
.Y(n_13758)
);

INVx2_ASAP7_75t_L g13759 ( 
.A(n_12488),
.Y(n_13759)
);

INVx1_ASAP7_75t_L g13760 ( 
.A(n_11996),
.Y(n_13760)
);

INVx3_ASAP7_75t_L g13761 ( 
.A(n_11803),
.Y(n_13761)
);

INVxp33_ASAP7_75t_L g13762 ( 
.A(n_12792),
.Y(n_13762)
);

HB1xp67_ASAP7_75t_L g13763 ( 
.A(n_11727),
.Y(n_13763)
);

OAI21x1_ASAP7_75t_L g13764 ( 
.A1(n_12285),
.A2(n_10826),
.B(n_10820),
.Y(n_13764)
);

INVx1_ASAP7_75t_L g13765 ( 
.A(n_12003),
.Y(n_13765)
);

BUFx3_ASAP7_75t_L g13766 ( 
.A(n_12605),
.Y(n_13766)
);

INVx1_ASAP7_75t_L g13767 ( 
.A(n_12003),
.Y(n_13767)
);

NAND2xp5_ASAP7_75t_L g13768 ( 
.A(n_11731),
.B(n_12026),
.Y(n_13768)
);

INVx2_ASAP7_75t_SL g13769 ( 
.A(n_12217),
.Y(n_13769)
);

OR2x6_ASAP7_75t_L g13770 ( 
.A(n_11955),
.B(n_9888),
.Y(n_13770)
);

INVx1_ASAP7_75t_L g13771 ( 
.A(n_12014),
.Y(n_13771)
);

INVx2_ASAP7_75t_L g13772 ( 
.A(n_12491),
.Y(n_13772)
);

INVx3_ASAP7_75t_L g13773 ( 
.A(n_11803),
.Y(n_13773)
);

AO21x2_ASAP7_75t_L g13774 ( 
.A1(n_12193),
.A2(n_10786),
.B(n_10776),
.Y(n_13774)
);

BUFx6f_ASAP7_75t_L g13775 ( 
.A(n_12454),
.Y(n_13775)
);

INVx2_ASAP7_75t_L g13776 ( 
.A(n_12493),
.Y(n_13776)
);

CKINVDCx6p67_ASAP7_75t_R g13777 ( 
.A(n_12099),
.Y(n_13777)
);

INVx2_ASAP7_75t_L g13778 ( 
.A(n_12499),
.Y(n_13778)
);

INVx1_ASAP7_75t_L g13779 ( 
.A(n_12014),
.Y(n_13779)
);

HB1xp67_ASAP7_75t_L g13780 ( 
.A(n_11727),
.Y(n_13780)
);

INVx1_ASAP7_75t_L g13781 ( 
.A(n_12024),
.Y(n_13781)
);

NAND2xp5_ASAP7_75t_L g13782 ( 
.A(n_11838),
.B(n_9671),
.Y(n_13782)
);

INVx1_ASAP7_75t_L g13783 ( 
.A(n_12024),
.Y(n_13783)
);

INVx4_ASAP7_75t_SL g13784 ( 
.A(n_12802),
.Y(n_13784)
);

AND2x2_ASAP7_75t_L g13785 ( 
.A(n_12279),
.B(n_10960),
.Y(n_13785)
);

INVx1_ASAP7_75t_L g13786 ( 
.A(n_12038),
.Y(n_13786)
);

INVx1_ASAP7_75t_L g13787 ( 
.A(n_12038),
.Y(n_13787)
);

INVx1_ASAP7_75t_L g13788 ( 
.A(n_12057),
.Y(n_13788)
);

OR2x2_ASAP7_75t_L g13789 ( 
.A(n_12553),
.B(n_10750),
.Y(n_13789)
);

INVx1_ASAP7_75t_L g13790 ( 
.A(n_12057),
.Y(n_13790)
);

INVx2_ASAP7_75t_L g13791 ( 
.A(n_12505),
.Y(n_13791)
);

INVx1_ASAP7_75t_L g13792 ( 
.A(n_12106),
.Y(n_13792)
);

AOI21x1_ASAP7_75t_L g13793 ( 
.A1(n_12667),
.A2(n_10818),
.B(n_10789),
.Y(n_13793)
);

INVx2_ASAP7_75t_L g13794 ( 
.A(n_12506),
.Y(n_13794)
);

INVx2_ASAP7_75t_L g13795 ( 
.A(n_12513),
.Y(n_13795)
);

HB1xp67_ASAP7_75t_L g13796 ( 
.A(n_12857),
.Y(n_13796)
);

OR2x2_ASAP7_75t_L g13797 ( 
.A(n_11920),
.B(n_10750),
.Y(n_13797)
);

HB1xp67_ASAP7_75t_L g13798 ( 
.A(n_12857),
.Y(n_13798)
);

NAND2xp5_ASAP7_75t_L g13799 ( 
.A(n_11718),
.B(n_11720),
.Y(n_13799)
);

HB1xp67_ASAP7_75t_L g13800 ( 
.A(n_12087),
.Y(n_13800)
);

AOI22xp33_ASAP7_75t_L g13801 ( 
.A1(n_11974),
.A2(n_10749),
.B1(n_10614),
.B2(n_10746),
.Y(n_13801)
);

OR2x2_ASAP7_75t_L g13802 ( 
.A(n_11922),
.B(n_10750),
.Y(n_13802)
);

INVx2_ASAP7_75t_L g13803 ( 
.A(n_12516),
.Y(n_13803)
);

INVx4_ASAP7_75t_L g13804 ( 
.A(n_12802),
.Y(n_13804)
);

OAI21x1_ASAP7_75t_SL g13805 ( 
.A1(n_11695),
.A2(n_10778),
.B(n_9083),
.Y(n_13805)
);

OAI21x1_ASAP7_75t_L g13806 ( 
.A1(n_12317),
.A2(n_12781),
.B(n_12685),
.Y(n_13806)
);

BUFx12f_ASAP7_75t_L g13807 ( 
.A(n_12722),
.Y(n_13807)
);

INVx2_ASAP7_75t_L g13808 ( 
.A(n_12526),
.Y(n_13808)
);

HB1xp67_ASAP7_75t_L g13809 ( 
.A(n_12087),
.Y(n_13809)
);

INVx2_ASAP7_75t_L g13810 ( 
.A(n_12533),
.Y(n_13810)
);

HB1xp67_ASAP7_75t_L g13811 ( 
.A(n_12087),
.Y(n_13811)
);

INVx2_ASAP7_75t_L g13812 ( 
.A(n_12536),
.Y(n_13812)
);

OR2x6_ASAP7_75t_L g13813 ( 
.A(n_11980),
.B(n_9888),
.Y(n_13813)
);

INVxp67_ASAP7_75t_SL g13814 ( 
.A(n_12900),
.Y(n_13814)
);

INVx1_ASAP7_75t_L g13815 ( 
.A(n_12106),
.Y(n_13815)
);

INVx1_ASAP7_75t_L g13816 ( 
.A(n_12119),
.Y(n_13816)
);

AO21x2_ASAP7_75t_L g13817 ( 
.A1(n_12197),
.A2(n_10819),
.B(n_10818),
.Y(n_13817)
);

INVx2_ASAP7_75t_L g13818 ( 
.A(n_12541),
.Y(n_13818)
);

OR2x2_ASAP7_75t_L g13819 ( 
.A(n_11835),
.B(n_10750),
.Y(n_13819)
);

INVx2_ASAP7_75t_L g13820 ( 
.A(n_12543),
.Y(n_13820)
);

INVx1_ASAP7_75t_L g13821 ( 
.A(n_12119),
.Y(n_13821)
);

INVx2_ASAP7_75t_L g13822 ( 
.A(n_12217),
.Y(n_13822)
);

BUFx10_ASAP7_75t_L g13823 ( 
.A(n_12503),
.Y(n_13823)
);

AO21x2_ASAP7_75t_L g13824 ( 
.A1(n_12430),
.A2(n_10836),
.B(n_10819),
.Y(n_13824)
);

INVx1_ASAP7_75t_L g13825 ( 
.A(n_12127),
.Y(n_13825)
);

INVx1_ASAP7_75t_L g13826 ( 
.A(n_12127),
.Y(n_13826)
);

INVx1_ASAP7_75t_L g13827 ( 
.A(n_12131),
.Y(n_13827)
);

INVx2_ASAP7_75t_L g13828 ( 
.A(n_12337),
.Y(n_13828)
);

INVx1_ASAP7_75t_L g13829 ( 
.A(n_12131),
.Y(n_13829)
);

BUFx3_ASAP7_75t_L g13830 ( 
.A(n_12722),
.Y(n_13830)
);

INVx1_ASAP7_75t_L g13831 ( 
.A(n_12173),
.Y(n_13831)
);

INVx4_ASAP7_75t_L g13832 ( 
.A(n_12061),
.Y(n_13832)
);

INVx1_ASAP7_75t_L g13833 ( 
.A(n_12173),
.Y(n_13833)
);

HB1xp67_ASAP7_75t_L g13834 ( 
.A(n_12321),
.Y(n_13834)
);

INVx2_ASAP7_75t_L g13835 ( 
.A(n_12337),
.Y(n_13835)
);

OR2x6_ASAP7_75t_L g13836 ( 
.A(n_11980),
.B(n_9888),
.Y(n_13836)
);

INVx1_ASAP7_75t_L g13837 ( 
.A(n_12194),
.Y(n_13837)
);

OR2x2_ASAP7_75t_L g13838 ( 
.A(n_12693),
.B(n_10750),
.Y(n_13838)
);

INVx1_ASAP7_75t_L g13839 ( 
.A(n_12194),
.Y(n_13839)
);

AND2x2_ASAP7_75t_L g13840 ( 
.A(n_12279),
.B(n_10960),
.Y(n_13840)
);

INVx3_ASAP7_75t_SL g13841 ( 
.A(n_12061),
.Y(n_13841)
);

OAI21x1_ASAP7_75t_L g13842 ( 
.A1(n_12317),
.A2(n_9406),
.B(n_9321),
.Y(n_13842)
);

AND2x2_ASAP7_75t_L g13843 ( 
.A(n_12301),
.B(n_12341),
.Y(n_13843)
);

INVx1_ASAP7_75t_L g13844 ( 
.A(n_12216),
.Y(n_13844)
);

AND2x4_ASAP7_75t_L g13845 ( 
.A(n_12655),
.B(n_10443),
.Y(n_13845)
);

INVx2_ASAP7_75t_L g13846 ( 
.A(n_12359),
.Y(n_13846)
);

INVx1_ASAP7_75t_L g13847 ( 
.A(n_12216),
.Y(n_13847)
);

NAND2xp5_ASAP7_75t_L g13848 ( 
.A(n_11712),
.B(n_9671),
.Y(n_13848)
);

OR2x2_ASAP7_75t_L g13849 ( 
.A(n_12697),
.B(n_9569),
.Y(n_13849)
);

BUFx6f_ASAP7_75t_L g13850 ( 
.A(n_12655),
.Y(n_13850)
);

INVx3_ASAP7_75t_L g13851 ( 
.A(n_11806),
.Y(n_13851)
);

INVx2_ASAP7_75t_L g13852 ( 
.A(n_12359),
.Y(n_13852)
);

INVx2_ASAP7_75t_L g13853 ( 
.A(n_12362),
.Y(n_13853)
);

INVx2_ASAP7_75t_L g13854 ( 
.A(n_12362),
.Y(n_13854)
);

AND2x2_ASAP7_75t_L g13855 ( 
.A(n_12301),
.B(n_10960),
.Y(n_13855)
);

INVx1_ASAP7_75t_L g13856 ( 
.A(n_12060),
.Y(n_13856)
);

INVx4_ASAP7_75t_L g13857 ( 
.A(n_12061),
.Y(n_13857)
);

INVx2_ASAP7_75t_L g13858 ( 
.A(n_12373),
.Y(n_13858)
);

BUFx2_ASAP7_75t_L g13859 ( 
.A(n_12400),
.Y(n_13859)
);

AO21x2_ASAP7_75t_L g13860 ( 
.A1(n_11751),
.A2(n_10837),
.B(n_10836),
.Y(n_13860)
);

INVx2_ASAP7_75t_L g13861 ( 
.A(n_12373),
.Y(n_13861)
);

OR2x2_ASAP7_75t_L g13862 ( 
.A(n_12701),
.B(n_9569),
.Y(n_13862)
);

INVx1_ASAP7_75t_L g13863 ( 
.A(n_12102),
.Y(n_13863)
);

INVx1_ASAP7_75t_L g13864 ( 
.A(n_12218),
.Y(n_13864)
);

INVx1_ASAP7_75t_L g13865 ( 
.A(n_12125),
.Y(n_13865)
);

NAND2xp5_ASAP7_75t_L g13866 ( 
.A(n_11717),
.B(n_9671),
.Y(n_13866)
);

OAI21x1_ASAP7_75t_L g13867 ( 
.A1(n_12700),
.A2(n_9406),
.B(n_9321),
.Y(n_13867)
);

INVx2_ASAP7_75t_L g13868 ( 
.A(n_12437),
.Y(n_13868)
);

INVxp67_ASAP7_75t_L g13869 ( 
.A(n_12548),
.Y(n_13869)
);

BUFx3_ASAP7_75t_L g13870 ( 
.A(n_12734),
.Y(n_13870)
);

INVx2_ASAP7_75t_L g13871 ( 
.A(n_12437),
.Y(n_13871)
);

AND2x2_ASAP7_75t_L g13872 ( 
.A(n_12301),
.B(n_10960),
.Y(n_13872)
);

OAI21x1_ASAP7_75t_L g13873 ( 
.A1(n_12705),
.A2(n_9406),
.B(n_9321),
.Y(n_13873)
);

INVx2_ASAP7_75t_L g13874 ( 
.A(n_12001),
.Y(n_13874)
);

OA21x2_ASAP7_75t_L g13875 ( 
.A1(n_12351),
.A2(n_11446),
.B(n_11416),
.Y(n_13875)
);

BUFx8_ASAP7_75t_SL g13876 ( 
.A(n_12734),
.Y(n_13876)
);

AND2x2_ASAP7_75t_L g13877 ( 
.A(n_12341),
.B(n_10960),
.Y(n_13877)
);

INVx1_ASAP7_75t_L g13878 ( 
.A(n_12202),
.Y(n_13878)
);

INVx3_ASAP7_75t_L g13879 ( 
.A(n_11806),
.Y(n_13879)
);

INVx1_ASAP7_75t_L g13880 ( 
.A(n_12053),
.Y(n_13880)
);

AND2x2_ASAP7_75t_L g13881 ( 
.A(n_12341),
.B(n_11043),
.Y(n_13881)
);

INVx1_ASAP7_75t_L g13882 ( 
.A(n_12834),
.Y(n_13882)
);

INVx1_ASAP7_75t_L g13883 ( 
.A(n_12840),
.Y(n_13883)
);

INVx2_ASAP7_75t_L g13884 ( 
.A(n_12025),
.Y(n_13884)
);

HB1xp67_ASAP7_75t_L g13885 ( 
.A(n_12321),
.Y(n_13885)
);

AND2x2_ASAP7_75t_L g13886 ( 
.A(n_12392),
.B(n_11043),
.Y(n_13886)
);

AND2x2_ASAP7_75t_L g13887 ( 
.A(n_12392),
.B(n_11043),
.Y(n_13887)
);

AO21x2_ASAP7_75t_L g13888 ( 
.A1(n_12338),
.A2(n_12715),
.B(n_12699),
.Y(n_13888)
);

AOI22xp33_ASAP7_75t_L g13889 ( 
.A1(n_11999),
.A2(n_10749),
.B1(n_10614),
.B2(n_10746),
.Y(n_13889)
);

INVx2_ASAP7_75t_L g13890 ( 
.A(n_12033),
.Y(n_13890)
);

INVx1_ASAP7_75t_L g13891 ( 
.A(n_12845),
.Y(n_13891)
);

OAI21xp5_ASAP7_75t_L g13892 ( 
.A1(n_11968),
.A2(n_11424),
.B(n_10281),
.Y(n_13892)
);

INVx1_ASAP7_75t_SL g13893 ( 
.A(n_12842),
.Y(n_13893)
);

NAND2xp5_ASAP7_75t_L g13894 ( 
.A(n_11863),
.B(n_11634),
.Y(n_13894)
);

INVx2_ASAP7_75t_L g13895 ( 
.A(n_12044),
.Y(n_13895)
);

AO21x2_ASAP7_75t_L g13896 ( 
.A1(n_12555),
.A2(n_10840),
.B(n_10837),
.Y(n_13896)
);

INVx1_ASAP7_75t_L g13897 ( 
.A(n_12847),
.Y(n_13897)
);

AOI21xp5_ASAP7_75t_SL g13898 ( 
.A1(n_11930),
.A2(n_10803),
.B(n_10626),
.Y(n_13898)
);

HB1xp67_ASAP7_75t_L g13899 ( 
.A(n_12321),
.Y(n_13899)
);

NAND2xp5_ASAP7_75t_L g13900 ( 
.A(n_11655),
.B(n_9671),
.Y(n_13900)
);

BUFx2_ASAP7_75t_SL g13901 ( 
.A(n_12718),
.Y(n_13901)
);

INVx1_ASAP7_75t_L g13902 ( 
.A(n_12654),
.Y(n_13902)
);

AO21x2_ASAP7_75t_L g13903 ( 
.A1(n_12558),
.A2(n_12880),
.B(n_11759),
.Y(n_13903)
);

INVx2_ASAP7_75t_SL g13904 ( 
.A(n_12655),
.Y(n_13904)
);

INVx1_ASAP7_75t_L g13905 ( 
.A(n_12654),
.Y(n_13905)
);

NAND2xp5_ASAP7_75t_L g13906 ( 
.A(n_11671),
.B(n_9671),
.Y(n_13906)
);

AOI21x1_ASAP7_75t_L g13907 ( 
.A1(n_12809),
.A2(n_10849),
.B(n_10840),
.Y(n_13907)
);

INVx1_ASAP7_75t_L g13908 ( 
.A(n_12665),
.Y(n_13908)
);

INVx1_ASAP7_75t_L g13909 ( 
.A(n_12665),
.Y(n_13909)
);

INVx2_ASAP7_75t_L g13910 ( 
.A(n_12049),
.Y(n_13910)
);

HB1xp67_ASAP7_75t_L g13911 ( 
.A(n_12322),
.Y(n_13911)
);

INVx1_ASAP7_75t_L g13912 ( 
.A(n_12676),
.Y(n_13912)
);

INVx2_ASAP7_75t_L g13913 ( 
.A(n_12070),
.Y(n_13913)
);

INVx2_ASAP7_75t_L g13914 ( 
.A(n_12075),
.Y(n_13914)
);

INVx1_ASAP7_75t_L g13915 ( 
.A(n_12676),
.Y(n_13915)
);

INVx1_ASAP7_75t_L g13916 ( 
.A(n_12682),
.Y(n_13916)
);

INVx1_ASAP7_75t_L g13917 ( 
.A(n_12682),
.Y(n_13917)
);

AND2x4_ASAP7_75t_L g13918 ( 
.A(n_12655),
.B(n_12759),
.Y(n_13918)
);

BUFx6f_ASAP7_75t_L g13919 ( 
.A(n_12593),
.Y(n_13919)
);

OR2x2_ASAP7_75t_L g13920 ( 
.A(n_12704),
.B(n_9569),
.Y(n_13920)
);

INVx3_ASAP7_75t_L g13921 ( 
.A(n_11806),
.Y(n_13921)
);

INVxp33_ASAP7_75t_L g13922 ( 
.A(n_11636),
.Y(n_13922)
);

INVx1_ASAP7_75t_L g13923 ( 
.A(n_12713),
.Y(n_13923)
);

AOI21xp5_ASAP7_75t_L g13924 ( 
.A1(n_11656),
.A2(n_10749),
.B(n_10746),
.Y(n_13924)
);

OAI21x1_ASAP7_75t_L g13925 ( 
.A1(n_12711),
.A2(n_9443),
.B(n_10876),
.Y(n_13925)
);

INVx1_ASAP7_75t_SL g13926 ( 
.A(n_12853),
.Y(n_13926)
);

INVx2_ASAP7_75t_L g13927 ( 
.A(n_12079),
.Y(n_13927)
);

INVx1_ASAP7_75t_L g13928 ( 
.A(n_12713),
.Y(n_13928)
);

BUFx3_ASAP7_75t_L g13929 ( 
.A(n_12548),
.Y(n_13929)
);

INVx4_ASAP7_75t_SL g13930 ( 
.A(n_12593),
.Y(n_13930)
);

INVx1_ASAP7_75t_L g13931 ( 
.A(n_12747),
.Y(n_13931)
);

INVx1_ASAP7_75t_L g13932 ( 
.A(n_12747),
.Y(n_13932)
);

NAND2xp5_ASAP7_75t_L g13933 ( 
.A(n_11708),
.B(n_10742),
.Y(n_13933)
);

BUFx3_ASAP7_75t_L g13934 ( 
.A(n_12472),
.Y(n_13934)
);

INVx1_ASAP7_75t_L g13935 ( 
.A(n_12769),
.Y(n_13935)
);

OR2x2_ASAP7_75t_L g13936 ( 
.A(n_12720),
.B(n_9569),
.Y(n_13936)
);

HB1xp67_ASAP7_75t_L g13937 ( 
.A(n_12322),
.Y(n_13937)
);

OAI21x1_ASAP7_75t_L g13938 ( 
.A1(n_11797),
.A2(n_9443),
.B(n_10876),
.Y(n_13938)
);

INVx1_ASAP7_75t_L g13939 ( 
.A(n_12769),
.Y(n_13939)
);

AND2x2_ASAP7_75t_L g13940 ( 
.A(n_12392),
.B(n_12798),
.Y(n_13940)
);

NOR2xp67_ASAP7_75t_SL g13941 ( 
.A(n_11640),
.B(n_9888),
.Y(n_13941)
);

BUFx2_ASAP7_75t_L g13942 ( 
.A(n_12400),
.Y(n_13942)
);

AND2x2_ASAP7_75t_L g13943 ( 
.A(n_12798),
.B(n_12818),
.Y(n_13943)
);

OA21x2_ASAP7_75t_L g13944 ( 
.A1(n_12351),
.A2(n_11446),
.B(n_11416),
.Y(n_13944)
);

INVx1_ASAP7_75t_L g13945 ( 
.A(n_12777),
.Y(n_13945)
);

INVx1_ASAP7_75t_L g13946 ( 
.A(n_12777),
.Y(n_13946)
);

BUFx6f_ASAP7_75t_L g13947 ( 
.A(n_12593),
.Y(n_13947)
);

INVxp67_ASAP7_75t_L g13948 ( 
.A(n_11871),
.Y(n_13948)
);

INVx3_ASAP7_75t_L g13949 ( 
.A(n_11810),
.Y(n_13949)
);

INVx1_ASAP7_75t_L g13950 ( 
.A(n_12803),
.Y(n_13950)
);

AND2x2_ASAP7_75t_L g13951 ( 
.A(n_12798),
.B(n_11043),
.Y(n_13951)
);

OA21x2_ASAP7_75t_L g13952 ( 
.A1(n_11797),
.A2(n_11533),
.B(n_11377),
.Y(n_13952)
);

OAI21x1_ASAP7_75t_L g13953 ( 
.A1(n_12612),
.A2(n_12623),
.B(n_12706),
.Y(n_13953)
);

INVx1_ASAP7_75t_L g13954 ( 
.A(n_12803),
.Y(n_13954)
);

INVx1_ASAP7_75t_L g13955 ( 
.A(n_12814),
.Y(n_13955)
);

INVx2_ASAP7_75t_L g13956 ( 
.A(n_12112),
.Y(n_13956)
);

OA21x2_ASAP7_75t_L g13957 ( 
.A1(n_12565),
.A2(n_11533),
.B(n_11377),
.Y(n_13957)
);

INVx2_ASAP7_75t_L g13958 ( 
.A(n_12113),
.Y(n_13958)
);

AOI21x1_ASAP7_75t_L g13959 ( 
.A1(n_11871),
.A2(n_10853),
.B(n_10849),
.Y(n_13959)
);

INVx1_ASAP7_75t_L g13960 ( 
.A(n_12814),
.Y(n_13960)
);

INVx2_ASAP7_75t_L g13961 ( 
.A(n_11674),
.Y(n_13961)
);

HB1xp67_ASAP7_75t_L g13962 ( 
.A(n_12322),
.Y(n_13962)
);

INVx1_ASAP7_75t_L g13963 ( 
.A(n_12735),
.Y(n_13963)
);

HB1xp67_ASAP7_75t_L g13964 ( 
.A(n_11646),
.Y(n_13964)
);

INVx1_ASAP7_75t_L g13965 ( 
.A(n_12833),
.Y(n_13965)
);

INVx2_ASAP7_75t_L g13966 ( 
.A(n_11734),
.Y(n_13966)
);

AND2x2_ASAP7_75t_L g13967 ( 
.A(n_12818),
.B(n_12018),
.Y(n_13967)
);

INVx2_ASAP7_75t_SL g13968 ( 
.A(n_11785),
.Y(n_13968)
);

HB1xp67_ASAP7_75t_L g13969 ( 
.A(n_11646),
.Y(n_13969)
);

INVx1_ASAP7_75t_L g13970 ( 
.A(n_12833),
.Y(n_13970)
);

INVx2_ASAP7_75t_SL g13971 ( 
.A(n_11823),
.Y(n_13971)
);

INVx2_ASAP7_75t_L g13972 ( 
.A(n_11810),
.Y(n_13972)
);

INVx2_ASAP7_75t_L g13973 ( 
.A(n_11810),
.Y(n_13973)
);

BUFx2_ASAP7_75t_L g13974 ( 
.A(n_11980),
.Y(n_13974)
);

INVx1_ASAP7_75t_L g13975 ( 
.A(n_12833),
.Y(n_13975)
);

OR2x6_ASAP7_75t_L g13976 ( 
.A(n_12502),
.B(n_9888),
.Y(n_13976)
);

INVx2_ASAP7_75t_SL g13977 ( 
.A(n_12076),
.Y(n_13977)
);

INVx2_ASAP7_75t_L g13978 ( 
.A(n_12124),
.Y(n_13978)
);

HB1xp67_ASAP7_75t_L g13979 ( 
.A(n_11659),
.Y(n_13979)
);

INVx1_ASAP7_75t_L g13980 ( 
.A(n_12836),
.Y(n_13980)
);

AND2x2_ASAP7_75t_L g13981 ( 
.A(n_12818),
.B(n_11043),
.Y(n_13981)
);

AND2x2_ASAP7_75t_L g13982 ( 
.A(n_12043),
.B(n_11163),
.Y(n_13982)
);

INVx2_ASAP7_75t_SL g13983 ( 
.A(n_12139),
.Y(n_13983)
);

INVx1_ASAP7_75t_L g13984 ( 
.A(n_12836),
.Y(n_13984)
);

INVx2_ASAP7_75t_L g13985 ( 
.A(n_12269),
.Y(n_13985)
);

INVx2_ASAP7_75t_L g13986 ( 
.A(n_12801),
.Y(n_13986)
);

INVx1_ASAP7_75t_L g13987 ( 
.A(n_12836),
.Y(n_13987)
);

HB1xp67_ASAP7_75t_L g13988 ( 
.A(n_11659),
.Y(n_13988)
);

INVx2_ASAP7_75t_L g13989 ( 
.A(n_12801),
.Y(n_13989)
);

OA21x2_ASAP7_75t_L g13990 ( 
.A1(n_12281),
.A2(n_11533),
.B(n_11377),
.Y(n_13990)
);

NAND3xp33_ASAP7_75t_L g13991 ( 
.A(n_13237),
.B(n_12052),
.C(n_11923),
.Y(n_13991)
);

O2A1O1Ixp33_ASAP7_75t_L g13992 ( 
.A1(n_13237),
.A2(n_12348),
.B(n_11977),
.C(n_11876),
.Y(n_13992)
);

OA21x2_ASAP7_75t_L g13993 ( 
.A1(n_13120),
.A2(n_12282),
.B(n_12281),
.Y(n_13993)
);

AND2x2_ASAP7_75t_L g13994 ( 
.A(n_13462),
.B(n_12502),
.Y(n_13994)
);

INVx2_ASAP7_75t_L g13995 ( 
.A(n_13766),
.Y(n_13995)
);

CKINVDCx5p33_ASAP7_75t_R g13996 ( 
.A(n_13876),
.Y(n_13996)
);

AND2x4_ASAP7_75t_L g13997 ( 
.A(n_13013),
.B(n_12502),
.Y(n_13997)
);

OAI22xp5_ASAP7_75t_L g13998 ( 
.A1(n_13552),
.A2(n_12436),
.B1(n_12205),
.B2(n_12207),
.Y(n_13998)
);

OAI21xp5_ASAP7_75t_L g13999 ( 
.A1(n_13544),
.A2(n_11876),
.B(n_12231),
.Y(n_13999)
);

OAI21xp5_ASAP7_75t_L g14000 ( 
.A1(n_13544),
.A2(n_12235),
.B(n_11829),
.Y(n_14000)
);

O2A1O1Ixp33_ASAP7_75t_SL g14001 ( 
.A1(n_12964),
.A2(n_12666),
.B(n_11844),
.C(n_11649),
.Y(n_14001)
);

OAI31xp33_ASAP7_75t_SL g14002 ( 
.A1(n_13093),
.A2(n_11726),
.A3(n_11651),
.B(n_11692),
.Y(n_14002)
);

AND2x2_ASAP7_75t_L g14003 ( 
.A(n_13118),
.B(n_11976),
.Y(n_14003)
);

INVx2_ASAP7_75t_L g14004 ( 
.A(n_12916),
.Y(n_14004)
);

OAI21xp33_ASAP7_75t_SL g14005 ( 
.A1(n_13077),
.A2(n_12056),
.B(n_12480),
.Y(n_14005)
);

AND2x4_ASAP7_75t_L g14006 ( 
.A(n_13026),
.B(n_12537),
.Y(n_14006)
);

AND2x4_ASAP7_75t_L g14007 ( 
.A(n_13057),
.B(n_12646),
.Y(n_14007)
);

INVxp33_ASAP7_75t_L g14008 ( 
.A(n_13876),
.Y(n_14008)
);

AND3x1_ASAP7_75t_L g14009 ( 
.A(n_13365),
.B(n_12472),
.C(n_12649),
.Y(n_14009)
);

OAI21x1_ASAP7_75t_SL g14010 ( 
.A1(n_13303),
.A2(n_12823),
.B(n_12670),
.Y(n_14010)
);

NAND3xp33_ASAP7_75t_L g14011 ( 
.A(n_12945),
.B(n_12122),
.C(n_11855),
.Y(n_14011)
);

OR2x2_ASAP7_75t_L g14012 ( 
.A(n_13893),
.B(n_12859),
.Y(n_14012)
);

INVx1_ASAP7_75t_L g14013 ( 
.A(n_13015),
.Y(n_14013)
);

NAND2xp33_ASAP7_75t_L g14014 ( 
.A(n_13211),
.B(n_12158),
.Y(n_14014)
);

INVx2_ASAP7_75t_L g14015 ( 
.A(n_12916),
.Y(n_14015)
);

AO32x2_ASAP7_75t_L g14016 ( 
.A1(n_13401),
.A2(n_11654),
.A3(n_11663),
.B1(n_11687),
.B2(n_11805),
.Y(n_14016)
);

AOI22xp33_ASAP7_75t_SL g14017 ( 
.A1(n_12949),
.A2(n_13308),
.B1(n_12945),
.B2(n_13401),
.Y(n_14017)
);

AND2x4_ASAP7_75t_L g14018 ( 
.A(n_13067),
.B(n_13100),
.Y(n_14018)
);

AOI221xp5_ASAP7_75t_L g14019 ( 
.A1(n_13296),
.A2(n_12468),
.B1(n_11950),
.B2(n_12035),
.C(n_11947),
.Y(n_14019)
);

NAND2xp5_ASAP7_75t_L g14020 ( 
.A(n_13118),
.B(n_11738),
.Y(n_14020)
);

AOI221xp5_ASAP7_75t_L g14021 ( 
.A1(n_13296),
.A2(n_11883),
.B1(n_12288),
.B2(n_12579),
.C(n_12424),
.Y(n_14021)
);

AND2x4_ASAP7_75t_SL g14022 ( 
.A(n_13756),
.B(n_12649),
.Y(n_14022)
);

INVx1_ASAP7_75t_L g14023 ( 
.A(n_13015),
.Y(n_14023)
);

AOI22xp5_ASAP7_75t_L g14024 ( 
.A1(n_13308),
.A2(n_11743),
.B1(n_11976),
.B2(n_11693),
.Y(n_14024)
);

AND2x2_ASAP7_75t_L g14025 ( 
.A(n_13274),
.B(n_12819),
.Y(n_14025)
);

BUFx6f_ASAP7_75t_L g14026 ( 
.A(n_12941),
.Y(n_14026)
);

INVx2_ASAP7_75t_L g14027 ( 
.A(n_12918),
.Y(n_14027)
);

INVx2_ASAP7_75t_L g14028 ( 
.A(n_12918),
.Y(n_14028)
);

AOI22xp5_ASAP7_75t_L g14029 ( 
.A1(n_13365),
.A2(n_11932),
.B1(n_11831),
.B2(n_12487),
.Y(n_14029)
);

AO32x2_ASAP7_75t_L g14030 ( 
.A1(n_13968),
.A2(n_11676),
.A3(n_11704),
.B1(n_11696),
.B2(n_12547),
.Y(n_14030)
);

AND2x2_ASAP7_75t_L g14031 ( 
.A(n_13274),
.B(n_12737),
.Y(n_14031)
);

BUFx12f_ASAP7_75t_L g14032 ( 
.A(n_13549),
.Y(n_14032)
);

BUFx6f_ASAP7_75t_L g14033 ( 
.A(n_12941),
.Y(n_14033)
);

OAI21xp5_ASAP7_75t_L g14034 ( 
.A1(n_13077),
.A2(n_11924),
.B(n_11842),
.Y(n_14034)
);

AND2x4_ASAP7_75t_L g14035 ( 
.A(n_13100),
.B(n_12750),
.Y(n_14035)
);

AND2x2_ASAP7_75t_L g14036 ( 
.A(n_13901),
.B(n_12737),
.Y(n_14036)
);

OA21x2_ASAP7_75t_L g14037 ( 
.A1(n_13120),
.A2(n_12282),
.B(n_12037),
.Y(n_14037)
);

OAI22xp5_ASAP7_75t_L g14038 ( 
.A1(n_13552),
.A2(n_12205),
.B1(n_12207),
.B2(n_12145),
.Y(n_14038)
);

AND2x2_ASAP7_75t_L g14039 ( 
.A(n_12964),
.B(n_13466),
.Y(n_14039)
);

AND2x2_ASAP7_75t_L g14040 ( 
.A(n_13471),
.B(n_12439),
.Y(n_14040)
);

AND2x2_ASAP7_75t_L g14041 ( 
.A(n_13474),
.B(n_12253),
.Y(n_14041)
);

AND2x2_ASAP7_75t_L g14042 ( 
.A(n_13363),
.B(n_12260),
.Y(n_14042)
);

OAI21x1_ASAP7_75t_L g14043 ( 
.A1(n_12917),
.A2(n_12810),
.B(n_12712),
.Y(n_14043)
);

INVx2_ASAP7_75t_L g14044 ( 
.A(n_12924),
.Y(n_14044)
);

NAND2xp5_ASAP7_75t_L g14045 ( 
.A(n_12998),
.B(n_11755),
.Y(n_14045)
);

INVx1_ASAP7_75t_L g14046 ( 
.A(n_13018),
.Y(n_14046)
);

NAND4xp25_ASAP7_75t_SL g14047 ( 
.A(n_13898),
.B(n_12305),
.C(n_11721),
.D(n_12324),
.Y(n_14047)
);

INVx1_ASAP7_75t_L g14048 ( 
.A(n_13018),
.Y(n_14048)
);

AND2x4_ASAP7_75t_L g14049 ( 
.A(n_13112),
.B(n_12924),
.Y(n_14049)
);

AND2x4_ASAP7_75t_L g14050 ( 
.A(n_13112),
.B(n_8183),
.Y(n_14050)
);

AOI221xp5_ASAP7_75t_L g14051 ( 
.A1(n_13688),
.A2(n_12115),
.B1(n_12111),
.B2(n_11924),
.C(n_11827),
.Y(n_14051)
);

AND2x4_ASAP7_75t_L g14052 ( 
.A(n_12936),
.B(n_12602),
.Y(n_14052)
);

OAI21x1_ASAP7_75t_L g14053 ( 
.A1(n_12932),
.A2(n_12850),
.B(n_12843),
.Y(n_14053)
);

OA21x2_ASAP7_75t_L g14054 ( 
.A1(n_12921),
.A2(n_12037),
.B(n_11961),
.Y(n_14054)
);

AOI21x1_ASAP7_75t_L g14055 ( 
.A1(n_12921),
.A2(n_11862),
.B(n_11832),
.Y(n_14055)
);

O2A1O1Ixp33_ASAP7_75t_L g14056 ( 
.A1(n_13948),
.A2(n_11638),
.B(n_12510),
.C(n_12754),
.Y(n_14056)
);

AOI22xp5_ASAP7_75t_L g14057 ( 
.A1(n_13903),
.A2(n_13622),
.B1(n_13358),
.B2(n_13396),
.Y(n_14057)
);

AND2x2_ASAP7_75t_L g14058 ( 
.A(n_13383),
.B(n_12278),
.Y(n_14058)
);

AND2x2_ASAP7_75t_L g14059 ( 
.A(n_13392),
.B(n_12286),
.Y(n_14059)
);

AOI21xp5_ASAP7_75t_L g14060 ( 
.A1(n_13062),
.A2(n_11912),
.B(n_11898),
.Y(n_14060)
);

OAI21xp5_ASAP7_75t_L g14061 ( 
.A1(n_13165),
.A2(n_11881),
.B(n_11949),
.Y(n_14061)
);

INVx1_ASAP7_75t_L g14062 ( 
.A(n_13060),
.Y(n_14062)
);

AND2x2_ASAP7_75t_L g14063 ( 
.A(n_13358),
.B(n_12295),
.Y(n_14063)
);

AND2x2_ASAP7_75t_L g14064 ( 
.A(n_13396),
.B(n_12302),
.Y(n_14064)
);

AO32x1_ASAP7_75t_L g14065 ( 
.A1(n_13904),
.A2(n_11707),
.A3(n_11733),
.B1(n_12458),
.B2(n_12457),
.Y(n_14065)
);

INVx1_ASAP7_75t_L g14066 ( 
.A(n_13060),
.Y(n_14066)
);

INVx1_ASAP7_75t_L g14067 ( 
.A(n_13075),
.Y(n_14067)
);

CKINVDCx6p67_ASAP7_75t_R g14068 ( 
.A(n_13254),
.Y(n_14068)
);

AO21x2_ASAP7_75t_L g14069 ( 
.A1(n_12934),
.A2(n_12860),
.B(n_12880),
.Y(n_14069)
);

AOI22x1_ASAP7_75t_SL g14070 ( 
.A1(n_13211),
.A2(n_8757),
.B1(n_12763),
.B2(n_11892),
.Y(n_14070)
);

CKINVDCx9p33_ASAP7_75t_R g14071 ( 
.A(n_13283),
.Y(n_14071)
);

CKINVDCx20_ASAP7_75t_R g14072 ( 
.A(n_13549),
.Y(n_14072)
);

NOR2x1_ASAP7_75t_SL g14073 ( 
.A(n_13413),
.B(n_10626),
.Y(n_14073)
);

INVx1_ASAP7_75t_L g14074 ( 
.A(n_13075),
.Y(n_14074)
);

OAI21x1_ASAP7_75t_L g14075 ( 
.A1(n_13267),
.A2(n_12904),
.B(n_12872),
.Y(n_14075)
);

AND2x2_ASAP7_75t_L g14076 ( 
.A(n_12936),
.B(n_12303),
.Y(n_14076)
);

INVxp67_ASAP7_75t_L g14077 ( 
.A(n_13101),
.Y(n_14077)
);

A2O1A1Ixp33_ASAP7_75t_L g14078 ( 
.A1(n_13922),
.A2(n_13062),
.B(n_13762),
.C(n_13721),
.Y(n_14078)
);

OR2x2_ASAP7_75t_L g14079 ( 
.A(n_13893),
.B(n_13926),
.Y(n_14079)
);

NAND2xp33_ASAP7_75t_L g14080 ( 
.A(n_13427),
.B(n_11845),
.Y(n_14080)
);

INVx1_ASAP7_75t_L g14081 ( 
.A(n_13083),
.Y(n_14081)
);

BUFx4f_ASAP7_75t_SL g14082 ( 
.A(n_13807),
.Y(n_14082)
);

INVx1_ASAP7_75t_L g14083 ( 
.A(n_13083),
.Y(n_14083)
);

NAND2xp5_ASAP7_75t_L g14084 ( 
.A(n_13000),
.B(n_11770),
.Y(n_14084)
);

AO32x2_ASAP7_75t_L g14085 ( 
.A1(n_13971),
.A2(n_11885),
.A3(n_11917),
.B1(n_12470),
.B2(n_11901),
.Y(n_14085)
);

OA21x2_ASAP7_75t_L g14086 ( 
.A1(n_12934),
.A2(n_11961),
.B(n_12111),
.Y(n_14086)
);

AND2x2_ASAP7_75t_L g14087 ( 
.A(n_13256),
.B(n_12308),
.Y(n_14087)
);

OR2x2_ASAP7_75t_L g14088 ( 
.A(n_13926),
.B(n_12861),
.Y(n_14088)
);

INVx1_ASAP7_75t_L g14089 ( 
.A(n_13091),
.Y(n_14089)
);

NAND4xp25_ASAP7_75t_L g14090 ( 
.A(n_13768),
.B(n_12115),
.C(n_11841),
.D(n_12423),
.Y(n_14090)
);

AND2x2_ASAP7_75t_L g14091 ( 
.A(n_13256),
.B(n_12311),
.Y(n_14091)
);

INVxp67_ASAP7_75t_L g14092 ( 
.A(n_13362),
.Y(n_14092)
);

INVx1_ASAP7_75t_L g14093 ( 
.A(n_13091),
.Y(n_14093)
);

AND2x4_ASAP7_75t_L g14094 ( 
.A(n_13189),
.B(n_12719),
.Y(n_14094)
);

AND2x2_ASAP7_75t_L g14095 ( 
.A(n_13458),
.B(n_12315),
.Y(n_14095)
);

AO32x2_ASAP7_75t_L g14096 ( 
.A1(n_13977),
.A2(n_12233),
.A3(n_11910),
.B1(n_12394),
.B2(n_12387),
.Y(n_14096)
);

INVx4_ASAP7_75t_L g14097 ( 
.A(n_12940),
.Y(n_14097)
);

AND2x2_ASAP7_75t_L g14098 ( 
.A(n_13458),
.B(n_12318),
.Y(n_14098)
);

OR2x2_ASAP7_75t_L g14099 ( 
.A(n_13269),
.B(n_11768),
.Y(n_14099)
);

AND2x4_ASAP7_75t_L g14100 ( 
.A(n_13189),
.B(n_12319),
.Y(n_14100)
);

NAND2xp5_ASAP7_75t_L g14101 ( 
.A(n_13869),
.B(n_11812),
.Y(n_14101)
);

OAI21xp5_ASAP7_75t_L g14102 ( 
.A1(n_13165),
.A2(n_11809),
.B(n_11853),
.Y(n_14102)
);

A2O1A1Ixp33_ASAP7_75t_L g14103 ( 
.A1(n_13922),
.A2(n_11780),
.B(n_11775),
.C(n_11841),
.Y(n_14103)
);

AND2x4_ASAP7_75t_L g14104 ( 
.A(n_13242),
.B(n_12323),
.Y(n_14104)
);

NAND4xp25_ASAP7_75t_L g14105 ( 
.A(n_13768),
.B(n_12410),
.C(n_12089),
.D(n_12629),
.Y(n_14105)
);

INVx4_ASAP7_75t_L g14106 ( 
.A(n_12940),
.Y(n_14106)
);

AND2x2_ASAP7_75t_L g14107 ( 
.A(n_13459),
.B(n_12554),
.Y(n_14107)
);

CKINVDCx20_ASAP7_75t_R g14108 ( 
.A(n_13038),
.Y(n_14108)
);

NOR2xp33_ASAP7_75t_L g14109 ( 
.A(n_13427),
.B(n_8757),
.Y(n_14109)
);

NAND2xp5_ASAP7_75t_L g14110 ( 
.A(n_13869),
.B(n_11821),
.Y(n_14110)
);

AND2x2_ASAP7_75t_L g14111 ( 
.A(n_13459),
.B(n_12566),
.Y(n_14111)
);

OR2x2_ASAP7_75t_L g14112 ( 
.A(n_13644),
.B(n_11792),
.Y(n_14112)
);

HB1xp67_ASAP7_75t_L g14113 ( 
.A(n_13109),
.Y(n_14113)
);

NOR2x1_ASAP7_75t_SL g14114 ( 
.A(n_13413),
.B(n_13541),
.Y(n_14114)
);

OAI21xp5_ASAP7_75t_L g14115 ( 
.A1(n_13438),
.A2(n_12291),
.B(n_12402),
.Y(n_14115)
);

AND2x2_ASAP7_75t_L g14116 ( 
.A(n_13014),
.B(n_12587),
.Y(n_14116)
);

AO21x2_ASAP7_75t_L g14117 ( 
.A1(n_12937),
.A2(n_11844),
.B(n_12510),
.Y(n_14117)
);

A2O1A1Ixp33_ASAP7_75t_L g14118 ( 
.A1(n_13762),
.A2(n_11739),
.B(n_12410),
.C(n_12402),
.Y(n_14118)
);

OR2x6_ASAP7_75t_L g14119 ( 
.A(n_13188),
.B(n_13242),
.Y(n_14119)
);

AND2x2_ASAP7_75t_L g14120 ( 
.A(n_13017),
.B(n_12600),
.Y(n_14120)
);

AND2x2_ASAP7_75t_L g14121 ( 
.A(n_13175),
.B(n_12608),
.Y(n_14121)
);

OAI22xp5_ASAP7_75t_L g14122 ( 
.A1(n_13129),
.A2(n_12145),
.B1(n_12298),
.B2(n_11649),
.Y(n_14122)
);

AND2x2_ASAP7_75t_L g14123 ( 
.A(n_13342),
.B(n_12611),
.Y(n_14123)
);

A2O1A1Ixp33_ASAP7_75t_L g14124 ( 
.A1(n_13688),
.A2(n_12147),
.B(n_12098),
.C(n_12754),
.Y(n_14124)
);

AND2x4_ASAP7_75t_L g14125 ( 
.A(n_13307),
.B(n_12874),
.Y(n_14125)
);

AND2x2_ASAP7_75t_L g14126 ( 
.A(n_13301),
.B(n_12617),
.Y(n_14126)
);

O2A1O1Ixp33_ASAP7_75t_L g14127 ( 
.A1(n_13948),
.A2(n_12709),
.B(n_11757),
.C(n_12067),
.Y(n_14127)
);

AND2x2_ASAP7_75t_L g14128 ( 
.A(n_13355),
.B(n_12620),
.Y(n_14128)
);

HB1xp67_ASAP7_75t_L g14129 ( 
.A(n_13109),
.Y(n_14129)
);

INVx3_ASAP7_75t_L g14130 ( 
.A(n_13352),
.Y(n_14130)
);

NAND2xp5_ASAP7_75t_L g14131 ( 
.A(n_13644),
.B(n_12752),
.Y(n_14131)
);

AOI221x1_ASAP7_75t_SL g14132 ( 
.A1(n_13622),
.A2(n_13129),
.B1(n_12969),
.B2(n_13400),
.C(n_13235),
.Y(n_14132)
);

OAI21xp5_ASAP7_75t_L g14133 ( 
.A1(n_13438),
.A2(n_12672),
.B(n_12660),
.Y(n_14133)
);

AND2x4_ASAP7_75t_L g14134 ( 
.A(n_13307),
.B(n_12939),
.Y(n_14134)
);

AND2x2_ASAP7_75t_L g14135 ( 
.A(n_13526),
.B(n_12627),
.Y(n_14135)
);

AND2x4_ASAP7_75t_L g14136 ( 
.A(n_12942),
.B(n_11163),
.Y(n_14136)
);

OAI21x1_ASAP7_75t_L g14137 ( 
.A1(n_12981),
.A2(n_12114),
.B(n_12101),
.Y(n_14137)
);

AND2x4_ASAP7_75t_L g14138 ( 
.A(n_13152),
.B(n_11163),
.Y(n_14138)
);

INVx2_ASAP7_75t_L g14139 ( 
.A(n_13352),
.Y(n_14139)
);

INVx1_ASAP7_75t_L g14140 ( 
.A(n_13116),
.Y(n_14140)
);

AND2x2_ASAP7_75t_L g14141 ( 
.A(n_13576),
.B(n_12628),
.Y(n_14141)
);

O2A1O1Ixp33_ASAP7_75t_L g14142 ( 
.A1(n_13721),
.A2(n_12709),
.B(n_11757),
.C(n_12067),
.Y(n_14142)
);

NAND4xp25_ASAP7_75t_L g14143 ( 
.A(n_13596),
.B(n_12639),
.C(n_12637),
.D(n_12344),
.Y(n_14143)
);

NAND2xp5_ASAP7_75t_L g14144 ( 
.A(n_13683),
.B(n_12762),
.Y(n_14144)
);

INVx1_ASAP7_75t_L g14145 ( 
.A(n_13116),
.Y(n_14145)
);

BUFx6f_ASAP7_75t_L g14146 ( 
.A(n_12962),
.Y(n_14146)
);

AND2x2_ASAP7_75t_SL g14147 ( 
.A(n_13304),
.B(n_11862),
.Y(n_14147)
);

NOR2xp33_ASAP7_75t_L g14148 ( 
.A(n_12966),
.B(n_11798),
.Y(n_14148)
);

INVx2_ASAP7_75t_L g14149 ( 
.A(n_13361),
.Y(n_14149)
);

AOI221xp5_ASAP7_75t_L g14150 ( 
.A1(n_12909),
.A2(n_11723),
.B1(n_12310),
.B2(n_12631),
.C(n_12263),
.Y(n_14150)
);

NOR2xp33_ASAP7_75t_L g14151 ( 
.A(n_12966),
.B(n_10460),
.Y(n_14151)
);

O2A1O1Ixp33_ASAP7_75t_L g14152 ( 
.A1(n_12947),
.A2(n_11795),
.B(n_11813),
.C(n_12298),
.Y(n_14152)
);

INVx1_ASAP7_75t_L g14153 ( 
.A(n_13133),
.Y(n_14153)
);

OR2x6_ASAP7_75t_L g14154 ( 
.A(n_13188),
.B(n_11762),
.Y(n_14154)
);

OAI21xp5_ASAP7_75t_L g14155 ( 
.A1(n_13924),
.A2(n_11661),
.B(n_11697),
.Y(n_14155)
);

NOR2xp33_ASAP7_75t_L g14156 ( 
.A(n_12972),
.B(n_10460),
.Y(n_14156)
);

OR2x2_ASAP7_75t_L g14157 ( 
.A(n_13683),
.B(n_11750),
.Y(n_14157)
);

INVx1_ASAP7_75t_L g14158 ( 
.A(n_13133),
.Y(n_14158)
);

AND2x2_ASAP7_75t_L g14159 ( 
.A(n_12946),
.B(n_12636),
.Y(n_14159)
);

AND2x2_ASAP7_75t_L g14160 ( 
.A(n_12967),
.B(n_12641),
.Y(n_14160)
);

NOR2x1_ASAP7_75t_SL g14161 ( 
.A(n_13413),
.B(n_9888),
.Y(n_14161)
);

NAND2xp5_ASAP7_75t_L g14162 ( 
.A(n_13520),
.B(n_12775),
.Y(n_14162)
);

OR2x2_ASAP7_75t_L g14163 ( 
.A(n_13933),
.B(n_11761),
.Y(n_14163)
);

AND2x2_ASAP7_75t_L g14164 ( 
.A(n_12985),
.B(n_12656),
.Y(n_14164)
);

OR2x2_ASAP7_75t_L g14165 ( 
.A(n_13933),
.B(n_11880),
.Y(n_14165)
);

AND2x4_ASAP7_75t_L g14166 ( 
.A(n_13157),
.B(n_13224),
.Y(n_14166)
);

OAI22xp5_ASAP7_75t_L g14167 ( 
.A1(n_12969),
.A2(n_12630),
.B1(n_12661),
.B2(n_12378),
.Y(n_14167)
);

A2O1A1Ixp33_ASAP7_75t_L g14168 ( 
.A1(n_13442),
.A2(n_12643),
.B(n_12716),
.C(n_12128),
.Y(n_14168)
);

OR2x2_ASAP7_75t_L g14169 ( 
.A(n_13733),
.B(n_11895),
.Y(n_14169)
);

OAI22xp5_ASAP7_75t_L g14170 ( 
.A1(n_13400),
.A2(n_12630),
.B1(n_12661),
.B2(n_12378),
.Y(n_14170)
);

AND2x2_ASAP7_75t_L g14171 ( 
.A(n_13007),
.B(n_12681),
.Y(n_14171)
);

AO21x1_ASAP7_75t_L g14172 ( 
.A1(n_12937),
.A2(n_13885),
.B(n_13834),
.Y(n_14172)
);

AND2x2_ASAP7_75t_L g14173 ( 
.A(n_13393),
.B(n_12689),
.Y(n_14173)
);

OAI22xp5_ASAP7_75t_L g14174 ( 
.A1(n_13235),
.A2(n_12382),
.B1(n_12198),
.B2(n_11813),
.Y(n_14174)
);

NAND2xp5_ASAP7_75t_L g14175 ( 
.A(n_13520),
.B(n_13734),
.Y(n_14175)
);

INVx2_ASAP7_75t_L g14176 ( 
.A(n_13361),
.Y(n_14176)
);

AND2x2_ASAP7_75t_L g14177 ( 
.A(n_13402),
.B(n_11741),
.Y(n_14177)
);

AND2x2_ASAP7_75t_L g14178 ( 
.A(n_13405),
.B(n_11843),
.Y(n_14178)
);

BUFx2_ASAP7_75t_L g14179 ( 
.A(n_13127),
.Y(n_14179)
);

AND2x2_ASAP7_75t_L g14180 ( 
.A(n_13484),
.B(n_11163),
.Y(n_14180)
);

HB1xp67_ASAP7_75t_L g14181 ( 
.A(n_12950),
.Y(n_14181)
);

AND2x2_ASAP7_75t_L g14182 ( 
.A(n_13492),
.B(n_11163),
.Y(n_14182)
);

BUFx12f_ASAP7_75t_L g14183 ( 
.A(n_12940),
.Y(n_14183)
);

A2O1A1Ixp33_ASAP7_75t_L g14184 ( 
.A1(n_13442),
.A2(n_12128),
.B(n_12191),
.C(n_12175),
.Y(n_14184)
);

AND2x2_ASAP7_75t_L g14185 ( 
.A(n_13037),
.B(n_11205),
.Y(n_14185)
);

INVx2_ASAP7_75t_L g14186 ( 
.A(n_12977),
.Y(n_14186)
);

AND2x4_ASAP7_75t_L g14187 ( 
.A(n_13246),
.B(n_11205),
.Y(n_14187)
);

AND2x2_ASAP7_75t_L g14188 ( 
.A(n_13037),
.B(n_11205),
.Y(n_14188)
);

AND2x2_ASAP7_75t_L g14189 ( 
.A(n_13841),
.B(n_11205),
.Y(n_14189)
);

AOI221xp5_ASAP7_75t_L g14190 ( 
.A1(n_12909),
.A2(n_12276),
.B1(n_12509),
.B2(n_12583),
.C(n_12581),
.Y(n_14190)
);

A2O1A1Ixp33_ASAP7_75t_L g14191 ( 
.A1(n_13924),
.A2(n_12560),
.B(n_12518),
.C(n_12817),
.Y(n_14191)
);

AND2x2_ASAP7_75t_L g14192 ( 
.A(n_13841),
.B(n_11205),
.Y(n_14192)
);

AOI22xp5_ASAP7_75t_L g14193 ( 
.A1(n_13903),
.A2(n_13105),
.B1(n_12972),
.B2(n_13335),
.Y(n_14193)
);

AND2x2_ASAP7_75t_L g14194 ( 
.A(n_13929),
.B(n_13481),
.Y(n_14194)
);

AND2x2_ASAP7_75t_L g14195 ( 
.A(n_13430),
.B(n_11238),
.Y(n_14195)
);

NOR2xp33_ASAP7_75t_L g14196 ( 
.A(n_13127),
.B(n_10460),
.Y(n_14196)
);

INVx1_ASAP7_75t_L g14197 ( 
.A(n_12950),
.Y(n_14197)
);

AO21x2_ASAP7_75t_L g14198 ( 
.A1(n_13335),
.A2(n_12666),
.B(n_12504),
.Y(n_14198)
);

OAI22xp5_ASAP7_75t_SL g14199 ( 
.A1(n_13651),
.A2(n_11862),
.B1(n_9984),
.B2(n_10086),
.Y(n_14199)
);

AND2x2_ASAP7_75t_L g14200 ( 
.A(n_13105),
.B(n_11238),
.Y(n_14200)
);

OR2x2_ASAP7_75t_L g14201 ( 
.A(n_13558),
.B(n_11630),
.Y(n_14201)
);

AND2x2_ASAP7_75t_L g14202 ( 
.A(n_13218),
.B(n_13096),
.Y(n_14202)
);

OR2x2_ASAP7_75t_L g14203 ( 
.A(n_13564),
.B(n_11632),
.Y(n_14203)
);

AND2x2_ASAP7_75t_L g14204 ( 
.A(n_13115),
.B(n_11238),
.Y(n_14204)
);

A2O1A1Ixp33_ASAP7_75t_L g14205 ( 
.A1(n_13941),
.A2(n_12892),
.B(n_12507),
.C(n_12464),
.Y(n_14205)
);

AND2x4_ASAP7_75t_L g14206 ( 
.A(n_13258),
.B(n_11238),
.Y(n_14206)
);

BUFx2_ASAP7_75t_L g14207 ( 
.A(n_13380),
.Y(n_14207)
);

OAI21xp5_ASAP7_75t_L g14208 ( 
.A1(n_13806),
.A2(n_12109),
.B(n_12108),
.Y(n_14208)
);

OAI22xp5_ASAP7_75t_L g14209 ( 
.A1(n_12927),
.A2(n_12382),
.B1(n_12198),
.B2(n_11795),
.Y(n_14209)
);

AND2x4_ASAP7_75t_L g14210 ( 
.A(n_13327),
.B(n_11238),
.Y(n_14210)
);

NAND3xp33_ASAP7_75t_L g14211 ( 
.A(n_13201),
.B(n_11969),
.C(n_11840),
.Y(n_14211)
);

INVxp67_ASAP7_75t_L g14212 ( 
.A(n_13607),
.Y(n_14212)
);

CKINVDCx6p67_ASAP7_75t_R g14213 ( 
.A(n_13518),
.Y(n_14213)
);

A2O1A1Ixp33_ASAP7_75t_L g14214 ( 
.A1(n_13093),
.A2(n_12200),
.B(n_12171),
.C(n_12575),
.Y(n_14214)
);

OA21x2_ASAP7_75t_L g14215 ( 
.A1(n_13834),
.A2(n_11778),
.B(n_11749),
.Y(n_14215)
);

AOI22x1_ASAP7_75t_SL g14216 ( 
.A1(n_13756),
.A2(n_10049),
.B1(n_10106),
.B2(n_10012),
.Y(n_14216)
);

OAI21xp5_ASAP7_75t_L g14217 ( 
.A1(n_13099),
.A2(n_12109),
.B(n_12108),
.Y(n_14217)
);

AND2x4_ASAP7_75t_L g14218 ( 
.A(n_13407),
.B(n_11299),
.Y(n_14218)
);

O2A1O1Ixp33_ASAP7_75t_L g14219 ( 
.A1(n_12947),
.A2(n_12680),
.B(n_12678),
.C(n_12406),
.Y(n_14219)
);

NAND2xp5_ASAP7_75t_L g14220 ( 
.A(n_13567),
.B(n_12815),
.Y(n_14220)
);

AND2x2_ASAP7_75t_L g14221 ( 
.A(n_13410),
.B(n_11299),
.Y(n_14221)
);

OAI21xp5_ASAP7_75t_L g14222 ( 
.A1(n_13099),
.A2(n_12927),
.B(n_13892),
.Y(n_14222)
);

OR2x2_ASAP7_75t_L g14223 ( 
.A(n_13702),
.B(n_12294),
.Y(n_14223)
);

AO32x2_ASAP7_75t_L g14224 ( 
.A1(n_13983),
.A2(n_12361),
.A3(n_12280),
.B1(n_12309),
.B2(n_11971),
.Y(n_14224)
);

INVx2_ASAP7_75t_L g14225 ( 
.A(n_12977),
.Y(n_14225)
);

INVx1_ASAP7_75t_L g14226 ( 
.A(n_12958),
.Y(n_14226)
);

A2O1A1Ixp33_ASAP7_75t_L g14227 ( 
.A1(n_13463),
.A2(n_12171),
.B(n_12200),
.C(n_12530),
.Y(n_14227)
);

AND2x2_ASAP7_75t_L g14228 ( 
.A(n_13435),
.B(n_11299),
.Y(n_14228)
);

AND2x4_ASAP7_75t_L g14229 ( 
.A(n_13040),
.B(n_11299),
.Y(n_14229)
);

AND2x4_ASAP7_75t_L g14230 ( 
.A(n_13040),
.B(n_11299),
.Y(n_14230)
);

AND2x2_ASAP7_75t_L g14231 ( 
.A(n_12938),
.B(n_11315),
.Y(n_14231)
);

INVx2_ASAP7_75t_L g14232 ( 
.A(n_12977),
.Y(n_14232)
);

AND2x2_ASAP7_75t_L g14233 ( 
.A(n_12938),
.B(n_11315),
.Y(n_14233)
);

AND2x4_ASAP7_75t_L g14234 ( 
.A(n_13043),
.B(n_11315),
.Y(n_14234)
);

INVx1_ASAP7_75t_L g14235 ( 
.A(n_12958),
.Y(n_14235)
);

OR2x2_ASAP7_75t_L g14236 ( 
.A(n_13706),
.B(n_12519),
.Y(n_14236)
);

NAND2xp5_ASAP7_75t_L g14237 ( 
.A(n_13882),
.B(n_12486),
.Y(n_14237)
);

AND2x2_ASAP7_75t_L g14238 ( 
.A(n_12938),
.B(n_11315),
.Y(n_14238)
);

AND2x4_ASAP7_75t_SL g14239 ( 
.A(n_13038),
.B(n_9608),
.Y(n_14239)
);

OR2x2_ASAP7_75t_L g14240 ( 
.A(n_13707),
.B(n_12520),
.Y(n_14240)
);

AO21x2_ASAP7_75t_L g14241 ( 
.A1(n_13885),
.A2(n_12616),
.B(n_12799),
.Y(n_14241)
);

AND2x2_ASAP7_75t_L g14242 ( 
.A(n_12992),
.B(n_11315),
.Y(n_14242)
);

INVx1_ASAP7_75t_L g14243 ( 
.A(n_12965),
.Y(n_14243)
);

NAND2xp5_ASAP7_75t_L g14244 ( 
.A(n_13883),
.B(n_12508),
.Y(n_14244)
);

INVx1_ASAP7_75t_L g14245 ( 
.A(n_12965),
.Y(n_14245)
);

HB1xp67_ASAP7_75t_L g14246 ( 
.A(n_12970),
.Y(n_14246)
);

INVx2_ASAP7_75t_L g14247 ( 
.A(n_13146),
.Y(n_14247)
);

AND2x2_ASAP7_75t_L g14248 ( 
.A(n_13184),
.B(n_11344),
.Y(n_14248)
);

BUFx3_ASAP7_75t_L g14249 ( 
.A(n_13573),
.Y(n_14249)
);

OAI211xp5_ASAP7_75t_L g14250 ( 
.A1(n_13201),
.A2(n_12871),
.B(n_12883),
.C(n_12531),
.Y(n_14250)
);

INVxp67_ASAP7_75t_L g14251 ( 
.A(n_13607),
.Y(n_14251)
);

AND2x4_ASAP7_75t_L g14252 ( 
.A(n_13043),
.B(n_11344),
.Y(n_14252)
);

INVx1_ASAP7_75t_L g14253 ( 
.A(n_12970),
.Y(n_14253)
);

BUFx10_ASAP7_75t_L g14254 ( 
.A(n_13146),
.Y(n_14254)
);

OA21x2_ASAP7_75t_L g14255 ( 
.A1(n_13899),
.A2(n_13937),
.B(n_13911),
.Y(n_14255)
);

O2A1O1Ixp5_ASAP7_75t_L g14256 ( 
.A1(n_13586),
.A2(n_12659),
.B(n_12668),
.C(n_12625),
.Y(n_14256)
);

AOI221xp5_ASAP7_75t_L g14257 ( 
.A1(n_13349),
.A2(n_12746),
.B1(n_12795),
.B2(n_11944),
.C(n_12743),
.Y(n_14257)
);

NAND2xp5_ASAP7_75t_L g14258 ( 
.A(n_13891),
.B(n_11946),
.Y(n_14258)
);

AO32x2_ASAP7_75t_L g14259 ( 
.A1(n_13769),
.A2(n_11970),
.A3(n_12574),
.B1(n_12441),
.B2(n_12571),
.Y(n_14259)
);

BUFx2_ASAP7_75t_L g14260 ( 
.A(n_13380),
.Y(n_14260)
);

NAND2xp5_ASAP7_75t_L g14261 ( 
.A(n_13897),
.B(n_12867),
.Y(n_14261)
);

O2A1O1Ixp33_ASAP7_75t_L g14262 ( 
.A1(n_13012),
.A2(n_12494),
.B(n_12675),
.C(n_12607),
.Y(n_14262)
);

INVx1_ASAP7_75t_L g14263 ( 
.A(n_12976),
.Y(n_14263)
);

INVx1_ASAP7_75t_L g14264 ( 
.A(n_12976),
.Y(n_14264)
);

NOR2xp33_ASAP7_75t_L g14265 ( 
.A(n_13061),
.B(n_10460),
.Y(n_14265)
);

AND2x2_ASAP7_75t_SL g14266 ( 
.A(n_13304),
.B(n_8546),
.Y(n_14266)
);

INVxp67_ASAP7_75t_L g14267 ( 
.A(n_13283),
.Y(n_14267)
);

NOR2xp33_ASAP7_75t_SL g14268 ( 
.A(n_12956),
.B(n_9968),
.Y(n_14268)
);

NAND4xp25_ASAP7_75t_L g14269 ( 
.A(n_13596),
.B(n_12776),
.C(n_12858),
.D(n_12829),
.Y(n_14269)
);

A2O1A1Ixp33_ASAP7_75t_L g14270 ( 
.A1(n_13463),
.A2(n_12782),
.B(n_12794),
.C(n_12863),
.Y(n_14270)
);

AND2x2_ASAP7_75t_L g14271 ( 
.A(n_13184),
.B(n_11344),
.Y(n_14271)
);

OAI21xp5_ASAP7_75t_L g14272 ( 
.A1(n_13892),
.A2(n_12494),
.B(n_12114),
.Y(n_14272)
);

AO21x2_ASAP7_75t_L g14273 ( 
.A1(n_13899),
.A2(n_12404),
.B(n_12399),
.Y(n_14273)
);

AOI21xp5_ASAP7_75t_L g14274 ( 
.A1(n_13056),
.A2(n_11763),
.B(n_12101),
.Y(n_14274)
);

AO21x2_ASAP7_75t_L g14275 ( 
.A1(n_13911),
.A2(n_11680),
.B(n_11668),
.Y(n_14275)
);

AOI21xp5_ASAP7_75t_L g14276 ( 
.A1(n_13056),
.A2(n_12429),
.B(n_12427),
.Y(n_14276)
);

O2A1O1Ixp33_ASAP7_75t_SL g14277 ( 
.A1(n_13012),
.A2(n_12902),
.B(n_12431),
.C(n_12398),
.Y(n_14277)
);

AO32x2_ASAP7_75t_L g14278 ( 
.A1(n_13354),
.A2(n_11918),
.A3(n_12258),
.B1(n_11850),
.B2(n_13832),
.Y(n_14278)
);

AND2x2_ASAP7_75t_L g14279 ( 
.A(n_13204),
.B(n_11344),
.Y(n_14279)
);

AND2x2_ASAP7_75t_L g14280 ( 
.A(n_13204),
.B(n_11344),
.Y(n_14280)
);

INVx5_ASAP7_75t_SL g14281 ( 
.A(n_13222),
.Y(n_14281)
);

INVx1_ASAP7_75t_L g14282 ( 
.A(n_12996),
.Y(n_14282)
);

AND2x4_ASAP7_75t_L g14283 ( 
.A(n_13830),
.B(n_11498),
.Y(n_14283)
);

OR2x6_ASAP7_75t_L g14284 ( 
.A(n_13532),
.B(n_9968),
.Y(n_14284)
);

AOI21xp5_ASAP7_75t_SL g14285 ( 
.A1(n_12956),
.A2(n_12592),
.B(n_12773),
.Y(n_14285)
);

AOI21x1_ASAP7_75t_L g14286 ( 
.A1(n_13937),
.A2(n_12726),
.B(n_12778),
.Y(n_14286)
);

OA21x2_ASAP7_75t_L g14287 ( 
.A1(n_13962),
.A2(n_11778),
.B(n_11749),
.Y(n_14287)
);

AOI21xp5_ASAP7_75t_SL g14288 ( 
.A1(n_13651),
.A2(n_12779),
.B(n_12714),
.Y(n_14288)
);

OAI211xp5_ASAP7_75t_L g14289 ( 
.A1(n_13349),
.A2(n_12894),
.B(n_12355),
.C(n_12866),
.Y(n_14289)
);

AND2x2_ASAP7_75t_L g14290 ( 
.A(n_13321),
.B(n_11498),
.Y(n_14290)
);

BUFx10_ASAP7_75t_L g14291 ( 
.A(n_13146),
.Y(n_14291)
);

AOI22xp33_ASAP7_75t_SL g14292 ( 
.A1(n_13660),
.A2(n_12684),
.B1(n_12882),
.B2(n_10803),
.Y(n_14292)
);

AND2x2_ASAP7_75t_L g14293 ( 
.A(n_13334),
.B(n_11498),
.Y(n_14293)
);

AOI22xp5_ASAP7_75t_L g14294 ( 
.A1(n_13777),
.A2(n_11857),
.B1(n_12220),
.B2(n_12225),
.Y(n_14294)
);

INVx2_ASAP7_75t_L g14295 ( 
.A(n_13221),
.Y(n_14295)
);

NOR2xp33_ASAP7_75t_L g14296 ( 
.A(n_13061),
.B(n_10862),
.Y(n_14296)
);

NOR2xp33_ASAP7_75t_SL g14297 ( 
.A(n_13573),
.B(n_13354),
.Y(n_14297)
);

AO32x2_ASAP7_75t_L g14298 ( 
.A1(n_13832),
.A2(n_12168),
.A3(n_12350),
.B1(n_12334),
.B2(n_12314),
.Y(n_14298)
);

AND2x4_ASAP7_75t_L g14299 ( 
.A(n_13830),
.B(n_11498),
.Y(n_14299)
);

AOI22xp5_ASAP7_75t_L g14300 ( 
.A1(n_13660),
.A2(n_12183),
.B1(n_12184),
.B2(n_12159),
.Y(n_14300)
);

AND2x2_ASAP7_75t_L g14301 ( 
.A(n_13356),
.B(n_11498),
.Y(n_14301)
);

NAND2xp5_ASAP7_75t_L g14302 ( 
.A(n_13113),
.B(n_12889),
.Y(n_14302)
);

INVx6_ASAP7_75t_L g14303 ( 
.A(n_13784),
.Y(n_14303)
);

BUFx3_ASAP7_75t_L g14304 ( 
.A(n_12987),
.Y(n_14304)
);

OR2x2_ASAP7_75t_L g14305 ( 
.A(n_13739),
.B(n_11869),
.Y(n_14305)
);

INVx5_ASAP7_75t_SL g14306 ( 
.A(n_13221),
.Y(n_14306)
);

OA21x2_ASAP7_75t_L g14307 ( 
.A1(n_13962),
.A2(n_11807),
.B(n_11786),
.Y(n_14307)
);

NOR2xp33_ASAP7_75t_L g14308 ( 
.A(n_13095),
.B(n_10862),
.Y(n_14308)
);

INVx2_ASAP7_75t_SL g14309 ( 
.A(n_13870),
.Y(n_14309)
);

CKINVDCx5p33_ASAP7_75t_R g14310 ( 
.A(n_13293),
.Y(n_14310)
);

INVx3_ASAP7_75t_L g14311 ( 
.A(n_13221),
.Y(n_14311)
);

NAND2xp5_ASAP7_75t_L g14312 ( 
.A(n_13138),
.B(n_12896),
.Y(n_14312)
);

NOR2x1_ASAP7_75t_SL g14313 ( 
.A(n_13541),
.B(n_9968),
.Y(n_14313)
);

INVx1_ASAP7_75t_L g14314 ( 
.A(n_12996),
.Y(n_14314)
);

AND2x2_ASAP7_75t_L g14315 ( 
.A(n_13364),
.B(n_11532),
.Y(n_14315)
);

OAI21xp5_ASAP7_75t_L g14316 ( 
.A1(n_13801),
.A2(n_12208),
.B(n_12203),
.Y(n_14316)
);

AND2x4_ASAP7_75t_L g14317 ( 
.A(n_13870),
.B(n_11532),
.Y(n_14317)
);

NOR2x1_ASAP7_75t_SL g14318 ( 
.A(n_13541),
.B(n_9968),
.Y(n_14318)
);

OAI211xp5_ASAP7_75t_SL g14319 ( 
.A1(n_13801),
.A2(n_12369),
.B(n_12452),
.C(n_12383),
.Y(n_14319)
);

O2A1O1Ixp33_ASAP7_75t_L g14320 ( 
.A1(n_13586),
.A2(n_12865),
.B(n_12455),
.C(n_12475),
.Y(n_14320)
);

OR2x6_ASAP7_75t_L g14321 ( 
.A(n_13532),
.B(n_9968),
.Y(n_14321)
);

OAI22xp5_ASAP7_75t_L g14322 ( 
.A1(n_13238),
.A2(n_12882),
.B1(n_12684),
.B2(n_11083),
.Y(n_14322)
);

AND2x2_ASAP7_75t_L g14323 ( 
.A(n_13367),
.B(n_11532),
.Y(n_14323)
);

AO22x2_ASAP7_75t_L g14324 ( 
.A1(n_13054),
.A2(n_12521),
.B1(n_11680),
.B2(n_11684),
.Y(n_14324)
);

AOI221xp5_ASAP7_75t_L g14325 ( 
.A1(n_13889),
.A2(n_12873),
.B1(n_10441),
.B2(n_10475),
.C(n_10474),
.Y(n_14325)
);

AND2x4_ASAP7_75t_L g14326 ( 
.A(n_13071),
.B(n_11532),
.Y(n_14326)
);

OAI22xp5_ASAP7_75t_L g14327 ( 
.A1(n_13238),
.A2(n_11083),
.B1(n_11390),
.B2(n_10862),
.Y(n_14327)
);

AND2x4_ASAP7_75t_L g14328 ( 
.A(n_13074),
.B(n_11532),
.Y(n_14328)
);

AO21x2_ASAP7_75t_L g14329 ( 
.A1(n_12908),
.A2(n_11684),
.B(n_11668),
.Y(n_14329)
);

OR2x2_ASAP7_75t_L g14330 ( 
.A(n_13746),
.B(n_11878),
.Y(n_14330)
);

INVx2_ASAP7_75t_L g14331 ( 
.A(n_13117),
.Y(n_14331)
);

AND2x4_ASAP7_75t_L g14332 ( 
.A(n_13309),
.B(n_11539),
.Y(n_14332)
);

NOR2x1_ASAP7_75t_SL g14333 ( 
.A(n_13276),
.B(n_9968),
.Y(n_14333)
);

OAI21x1_ASAP7_75t_SL g14334 ( 
.A1(n_13260),
.A2(n_10778),
.B(n_12296),
.Y(n_14334)
);

INVx1_ASAP7_75t_L g14335 ( 
.A(n_13001),
.Y(n_14335)
);

AND2x4_ASAP7_75t_L g14336 ( 
.A(n_13470),
.B(n_11539),
.Y(n_14336)
);

INVx1_ASAP7_75t_L g14337 ( 
.A(n_13001),
.Y(n_14337)
);

OAI21x1_ASAP7_75t_SL g14338 ( 
.A1(n_13177),
.A2(n_10778),
.B(n_12296),
.Y(n_14338)
);

AND2x2_ASAP7_75t_L g14339 ( 
.A(n_13409),
.B(n_11539),
.Y(n_14339)
);

OAI22xp5_ASAP7_75t_L g14340 ( 
.A1(n_13382),
.A2(n_11083),
.B1(n_11390),
.B2(n_10862),
.Y(n_14340)
);

OAI21xp5_ASAP7_75t_L g14341 ( 
.A1(n_13889),
.A2(n_11994),
.B(n_12692),
.Y(n_14341)
);

OAI21xp5_ASAP7_75t_L g14342 ( 
.A1(n_13691),
.A2(n_12032),
.B(n_12017),
.Y(n_14342)
);

INVx1_ASAP7_75t_L g14343 ( 
.A(n_13008),
.Y(n_14343)
);

OAI22xp5_ASAP7_75t_L g14344 ( 
.A1(n_13382),
.A2(n_13651),
.B1(n_13288),
.B2(n_13137),
.Y(n_14344)
);

BUFx6f_ASAP7_75t_L g14345 ( 
.A(n_13532),
.Y(n_14345)
);

AND2x2_ASAP7_75t_L g14346 ( 
.A(n_13447),
.B(n_11539),
.Y(n_14346)
);

OR2x2_ASAP7_75t_L g14347 ( 
.A(n_13747),
.B(n_11701),
.Y(n_14347)
);

INVx1_ASAP7_75t_L g14348 ( 
.A(n_13008),
.Y(n_14348)
);

AND2x2_ASAP7_75t_L g14349 ( 
.A(n_13448),
.B(n_11539),
.Y(n_14349)
);

OAI21xp5_ASAP7_75t_L g14350 ( 
.A1(n_13691),
.A2(n_12062),
.B(n_12050),
.Y(n_14350)
);

A2O1A1Ixp33_ASAP7_75t_L g14351 ( 
.A1(n_13953),
.A2(n_12789),
.B(n_12467),
.C(n_12552),
.Y(n_14351)
);

AO32x2_ASAP7_75t_L g14352 ( 
.A1(n_13857),
.A2(n_12376),
.A3(n_12745),
.B1(n_12732),
.B2(n_12780),
.Y(n_14352)
);

AND2x2_ASAP7_75t_L g14353 ( 
.A(n_13451),
.B(n_11549),
.Y(n_14353)
);

NAND2xp5_ASAP7_75t_L g14354 ( 
.A(n_13142),
.B(n_12653),
.Y(n_14354)
);

AO21x1_ASAP7_75t_L g14355 ( 
.A1(n_13059),
.A2(n_12521),
.B(n_11807),
.Y(n_14355)
);

AOI221xp5_ASAP7_75t_L g14356 ( 
.A1(n_13537),
.A2(n_10474),
.B1(n_10481),
.B2(n_10475),
.C(n_10452),
.Y(n_14356)
);

NAND2xp33_ASAP7_75t_L g14357 ( 
.A(n_13538),
.B(n_9668),
.Y(n_14357)
);

AND2x2_ASAP7_75t_L g14358 ( 
.A(n_13102),
.B(n_11549),
.Y(n_14358)
);

OA21x2_ASAP7_75t_L g14359 ( 
.A1(n_13800),
.A2(n_11817),
.B(n_11786),
.Y(n_14359)
);

AND2x2_ASAP7_75t_L g14360 ( 
.A(n_13122),
.B(n_11549),
.Y(n_14360)
);

OR2x2_ASAP7_75t_L g14361 ( 
.A(n_13002),
.B(n_11725),
.Y(n_14361)
);

INVx1_ASAP7_75t_L g14362 ( 
.A(n_13153),
.Y(n_14362)
);

AND2x4_ASAP7_75t_L g14363 ( 
.A(n_13588),
.B(n_11549),
.Y(n_14363)
);

INVx1_ASAP7_75t_SL g14364 ( 
.A(n_13735),
.Y(n_14364)
);

OR2x2_ASAP7_75t_L g14365 ( 
.A(n_13009),
.B(n_11907),
.Y(n_14365)
);

CKINVDCx5p33_ASAP7_75t_R g14366 ( 
.A(n_13518),
.Y(n_14366)
);

AND2x2_ASAP7_75t_L g14367 ( 
.A(n_13124),
.B(n_11549),
.Y(n_14367)
);

OA21x2_ASAP7_75t_L g14368 ( 
.A1(n_13800),
.A2(n_11866),
.B(n_11817),
.Y(n_14368)
);

AND2x2_ASAP7_75t_L g14369 ( 
.A(n_12943),
.B(n_12960),
.Y(n_14369)
);

NAND2xp5_ASAP7_75t_SL g14370 ( 
.A(n_13385),
.B(n_12091),
.Y(n_14370)
);

AND2x2_ASAP7_75t_L g14371 ( 
.A(n_13384),
.B(n_11269),
.Y(n_14371)
);

OR2x2_ASAP7_75t_L g14372 ( 
.A(n_13011),
.B(n_11914),
.Y(n_14372)
);

INVx4_ASAP7_75t_L g14373 ( 
.A(n_13538),
.Y(n_14373)
);

HB1xp67_ASAP7_75t_L g14374 ( 
.A(n_13153),
.Y(n_14374)
);

AOI221x1_ASAP7_75t_L g14375 ( 
.A1(n_13385),
.A2(n_12820),
.B1(n_12881),
.B2(n_12804),
.C(n_12784),
.Y(n_14375)
);

OR2x2_ASAP7_75t_L g14376 ( 
.A(n_13894),
.B(n_11934),
.Y(n_14376)
);

AND2x2_ASAP7_75t_L g14377 ( 
.A(n_13384),
.B(n_11269),
.Y(n_14377)
);

OAI21xp5_ASAP7_75t_L g14378 ( 
.A1(n_13537),
.A2(n_12133),
.B(n_12132),
.Y(n_14378)
);

INVx1_ASAP7_75t_L g14379 ( 
.A(n_13154),
.Y(n_14379)
);

AO21x2_ASAP7_75t_L g14380 ( 
.A1(n_12908),
.A2(n_11694),
.B(n_11691),
.Y(n_14380)
);

NOR2x1_ASAP7_75t_SL g14381 ( 
.A(n_13276),
.B(n_9984),
.Y(n_14381)
);

OAI21xp5_ASAP7_75t_L g14382 ( 
.A1(n_13959),
.A2(n_12137),
.B(n_10281),
.Y(n_14382)
);

AO21x1_ASAP7_75t_L g14383 ( 
.A1(n_13059),
.A2(n_11897),
.B(n_11866),
.Y(n_14383)
);

AOI22xp5_ASAP7_75t_L g14384 ( 
.A1(n_13137),
.A2(n_11585),
.B1(n_11057),
.B2(n_11083),
.Y(n_14384)
);

OAI21xp5_ASAP7_75t_L g14385 ( 
.A1(n_13137),
.A2(n_10281),
.B(n_10700),
.Y(n_14385)
);

AO32x2_ASAP7_75t_L g14386 ( 
.A1(n_13857),
.A2(n_12890),
.A3(n_12264),
.B1(n_12241),
.B2(n_9781),
.Y(n_14386)
);

OAI211xp5_ASAP7_75t_SL g14387 ( 
.A1(n_13799),
.A2(n_12787),
.B(n_12788),
.C(n_12742),
.Y(n_14387)
);

AND2x4_ASAP7_75t_L g14388 ( 
.A(n_13611),
.B(n_10012),
.Y(n_14388)
);

OAI22xp5_ASAP7_75t_SL g14389 ( 
.A1(n_13288),
.A2(n_10086),
.B1(n_9984),
.B2(n_10862),
.Y(n_14389)
);

OA21x2_ASAP7_75t_L g14390 ( 
.A1(n_13809),
.A2(n_11902),
.B(n_11897),
.Y(n_14390)
);

AND2x4_ASAP7_75t_L g14391 ( 
.A(n_13617),
.B(n_13556),
.Y(n_14391)
);

OAI21xp5_ASAP7_75t_L g14392 ( 
.A1(n_13288),
.A2(n_10712),
.B(n_10700),
.Y(n_14392)
);

AOI22xp33_ASAP7_75t_SL g14393 ( 
.A1(n_13888),
.A2(n_10803),
.B1(n_9838),
.B2(n_9892),
.Y(n_14393)
);

NAND2xp5_ASAP7_75t_L g14394 ( 
.A(n_13147),
.B(n_12796),
.Y(n_14394)
);

INVx1_ASAP7_75t_L g14395 ( 
.A(n_13154),
.Y(n_14395)
);

OA21x2_ASAP7_75t_L g14396 ( 
.A1(n_13809),
.A2(n_11913),
.B(n_11902),
.Y(n_14396)
);

NAND3xp33_ASAP7_75t_L g14397 ( 
.A(n_13802),
.B(n_10803),
.C(n_11464),
.Y(n_14397)
);

AND2x4_ASAP7_75t_L g14398 ( 
.A(n_13571),
.B(n_10012),
.Y(n_14398)
);

OAI21xp5_ASAP7_75t_L g14399 ( 
.A1(n_13642),
.A2(n_10712),
.B(n_10700),
.Y(n_14399)
);

HB1xp67_ASAP7_75t_L g14400 ( 
.A(n_13553),
.Y(n_14400)
);

INVx2_ASAP7_75t_SL g14401 ( 
.A(n_13538),
.Y(n_14401)
);

INVx4_ASAP7_75t_L g14402 ( 
.A(n_13784),
.Y(n_14402)
);

AND2x2_ASAP7_75t_L g14403 ( 
.A(n_13390),
.B(n_11269),
.Y(n_14403)
);

NOR2x1_ASAP7_75t_SL g14404 ( 
.A(n_13123),
.B(n_9984),
.Y(n_14404)
);

NOR2xp33_ASAP7_75t_L g14405 ( 
.A(n_13095),
.B(n_11083),
.Y(n_14405)
);

INVx1_ASAP7_75t_L g14406 ( 
.A(n_13054),
.Y(n_14406)
);

INVx3_ASAP7_75t_L g14407 ( 
.A(n_13845),
.Y(n_14407)
);

INVx1_ASAP7_75t_L g14408 ( 
.A(n_13051),
.Y(n_14408)
);

AND2x2_ASAP7_75t_L g14409 ( 
.A(n_13390),
.B(n_11269),
.Y(n_14409)
);

AND2x4_ASAP7_75t_L g14410 ( 
.A(n_13608),
.B(n_10049),
.Y(n_14410)
);

INVx2_ASAP7_75t_L g14411 ( 
.A(n_13350),
.Y(n_14411)
);

AND2x2_ASAP7_75t_L g14412 ( 
.A(n_13729),
.B(n_11269),
.Y(n_14412)
);

NOR2xp33_ASAP7_75t_L g14413 ( 
.A(n_12978),
.B(n_11083),
.Y(n_14413)
);

AND2x4_ASAP7_75t_L g14414 ( 
.A(n_13609),
.B(n_10049),
.Y(n_14414)
);

OAI211xp5_ASAP7_75t_L g14415 ( 
.A1(n_13797),
.A2(n_10481),
.B(n_10631),
.C(n_10612),
.Y(n_14415)
);

INVx1_ASAP7_75t_L g14416 ( 
.A(n_13052),
.Y(n_14416)
);

NOR2x1_ASAP7_75t_L g14417 ( 
.A(n_13934),
.B(n_13053),
.Y(n_14417)
);

NAND2x1_ASAP7_75t_L g14418 ( 
.A(n_13616),
.B(n_13581),
.Y(n_14418)
);

AOI211xp5_ASAP7_75t_L g14419 ( 
.A1(n_13671),
.A2(n_11465),
.B(n_11464),
.C(n_10631),
.Y(n_14419)
);

HB1xp67_ASAP7_75t_L g14420 ( 
.A(n_13553),
.Y(n_14420)
);

NAND3xp33_ASAP7_75t_L g14421 ( 
.A(n_13859),
.B(n_10803),
.C(n_11465),
.Y(n_14421)
);

INVx2_ASAP7_75t_L g14422 ( 
.A(n_13350),
.Y(n_14422)
);

AND2x2_ASAP7_75t_L g14423 ( 
.A(n_13740),
.B(n_13378),
.Y(n_14423)
);

NOR2x1_ASAP7_75t_L g14424 ( 
.A(n_13934),
.B(n_12296),
.Y(n_14424)
);

NOR2xp33_ASAP7_75t_L g14425 ( 
.A(n_12978),
.B(n_11390),
.Y(n_14425)
);

NAND2xp5_ASAP7_75t_L g14426 ( 
.A(n_13637),
.B(n_12807),
.Y(n_14426)
);

OR2x2_ASAP7_75t_L g14427 ( 
.A(n_13894),
.B(n_11965),
.Y(n_14427)
);

AOI221xp5_ASAP7_75t_L g14428 ( 
.A1(n_13639),
.A2(n_10641),
.B1(n_10784),
.B2(n_10661),
.C(n_10612),
.Y(n_14428)
);

AOI221xp5_ASAP7_75t_L g14429 ( 
.A1(n_13643),
.A2(n_13657),
.B1(n_13656),
.B2(n_13648),
.C(n_13799),
.Y(n_14429)
);

AND2x4_ASAP7_75t_L g14430 ( 
.A(n_13664),
.B(n_10049),
.Y(n_14430)
);

INVx11_ASAP7_75t_L g14431 ( 
.A(n_13023),
.Y(n_14431)
);

AND2x4_ASAP7_75t_L g14432 ( 
.A(n_13718),
.B(n_10049),
.Y(n_14432)
);

AND2x4_ASAP7_75t_L g14433 ( 
.A(n_13023),
.B(n_10049),
.Y(n_14433)
);

AO32x2_ASAP7_75t_L g14434 ( 
.A1(n_13804),
.A2(n_9781),
.A3(n_9851),
.B1(n_9759),
.B2(n_9706),
.Y(n_14434)
);

OR2x2_ASAP7_75t_L g14435 ( 
.A(n_13699),
.B(n_11984),
.Y(n_14435)
);

NOR2xp33_ASAP7_75t_L g14436 ( 
.A(n_13024),
.B(n_11390),
.Y(n_14436)
);

AND2x2_ASAP7_75t_L g14437 ( 
.A(n_13031),
.B(n_11275),
.Y(n_14437)
);

INVx2_ASAP7_75t_L g14438 ( 
.A(n_13366),
.Y(n_14438)
);

NOR2xp33_ASAP7_75t_L g14439 ( 
.A(n_13024),
.B(n_13735),
.Y(n_14439)
);

INVx2_ASAP7_75t_L g14440 ( 
.A(n_13366),
.Y(n_14440)
);

O2A1O1Ixp33_ASAP7_75t_SL g14441 ( 
.A1(n_13259),
.A2(n_11383),
.B(n_11926),
.C(n_11913),
.Y(n_14441)
);

OR2x2_ASAP7_75t_L g14442 ( 
.A(n_13700),
.B(n_11998),
.Y(n_14442)
);

AND2x2_ASAP7_75t_L g14443 ( 
.A(n_13042),
.B(n_11275),
.Y(n_14443)
);

AO21x2_ASAP7_75t_L g14444 ( 
.A1(n_13811),
.A2(n_11694),
.B(n_11691),
.Y(n_14444)
);

OAI21xp5_ASAP7_75t_L g14445 ( 
.A1(n_13642),
.A2(n_10723),
.B(n_10712),
.Y(n_14445)
);

NOR2x1_ASAP7_75t_L g14446 ( 
.A(n_13053),
.B(n_12838),
.Y(n_14446)
);

NAND2xp5_ASAP7_75t_L g14447 ( 
.A(n_13942),
.B(n_12878),
.Y(n_14447)
);

INVx3_ASAP7_75t_L g14448 ( 
.A(n_13845),
.Y(n_14448)
);

O2A1O1Ixp33_ASAP7_75t_L g14449 ( 
.A1(n_13642),
.A2(n_10641),
.B(n_10784),
.C(n_10661),
.Y(n_14449)
);

AO21x2_ASAP7_75t_L g14450 ( 
.A1(n_13811),
.A2(n_11715),
.B(n_11926),
.Y(n_14450)
);

OAI21xp5_ASAP7_75t_L g14451 ( 
.A1(n_13244),
.A2(n_13250),
.B(n_13130),
.Y(n_14451)
);

AO21x1_ASAP7_75t_L g14452 ( 
.A1(n_13404),
.A2(n_11960),
.B(n_11715),
.Y(n_14452)
);

AOI221xp5_ASAP7_75t_L g14453 ( 
.A1(n_13055),
.A2(n_11080),
.B1(n_11239),
.B2(n_11210),
.C(n_11065),
.Y(n_14453)
);

O2A1O1Ixp33_ASAP7_75t_SL g14454 ( 
.A1(n_13294),
.A2(n_11383),
.B(n_11960),
.C(n_12265),
.Y(n_14454)
);

OR2x2_ASAP7_75t_L g14455 ( 
.A(n_13072),
.B(n_12580),
.Y(n_14455)
);

BUFx3_ASAP7_75t_L g14456 ( 
.A(n_13919),
.Y(n_14456)
);

OR2x6_ASAP7_75t_L g14457 ( 
.A(n_13804),
.B(n_9984),
.Y(n_14457)
);

OAI211xp5_ASAP7_75t_SL g14458 ( 
.A1(n_13819),
.A2(n_12613),
.B(n_12645),
.C(n_12610),
.Y(n_14458)
);

AND2x4_ASAP7_75t_L g14459 ( 
.A(n_13930),
.B(n_10106),
.Y(n_14459)
);

AOI22xp5_ASAP7_75t_L g14460 ( 
.A1(n_12923),
.A2(n_11585),
.B1(n_11057),
.B2(n_11390),
.Y(n_14460)
);

NOR2xp33_ASAP7_75t_L g14461 ( 
.A(n_13671),
.B(n_11390),
.Y(n_14461)
);

INVx1_ASAP7_75t_L g14462 ( 
.A(n_13058),
.Y(n_14462)
);

AND2x2_ASAP7_75t_L g14463 ( 
.A(n_13070),
.B(n_11275),
.Y(n_14463)
);

OA21x2_ASAP7_75t_L g14464 ( 
.A1(n_13404),
.A2(n_12330),
.B(n_12265),
.Y(n_14464)
);

AO32x2_ASAP7_75t_L g14465 ( 
.A1(n_13750),
.A2(n_9851),
.A3(n_9860),
.B1(n_9781),
.B2(n_9759),
.Y(n_14465)
);

NOR2x1_ASAP7_75t_SL g14466 ( 
.A(n_13123),
.B(n_9984),
.Y(n_14466)
);

AO32x2_ASAP7_75t_L g14467 ( 
.A1(n_13750),
.A2(n_9851),
.A3(n_9860),
.B1(n_9781),
.B2(n_9759),
.Y(n_14467)
);

AND2x2_ASAP7_75t_L g14468 ( 
.A(n_13080),
.B(n_11275),
.Y(n_14468)
);

AND2x2_ASAP7_75t_L g14469 ( 
.A(n_13082),
.B(n_11275),
.Y(n_14469)
);

AOI21xp5_ASAP7_75t_L g14470 ( 
.A1(n_13053),
.A2(n_10773),
.B(n_10746),
.Y(n_14470)
);

AND2x2_ASAP7_75t_L g14471 ( 
.A(n_12979),
.B(n_11320),
.Y(n_14471)
);

INVx1_ASAP7_75t_L g14472 ( 
.A(n_13064),
.Y(n_14472)
);

HB1xp67_ASAP7_75t_L g14473 ( 
.A(n_13602),
.Y(n_14473)
);

AND2x2_ASAP7_75t_L g14474 ( 
.A(n_13696),
.B(n_11320),
.Y(n_14474)
);

OAI21x1_ASAP7_75t_SL g14475 ( 
.A1(n_13589),
.A2(n_13805),
.B(n_13511),
.Y(n_14475)
);

AOI221xp5_ASAP7_75t_L g14476 ( 
.A1(n_13066),
.A2(n_11210),
.B1(n_11239),
.B2(n_11080),
.C(n_11065),
.Y(n_14476)
);

HB1xp67_ASAP7_75t_L g14477 ( 
.A(n_13602),
.Y(n_14477)
);

OR2x2_ASAP7_75t_L g14478 ( 
.A(n_13078),
.B(n_12597),
.Y(n_14478)
);

NOR2x1_ASAP7_75t_SL g14479 ( 
.A(n_13172),
.B(n_10086),
.Y(n_14479)
);

AOI221xp5_ASAP7_75t_L g14480 ( 
.A1(n_13073),
.A2(n_11392),
.B1(n_11421),
.B2(n_11370),
.C(n_11314),
.Y(n_14480)
);

AOI21xp5_ASAP7_75t_SL g14481 ( 
.A1(n_12986),
.A2(n_13041),
.B(n_12995),
.Y(n_14481)
);

OAI21xp5_ASAP7_75t_L g14482 ( 
.A1(n_13130),
.A2(n_10731),
.B(n_10723),
.Y(n_14482)
);

BUFx6f_ASAP7_75t_L g14483 ( 
.A(n_13919),
.Y(n_14483)
);

OR2x6_ASAP7_75t_L g14484 ( 
.A(n_13919),
.B(n_10086),
.Y(n_14484)
);

AND2x2_ASAP7_75t_L g14485 ( 
.A(n_13843),
.B(n_13940),
.Y(n_14485)
);

OR2x2_ASAP7_75t_L g14486 ( 
.A(n_13081),
.B(n_12652),
.Y(n_14486)
);

OR2x2_ASAP7_75t_L g14487 ( 
.A(n_13085),
.B(n_12261),
.Y(n_14487)
);

INVx1_ASAP7_75t_L g14488 ( 
.A(n_13084),
.Y(n_14488)
);

A2O1A1Ixp33_ASAP7_75t_L g14489 ( 
.A1(n_13094),
.A2(n_13457),
.B(n_13525),
.C(n_13450),
.Y(n_14489)
);

AND2x2_ASAP7_75t_L g14490 ( 
.A(n_13943),
.B(n_11320),
.Y(n_14490)
);

AND2x2_ASAP7_75t_L g14491 ( 
.A(n_13128),
.B(n_11320),
.Y(n_14491)
);

AND2x4_ASAP7_75t_SL g14492 ( 
.A(n_13754),
.B(n_13823),
.Y(n_14492)
);

OAI21xp5_ASAP7_75t_L g14493 ( 
.A1(n_13005),
.A2(n_13842),
.B(n_13339),
.Y(n_14493)
);

INVx2_ASAP7_75t_L g14494 ( 
.A(n_13377),
.Y(n_14494)
);

NOR2x1_ASAP7_75t_SL g14495 ( 
.A(n_13172),
.B(n_10086),
.Y(n_14495)
);

NOR2xp33_ASAP7_75t_L g14496 ( 
.A(n_13754),
.B(n_10086),
.Y(n_14496)
);

OR2x2_ASAP7_75t_L g14497 ( 
.A(n_13661),
.B(n_12283),
.Y(n_14497)
);

AND2x2_ASAP7_75t_L g14498 ( 
.A(n_13132),
.B(n_11320),
.Y(n_14498)
);

AND2x2_ASAP7_75t_L g14499 ( 
.A(n_13136),
.B(n_13164),
.Y(n_14499)
);

INVxp33_ASAP7_75t_L g14500 ( 
.A(n_13503),
.Y(n_14500)
);

NAND2xp5_ASAP7_75t_L g14501 ( 
.A(n_13822),
.B(n_12696),
.Y(n_14501)
);

BUFx8_ASAP7_75t_SL g14502 ( 
.A(n_13947),
.Y(n_14502)
);

INVx1_ASAP7_75t_L g14503 ( 
.A(n_13086),
.Y(n_14503)
);

OAI22xp5_ASAP7_75t_SL g14504 ( 
.A1(n_12928),
.A2(n_10583),
.B1(n_9167),
.B2(n_9169),
.Y(n_14504)
);

OA21x2_ASAP7_75t_L g14505 ( 
.A1(n_13763),
.A2(n_13780),
.B(n_13764),
.Y(n_14505)
);

O2A1O1Ixp33_ASAP7_75t_SL g14506 ( 
.A1(n_13483),
.A2(n_11383),
.B(n_12352),
.C(n_12330),
.Y(n_14506)
);

OAI21x1_ASAP7_75t_SL g14507 ( 
.A1(n_13420),
.A2(n_9662),
.B(n_11660),
.Y(n_14507)
);

AOI21xp33_ASAP7_75t_SL g14508 ( 
.A1(n_12928),
.A2(n_13510),
.B(n_13503),
.Y(n_14508)
);

INVx1_ASAP7_75t_L g14509 ( 
.A(n_13098),
.Y(n_14509)
);

A2O1A1Ixp33_ASAP7_75t_L g14510 ( 
.A1(n_13527),
.A2(n_11370),
.B(n_11392),
.C(n_11314),
.Y(n_14510)
);

AND2x4_ASAP7_75t_L g14511 ( 
.A(n_13930),
.B(n_10106),
.Y(n_14511)
);

AND2x2_ASAP7_75t_L g14512 ( 
.A(n_13183),
.B(n_10199),
.Y(n_14512)
);

AO21x2_ASAP7_75t_L g14513 ( 
.A1(n_13036),
.A2(n_12364),
.B(n_12352),
.Y(n_14513)
);

INVx2_ASAP7_75t_SL g14514 ( 
.A(n_13377),
.Y(n_14514)
);

AOI21xp5_ASAP7_75t_L g14515 ( 
.A1(n_12928),
.A2(n_10773),
.B(n_10707),
.Y(n_14515)
);

AND2x4_ASAP7_75t_L g14516 ( 
.A(n_13930),
.B(n_10106),
.Y(n_14516)
);

NOR2x1_ASAP7_75t_SL g14517 ( 
.A(n_12993),
.B(n_9004),
.Y(n_14517)
);

AND2x2_ASAP7_75t_L g14518 ( 
.A(n_13191),
.B(n_10199),
.Y(n_14518)
);

AND2x6_ASAP7_75t_L g14519 ( 
.A(n_13947),
.B(n_10435),
.Y(n_14519)
);

AOI21xp5_ASAP7_75t_L g14520 ( 
.A1(n_13646),
.A2(n_10773),
.B(n_10707),
.Y(n_14520)
);

OAI21xp5_ASAP7_75t_L g14521 ( 
.A1(n_13938),
.A2(n_10731),
.B(n_10723),
.Y(n_14521)
);

OAI21xp5_ASAP7_75t_L g14522 ( 
.A1(n_13647),
.A2(n_10733),
.B(n_10731),
.Y(n_14522)
);

AND2x2_ASAP7_75t_L g14523 ( 
.A(n_13193),
.B(n_10199),
.Y(n_14523)
);

AOI22xp5_ASAP7_75t_L g14524 ( 
.A1(n_13228),
.A2(n_11585),
.B1(n_11057),
.B2(n_10424),
.Y(n_14524)
);

BUFx2_ASAP7_75t_L g14525 ( 
.A(n_13003),
.Y(n_14525)
);

INVx1_ASAP7_75t_L g14526 ( 
.A(n_13103),
.Y(n_14526)
);

INVx2_ASAP7_75t_L g14527 ( 
.A(n_13529),
.Y(n_14527)
);

NOR2x1_ASAP7_75t_SL g14528 ( 
.A(n_12993),
.B(n_9004),
.Y(n_14528)
);

AO32x2_ASAP7_75t_L g14529 ( 
.A1(n_13750),
.A2(n_9851),
.A3(n_9860),
.B1(n_9781),
.B2(n_9759),
.Y(n_14529)
);

NOR2xp33_ASAP7_75t_L g14530 ( 
.A(n_13823),
.B(n_13510),
.Y(n_14530)
);

NAND2xp5_ASAP7_75t_L g14531 ( 
.A(n_13828),
.B(n_12703),
.Y(n_14531)
);

BUFx6f_ASAP7_75t_L g14532 ( 
.A(n_13947),
.Y(n_14532)
);

AND2x4_ASAP7_75t_L g14533 ( 
.A(n_13784),
.B(n_10106),
.Y(n_14533)
);

AND2x2_ASAP7_75t_L g14534 ( 
.A(n_13200),
.B(n_10199),
.Y(n_14534)
);

A2O1A1Ixp33_ASAP7_75t_L g14535 ( 
.A1(n_13540),
.A2(n_11527),
.B(n_11543),
.C(n_11421),
.Y(n_14535)
);

AND2x2_ASAP7_75t_L g14536 ( 
.A(n_13215),
.B(n_10199),
.Y(n_14536)
);

OAI22xp5_ASAP7_75t_L g14537 ( 
.A1(n_12974),
.A2(n_13049),
.B1(n_13029),
.B2(n_13565),
.Y(n_14537)
);

A2O1A1Ixp33_ASAP7_75t_L g14538 ( 
.A1(n_13737),
.A2(n_11543),
.B(n_11566),
.C(n_11527),
.Y(n_14538)
);

AO32x2_ASAP7_75t_L g14539 ( 
.A1(n_12961),
.A2(n_9860),
.A3(n_9891),
.B1(n_9851),
.B2(n_9759),
.Y(n_14539)
);

OAI21xp5_ASAP7_75t_L g14540 ( 
.A1(n_13745),
.A2(n_10733),
.B(n_10651),
.Y(n_14540)
);

NOR2x1_ASAP7_75t_SL g14541 ( 
.A(n_13278),
.B(n_9004),
.Y(n_14541)
);

INVx1_ASAP7_75t_L g14542 ( 
.A(n_13106),
.Y(n_14542)
);

AND2x2_ASAP7_75t_L g14543 ( 
.A(n_13223),
.B(n_10223),
.Y(n_14543)
);

NOR2x1_ASAP7_75t_SL g14544 ( 
.A(n_13278),
.B(n_9004),
.Y(n_14544)
);

INVx1_ASAP7_75t_L g14545 ( 
.A(n_13107),
.Y(n_14545)
);

OAI22xp5_ASAP7_75t_SL g14546 ( 
.A1(n_13677),
.A2(n_10583),
.B1(n_9167),
.B2(n_9169),
.Y(n_14546)
);

INVx1_ASAP7_75t_L g14547 ( 
.A(n_13111),
.Y(n_14547)
);

INVx4_ASAP7_75t_L g14548 ( 
.A(n_13476),
.Y(n_14548)
);

INVx1_ASAP7_75t_L g14549 ( 
.A(n_13114),
.Y(n_14549)
);

AND2x2_ASAP7_75t_L g14550 ( 
.A(n_13265),
.B(n_10223),
.Y(n_14550)
);

O2A1O1Ixp33_ASAP7_75t_L g14551 ( 
.A1(n_13625),
.A2(n_11590),
.B(n_11612),
.C(n_11566),
.Y(n_14551)
);

AND2x2_ASAP7_75t_L g14552 ( 
.A(n_13271),
.B(n_10223),
.Y(n_14552)
);

AND2x2_ASAP7_75t_L g14553 ( 
.A(n_13494),
.B(n_10223),
.Y(n_14553)
);

NAND2xp33_ASAP7_75t_L g14554 ( 
.A(n_13775),
.B(n_9965),
.Y(n_14554)
);

CKINVDCx5p33_ASAP7_75t_R g14555 ( 
.A(n_13677),
.Y(n_14555)
);

AOI22xp5_ASAP7_75t_L g14556 ( 
.A1(n_13228),
.A2(n_11585),
.B1(n_11057),
.B2(n_10424),
.Y(n_14556)
);

HB1xp67_ASAP7_75t_L g14557 ( 
.A(n_13625),
.Y(n_14557)
);

AND2x2_ASAP7_75t_L g14558 ( 
.A(n_13499),
.B(n_10223),
.Y(n_14558)
);

INVx1_ASAP7_75t_L g14559 ( 
.A(n_13119),
.Y(n_14559)
);

AND2x2_ASAP7_75t_L g14560 ( 
.A(n_13508),
.B(n_10232),
.Y(n_14560)
);

AND2x2_ASAP7_75t_L g14561 ( 
.A(n_13524),
.B(n_10232),
.Y(n_14561)
);

AOI21xp5_ASAP7_75t_L g14562 ( 
.A1(n_13646),
.A2(n_10707),
.B(n_10657),
.Y(n_14562)
);

AND2x2_ASAP7_75t_L g14563 ( 
.A(n_13533),
.B(n_10232),
.Y(n_14563)
);

HB1xp67_ASAP7_75t_L g14564 ( 
.A(n_13627),
.Y(n_14564)
);

AO32x2_ASAP7_75t_L g14565 ( 
.A1(n_13860),
.A2(n_9956),
.A3(n_9891),
.B1(n_9860),
.B2(n_12517),
.Y(n_14565)
);

INVx1_ASAP7_75t_L g14566 ( 
.A(n_13125),
.Y(n_14566)
);

OR2x2_ASAP7_75t_L g14567 ( 
.A(n_13662),
.B(n_12232),
.Y(n_14567)
);

NOR2xp33_ASAP7_75t_SL g14568 ( 
.A(n_13546),
.B(n_10625),
.Y(n_14568)
);

OA21x2_ASAP7_75t_L g14569 ( 
.A1(n_13763),
.A2(n_12375),
.B(n_12364),
.Y(n_14569)
);

AND2x2_ASAP7_75t_L g14570 ( 
.A(n_13967),
.B(n_13545),
.Y(n_14570)
);

INVx2_ASAP7_75t_L g14571 ( 
.A(n_13529),
.Y(n_14571)
);

AND2x2_ASAP7_75t_L g14572 ( 
.A(n_13557),
.B(n_10232),
.Y(n_14572)
);

CKINVDCx5p33_ASAP7_75t_R g14573 ( 
.A(n_13677),
.Y(n_14573)
);

NAND2xp5_ASAP7_75t_L g14574 ( 
.A(n_13835),
.B(n_12717),
.Y(n_14574)
);

AND2x2_ASAP7_75t_L g14575 ( 
.A(n_13575),
.B(n_10232),
.Y(n_14575)
);

INVx2_ASAP7_75t_L g14576 ( 
.A(n_13551),
.Y(n_14576)
);

A2O1A1Ixp33_ASAP7_75t_L g14577 ( 
.A1(n_13748),
.A2(n_11612),
.B(n_11590),
.C(n_9167),
.Y(n_14577)
);

AND2x2_ASAP7_75t_L g14578 ( 
.A(n_13618),
.B(n_10370),
.Y(n_14578)
);

OAI21xp5_ASAP7_75t_L g14579 ( 
.A1(n_13720),
.A2(n_10733),
.B(n_10651),
.Y(n_14579)
);

INVx3_ASAP7_75t_L g14580 ( 
.A(n_13752),
.Y(n_14580)
);

AOI22xp5_ASAP7_75t_L g14581 ( 
.A1(n_13516),
.A2(n_13542),
.B1(n_13974),
.B2(n_13467),
.Y(n_14581)
);

AND2x4_ASAP7_75t_L g14582 ( 
.A(n_12980),
.B(n_10106),
.Y(n_14582)
);

A2O1A1Ixp33_ASAP7_75t_L g14583 ( 
.A1(n_13579),
.A2(n_9167),
.B(n_9169),
.C(n_9158),
.Y(n_14583)
);

OR2x2_ASAP7_75t_L g14584 ( 
.A(n_13666),
.B(n_11594),
.Y(n_14584)
);

NAND2xp5_ASAP7_75t_L g14585 ( 
.A(n_13846),
.B(n_12721),
.Y(n_14585)
);

OR2x2_ASAP7_75t_L g14586 ( 
.A(n_13668),
.B(n_11594),
.Y(n_14586)
);

OR2x6_ASAP7_75t_L g14587 ( 
.A(n_13685),
.B(n_10178),
.Y(n_14587)
);

AND2x2_ASAP7_75t_L g14588 ( 
.A(n_13618),
.B(n_10370),
.Y(n_14588)
);

OAI22xp5_ASAP7_75t_L g14589 ( 
.A1(n_12974),
.A2(n_10583),
.B1(n_9443),
.B2(n_9167),
.Y(n_14589)
);

AND2x4_ASAP7_75t_L g14590 ( 
.A(n_12980),
.B(n_10106),
.Y(n_14590)
);

OR2x6_ASAP7_75t_L g14591 ( 
.A(n_13685),
.B(n_10178),
.Y(n_14591)
);

AND2x4_ASAP7_75t_L g14592 ( 
.A(n_13852),
.B(n_10106),
.Y(n_14592)
);

AND2x4_ASAP7_75t_L g14593 ( 
.A(n_13853),
.B(n_13854),
.Y(n_14593)
);

INVx2_ASAP7_75t_L g14594 ( 
.A(n_13551),
.Y(n_14594)
);

OAI22xp5_ASAP7_75t_L g14595 ( 
.A1(n_13029),
.A2(n_9167),
.B1(n_9169),
.B2(n_9158),
.Y(n_14595)
);

O2A1O1Ixp33_ASAP7_75t_L g14596 ( 
.A1(n_13627),
.A2(n_10651),
.B(n_10688),
.C(n_10568),
.Y(n_14596)
);

OA21x2_ASAP7_75t_L g14597 ( 
.A1(n_13780),
.A2(n_12527),
.B(n_12375),
.Y(n_14597)
);

OAI21xp5_ASAP7_75t_L g14598 ( 
.A1(n_13867),
.A2(n_10651),
.B(n_10568),
.Y(n_14598)
);

INVx11_ASAP7_75t_L g14599 ( 
.A(n_13685),
.Y(n_14599)
);

OAI22xp5_ASAP7_75t_L g14600 ( 
.A1(n_13049),
.A2(n_9169),
.B1(n_9204),
.B2(n_9158),
.Y(n_14600)
);

A2O1A1Ixp33_ASAP7_75t_L g14601 ( 
.A1(n_13028),
.A2(n_9169),
.B(n_9204),
.C(n_9158),
.Y(n_14601)
);

NAND2xp5_ASAP7_75t_L g14602 ( 
.A(n_13858),
.B(n_12727),
.Y(n_14602)
);

OAI21xp5_ASAP7_75t_L g14603 ( 
.A1(n_13873),
.A2(n_10688),
.B(n_10568),
.Y(n_14603)
);

AOI21xp5_ASAP7_75t_L g14604 ( 
.A1(n_13888),
.A2(n_13328),
.B(n_13555),
.Y(n_14604)
);

HB1xp67_ASAP7_75t_L g14605 ( 
.A(n_13126),
.Y(n_14605)
);

AND2x2_ASAP7_75t_L g14606 ( 
.A(n_13630),
.B(n_10370),
.Y(n_14606)
);

INVx3_ASAP7_75t_L g14607 ( 
.A(n_13752),
.Y(n_14607)
);

AND2x2_ASAP7_75t_L g14608 ( 
.A(n_13630),
.B(n_10370),
.Y(n_14608)
);

AND2x2_ASAP7_75t_L g14609 ( 
.A(n_13652),
.B(n_10370),
.Y(n_14609)
);

A2O1A1Ixp33_ASAP7_75t_L g14610 ( 
.A1(n_13665),
.A2(n_9204),
.B(n_9237),
.C(n_9158),
.Y(n_14610)
);

AND2x2_ASAP7_75t_L g14611 ( 
.A(n_13652),
.B(n_12728),
.Y(n_14611)
);

INVx2_ASAP7_75t_SL g14612 ( 
.A(n_13775),
.Y(n_14612)
);

O2A1O1Ixp33_ASAP7_75t_SL g14613 ( 
.A1(n_13487),
.A2(n_12538),
.B(n_12539),
.C(n_12527),
.Y(n_14613)
);

OAI22xp5_ASAP7_75t_L g14614 ( 
.A1(n_13782),
.A2(n_9204),
.B1(n_9237),
.B2(n_9158),
.Y(n_14614)
);

O2A1O1Ixp33_ASAP7_75t_SL g14615 ( 
.A1(n_13487),
.A2(n_12539),
.B(n_12538),
.C(n_11033),
.Y(n_14615)
);

NAND2xp5_ASAP7_75t_L g14616 ( 
.A(n_13861),
.B(n_12738),
.Y(n_14616)
);

BUFx12f_ASAP7_75t_L g14617 ( 
.A(n_12986),
.Y(n_14617)
);

AND2x2_ASAP7_75t_L g14618 ( 
.A(n_13676),
.B(n_13701),
.Y(n_14618)
);

AOI22xp5_ASAP7_75t_L g14619 ( 
.A1(n_13516),
.A2(n_13542),
.B1(n_13467),
.B2(n_13460),
.Y(n_14619)
);

OA21x2_ASAP7_75t_L g14620 ( 
.A1(n_13036),
.A2(n_12613),
.B(n_12610),
.Y(n_14620)
);

AO32x2_ASAP7_75t_L g14621 ( 
.A1(n_13860),
.A2(n_9956),
.A3(n_9891),
.B1(n_9349),
.B2(n_8568),
.Y(n_14621)
);

O2A1O1Ixp33_ASAP7_75t_SL g14622 ( 
.A1(n_13495),
.A2(n_11033),
.B(n_11215),
.C(n_11066),
.Y(n_14622)
);

AOI221xp5_ASAP7_75t_L g14623 ( 
.A1(n_13131),
.A2(n_11057),
.B1(n_11585),
.B2(n_11579),
.C(n_11569),
.Y(n_14623)
);

NOR2xp33_ASAP7_75t_L g14624 ( 
.A(n_12995),
.B(n_10625),
.Y(n_14624)
);

AOI211xp5_ASAP7_75t_L g14625 ( 
.A1(n_13041),
.A2(n_10670),
.B(n_10753),
.C(n_10711),
.Y(n_14625)
);

AND2x4_ASAP7_75t_L g14626 ( 
.A(n_13868),
.B(n_11577),
.Y(n_14626)
);

AOI22xp5_ASAP7_75t_L g14627 ( 
.A1(n_13460),
.A2(n_10424),
.B1(n_11137),
.B2(n_11118),
.Y(n_14627)
);

INVx2_ASAP7_75t_L g14628 ( 
.A(n_13574),
.Y(n_14628)
);

AND2x4_ASAP7_75t_SL g14629 ( 
.A(n_13770),
.B(n_13813),
.Y(n_14629)
);

AND2x4_ASAP7_75t_L g14630 ( 
.A(n_13871),
.B(n_13089),
.Y(n_14630)
);

O2A1O1Ixp33_ASAP7_75t_L g14631 ( 
.A1(n_13135),
.A2(n_10688),
.B(n_10568),
.C(n_12645),
.Y(n_14631)
);

AND2x2_ASAP7_75t_L g14632 ( 
.A(n_13676),
.B(n_13701),
.Y(n_14632)
);

OR2x2_ASAP7_75t_L g14633 ( 
.A(n_13669),
.B(n_13670),
.Y(n_14633)
);

AND2x4_ASAP7_75t_L g14634 ( 
.A(n_13089),
.B(n_11577),
.Y(n_14634)
);

AOI21xp5_ASAP7_75t_L g14635 ( 
.A1(n_13328),
.A2(n_10707),
.B(n_10657),
.Y(n_14635)
);

INVx1_ASAP7_75t_L g14636 ( 
.A(n_13139),
.Y(n_14636)
);

INVx1_ASAP7_75t_L g14637 ( 
.A(n_13143),
.Y(n_14637)
);

BUFx2_ASAP7_75t_L g14638 ( 
.A(n_13003),
.Y(n_14638)
);

AND2x2_ASAP7_75t_L g14639 ( 
.A(n_13708),
.B(n_12739),
.Y(n_14639)
);

NOR2xp33_ASAP7_75t_L g14640 ( 
.A(n_13770),
.B(n_10625),
.Y(n_14640)
);

OR2x6_ASAP7_75t_L g14641 ( 
.A(n_13770),
.B(n_10178),
.Y(n_14641)
);

CKINVDCx5p33_ASAP7_75t_R g14642 ( 
.A(n_13813),
.Y(n_14642)
);

AO32x2_ASAP7_75t_L g14643 ( 
.A1(n_13682),
.A2(n_9891),
.A3(n_9956),
.B1(n_9349),
.B2(n_13743),
.Y(n_14643)
);

NOR2x1_ASAP7_75t_SL g14644 ( 
.A(n_13065),
.B(n_9004),
.Y(n_14644)
);

AND2x2_ASAP7_75t_L g14645 ( 
.A(n_13708),
.B(n_12325),
.Y(n_14645)
);

AOI22xp5_ASAP7_75t_L g14646 ( 
.A1(n_13397),
.A2(n_10424),
.B1(n_11137),
.B2(n_11118),
.Y(n_14646)
);

NOR2xp33_ASAP7_75t_L g14647 ( 
.A(n_13813),
.B(n_10625),
.Y(n_14647)
);

NAND2xp33_ASAP7_75t_L g14648 ( 
.A(n_13775),
.B(n_9965),
.Y(n_14648)
);

AND2x2_ASAP7_75t_L g14649 ( 
.A(n_13722),
.B(n_12329),
.Y(n_14649)
);

AND2x2_ASAP7_75t_L g14650 ( 
.A(n_13722),
.B(n_12339),
.Y(n_14650)
);

BUFx3_ASAP7_75t_L g14651 ( 
.A(n_13476),
.Y(n_14651)
);

AOI221xp5_ASAP7_75t_L g14652 ( 
.A1(n_13144),
.A2(n_11579),
.B1(n_11569),
.B2(n_11137),
.C(n_11118),
.Y(n_14652)
);

NAND2xp5_ASAP7_75t_L g14653 ( 
.A(n_13678),
.B(n_9514),
.Y(n_14653)
);

INVx1_ASAP7_75t_L g14654 ( 
.A(n_13145),
.Y(n_14654)
);

A2O1A1Ixp33_ASAP7_75t_L g14655 ( 
.A1(n_13789),
.A2(n_9237),
.B(n_9256),
.C(n_9204),
.Y(n_14655)
);

OA21x2_ASAP7_75t_L g14656 ( 
.A1(n_13090),
.A2(n_11626),
.B(n_11609),
.Y(n_14656)
);

INVx2_ASAP7_75t_L g14657 ( 
.A(n_13574),
.Y(n_14657)
);

AND4x1_ASAP7_75t_L g14658 ( 
.A(n_13148),
.B(n_8611),
.C(n_8546),
.D(n_8151),
.Y(n_14658)
);

OAI21xp5_ASAP7_75t_L g14659 ( 
.A1(n_13925),
.A2(n_10688),
.B(n_10670),
.Y(n_14659)
);

AOI22xp33_ASAP7_75t_L g14660 ( 
.A1(n_13874),
.A2(n_9965),
.B1(n_10345),
.B2(n_10810),
.Y(n_14660)
);

AO21x2_ASAP7_75t_L g14661 ( 
.A1(n_13090),
.A2(n_11249),
.B(n_10742),
.Y(n_14661)
);

NOR2xp33_ASAP7_75t_L g14662 ( 
.A(n_13836),
.B(n_10625),
.Y(n_14662)
);

AND2x2_ASAP7_75t_L g14663 ( 
.A(n_13724),
.B(n_12354),
.Y(n_14663)
);

AO21x1_ASAP7_75t_L g14664 ( 
.A1(n_13134),
.A2(n_10340),
.B(n_10742),
.Y(n_14664)
);

OAI22xp5_ASAP7_75t_L g14665 ( 
.A1(n_13782),
.A2(n_9237),
.B1(n_9256),
.B2(n_9204),
.Y(n_14665)
);

INVx1_ASAP7_75t_L g14666 ( 
.A(n_13149),
.Y(n_14666)
);

INVx1_ASAP7_75t_L g14667 ( 
.A(n_12912),
.Y(n_14667)
);

OAI21x1_ASAP7_75t_SL g14668 ( 
.A1(n_13659),
.A2(n_9662),
.B(n_11660),
.Y(n_14668)
);

INVx2_ASAP7_75t_L g14669 ( 
.A(n_13761),
.Y(n_14669)
);

AND2x4_ASAP7_75t_L g14670 ( 
.A(n_13836),
.B(n_11577),
.Y(n_14670)
);

AND2x2_ASAP7_75t_L g14671 ( 
.A(n_13724),
.B(n_12356),
.Y(n_14671)
);

OAI22xp5_ASAP7_75t_L g14672 ( 
.A1(n_13495),
.A2(n_13505),
.B1(n_13522),
.B2(n_13519),
.Y(n_14672)
);

BUFx2_ASAP7_75t_L g14673 ( 
.A(n_13003),
.Y(n_14673)
);

AND2x2_ASAP7_75t_L g14674 ( 
.A(n_13580),
.B(n_12379),
.Y(n_14674)
);

AND2x6_ASAP7_75t_L g14675 ( 
.A(n_13850),
.B(n_13476),
.Y(n_14675)
);

AND2x2_ASAP7_75t_L g14676 ( 
.A(n_13592),
.B(n_12381),
.Y(n_14676)
);

AND2x2_ASAP7_75t_L g14677 ( 
.A(n_13603),
.B(n_12386),
.Y(n_14677)
);

AND2x2_ASAP7_75t_L g14678 ( 
.A(n_13655),
.B(n_12390),
.Y(n_14678)
);

AO32x2_ASAP7_75t_L g14679 ( 
.A1(n_13682),
.A2(n_9956),
.A3(n_9891),
.B1(n_8589),
.B2(n_12187),
.Y(n_14679)
);

AND2x2_ASAP7_75t_L g14680 ( 
.A(n_13045),
.B(n_12403),
.Y(n_14680)
);

OAI21xp5_ASAP7_75t_L g14681 ( 
.A1(n_13253),
.A2(n_10670),
.B(n_10803),
.Y(n_14681)
);

AND2x2_ASAP7_75t_L g14682 ( 
.A(n_13045),
.B(n_12413),
.Y(n_14682)
);

OR2x2_ASAP7_75t_L g14683 ( 
.A(n_13680),
.B(n_11594),
.Y(n_14683)
);

AOI22xp5_ASAP7_75t_L g14684 ( 
.A1(n_13273),
.A2(n_10424),
.B1(n_11137),
.B2(n_11118),
.Y(n_14684)
);

OA21x2_ASAP7_75t_L g14685 ( 
.A1(n_13134),
.A2(n_11626),
.B(n_11609),
.Y(n_14685)
);

OR2x2_ASAP7_75t_L g14686 ( 
.A(n_13684),
.B(n_11594),
.Y(n_14686)
);

INVx1_ASAP7_75t_L g14687 ( 
.A(n_12914),
.Y(n_14687)
);

OR2x2_ASAP7_75t_L g14688 ( 
.A(n_13687),
.B(n_11594),
.Y(n_14688)
);

OR2x2_ASAP7_75t_L g14689 ( 
.A(n_13560),
.B(n_11594),
.Y(n_14689)
);

AND2x2_ASAP7_75t_L g14690 ( 
.A(n_13068),
.B(n_12417),
.Y(n_14690)
);

AND2x2_ASAP7_75t_L g14691 ( 
.A(n_13068),
.B(n_12425),
.Y(n_14691)
);

BUFx3_ASAP7_75t_L g14692 ( 
.A(n_13836),
.Y(n_14692)
);

AND2x2_ASAP7_75t_L g14693 ( 
.A(n_13087),
.B(n_12432),
.Y(n_14693)
);

AND2x4_ASAP7_75t_L g14694 ( 
.A(n_13976),
.B(n_11591),
.Y(n_14694)
);

OAI22xp5_ASAP7_75t_L g14695 ( 
.A1(n_13505),
.A2(n_9256),
.B1(n_9267),
.B2(n_9237),
.Y(n_14695)
);

INVx2_ASAP7_75t_L g14696 ( 
.A(n_13761),
.Y(n_14696)
);

AOI22x1_ASAP7_75t_SL g14697 ( 
.A1(n_13961),
.A2(n_10907),
.B1(n_10986),
.B2(n_10759),
.Y(n_14697)
);

OAI22xp5_ASAP7_75t_L g14698 ( 
.A1(n_13519),
.A2(n_9256),
.B1(n_9267),
.B2(n_9237),
.Y(n_14698)
);

OR2x2_ASAP7_75t_L g14699 ( 
.A(n_13692),
.B(n_11594),
.Y(n_14699)
);

OR2x6_ASAP7_75t_L g14700 ( 
.A(n_13976),
.B(n_13850),
.Y(n_14700)
);

OR2x2_ASAP7_75t_L g14701 ( 
.A(n_13693),
.B(n_11594),
.Y(n_14701)
);

OA21x2_ASAP7_75t_L g14702 ( 
.A1(n_13210),
.A2(n_11626),
.B(n_11609),
.Y(n_14702)
);

OR2x2_ASAP7_75t_L g14703 ( 
.A(n_13694),
.B(n_10211),
.Y(n_14703)
);

NAND2xp5_ASAP7_75t_L g14704 ( 
.A(n_13715),
.B(n_9514),
.Y(n_14704)
);

OAI22xp5_ASAP7_75t_L g14705 ( 
.A1(n_13522),
.A2(n_13441),
.B1(n_13976),
.B2(n_13372),
.Y(n_14705)
);

BUFx3_ASAP7_75t_L g14706 ( 
.A(n_13966),
.Y(n_14706)
);

A2O1A1Ixp33_ASAP7_75t_L g14707 ( 
.A1(n_13838),
.A2(n_13422),
.B(n_13449),
.C(n_13433),
.Y(n_14707)
);

AND2x4_ASAP7_75t_SL g14708 ( 
.A(n_13918),
.B(n_9608),
.Y(n_14708)
);

A2O1A1Ixp33_ASAP7_75t_L g14709 ( 
.A1(n_13506),
.A2(n_9267),
.B(n_9297),
.C(n_9256),
.Y(n_14709)
);

AND2x2_ASAP7_75t_L g14710 ( 
.A(n_13087),
.B(n_12438),
.Y(n_14710)
);

AND2x2_ASAP7_75t_L g14711 ( 
.A(n_13097),
.B(n_10443),
.Y(n_14711)
);

OR2x2_ASAP7_75t_L g14712 ( 
.A(n_13716),
.B(n_10211),
.Y(n_14712)
);

BUFx12f_ASAP7_75t_L g14713 ( 
.A(n_13850),
.Y(n_14713)
);

AO21x2_ASAP7_75t_L g14714 ( 
.A1(n_13210),
.A2(n_13814),
.B(n_13743),
.Y(n_14714)
);

OR2x2_ASAP7_75t_L g14715 ( 
.A(n_13725),
.B(n_10211),
.Y(n_14715)
);

AOI221xp5_ASAP7_75t_L g14716 ( 
.A1(n_13728),
.A2(n_11569),
.B1(n_11579),
.B2(n_11137),
.C(n_11118),
.Y(n_14716)
);

A2O1A1Ixp33_ASAP7_75t_L g14717 ( 
.A1(n_13523),
.A2(n_13234),
.B(n_13198),
.C(n_13162),
.Y(n_14717)
);

OAI22xp5_ASAP7_75t_SL g14718 ( 
.A1(n_13918),
.A2(n_9267),
.B1(n_9297),
.B2(n_9256),
.Y(n_14718)
);

OR2x2_ASAP7_75t_L g14719 ( 
.A(n_13731),
.B(n_10211),
.Y(n_14719)
);

INVx1_ASAP7_75t_L g14720 ( 
.A(n_12915),
.Y(n_14720)
);

INVxp67_ASAP7_75t_L g14721 ( 
.A(n_13978),
.Y(n_14721)
);

INVxp33_ASAP7_75t_L g14722 ( 
.A(n_13663),
.Y(n_14722)
);

AND2x4_ASAP7_75t_SL g14723 ( 
.A(n_13581),
.B(n_9608),
.Y(n_14723)
);

AOI22xp5_ASAP7_75t_L g14724 ( 
.A1(n_13273),
.A2(n_13972),
.B1(n_13973),
.B2(n_13496),
.Y(n_14724)
);

INVx2_ASAP7_75t_L g14725 ( 
.A(n_13773),
.Y(n_14725)
);

NOR2xp33_ASAP7_75t_L g14726 ( 
.A(n_13963),
.B(n_13039),
.Y(n_14726)
);

OAI21xp5_ASAP7_75t_L g14727 ( 
.A1(n_13046),
.A2(n_10799),
.B(n_10769),
.Y(n_14727)
);

AO32x2_ASAP7_75t_L g14728 ( 
.A1(n_13539),
.A2(n_9956),
.A3(n_8589),
.B1(n_12215),
.B2(n_8657),
.Y(n_14728)
);

A2O1A1Ixp33_ASAP7_75t_L g14729 ( 
.A1(n_13530),
.A2(n_9297),
.B(n_9350),
.C(n_9267),
.Y(n_14729)
);

A2O1A1Ixp33_ASAP7_75t_L g14730 ( 
.A1(n_13543),
.A2(n_9297),
.B(n_9350),
.C(n_9267),
.Y(n_14730)
);

NOR2xp33_ASAP7_75t_L g14731 ( 
.A(n_13048),
.B(n_10759),
.Y(n_14731)
);

AND2x2_ASAP7_75t_L g14732 ( 
.A(n_13097),
.B(n_10443),
.Y(n_14732)
);

OR2x2_ASAP7_75t_L g14733 ( 
.A(n_13856),
.B(n_10211),
.Y(n_14733)
);

NOR2xp33_ASAP7_75t_L g14734 ( 
.A(n_13985),
.B(n_13863),
.Y(n_14734)
);

AND2x4_ASAP7_75t_L g14735 ( 
.A(n_13773),
.B(n_11591),
.Y(n_14735)
);

INVx1_ASAP7_75t_L g14736 ( 
.A(n_12920),
.Y(n_14736)
);

AND2x2_ASAP7_75t_L g14737 ( 
.A(n_13272),
.B(n_10443),
.Y(n_14737)
);

AND2x4_ASAP7_75t_L g14738 ( 
.A(n_13851),
.B(n_11591),
.Y(n_14738)
);

OAI21x1_ASAP7_75t_L g14739 ( 
.A1(n_13742),
.A2(n_12786),
.B(n_12694),
.Y(n_14739)
);

BUFx3_ASAP7_75t_L g14740 ( 
.A(n_13851),
.Y(n_14740)
);

A2O1A1Ixp33_ASAP7_75t_L g14741 ( 
.A1(n_13156),
.A2(n_9350),
.B(n_9297),
.C(n_9845),
.Y(n_14741)
);

CKINVDCx6p67_ASAP7_75t_R g14742 ( 
.A(n_13496),
.Y(n_14742)
);

OA21x2_ASAP7_75t_L g14743 ( 
.A1(n_13970),
.A2(n_11249),
.B(n_10944),
.Y(n_14743)
);

INVx1_ASAP7_75t_L g14744 ( 
.A(n_12925),
.Y(n_14744)
);

OR2x2_ASAP7_75t_L g14745 ( 
.A(n_13864),
.B(n_10211),
.Y(n_14745)
);

OAI21xp5_ASAP7_75t_L g14746 ( 
.A1(n_12984),
.A2(n_10799),
.B(n_10769),
.Y(n_14746)
);

NOR2x1_ASAP7_75t_L g14747 ( 
.A(n_13555),
.B(n_13614),
.Y(n_14747)
);

AND2x4_ASAP7_75t_L g14748 ( 
.A(n_13879),
.B(n_11591),
.Y(n_14748)
);

AO32x2_ASAP7_75t_L g14749 ( 
.A1(n_13539),
.A2(n_8657),
.A3(n_11911),
.B1(n_11847),
.B2(n_11824),
.Y(n_14749)
);

INVx1_ASAP7_75t_L g14750 ( 
.A(n_12926),
.Y(n_14750)
);

AO32x1_ASAP7_75t_L g14751 ( 
.A1(n_13025),
.A2(n_11249),
.A3(n_9787),
.B1(n_9843),
.B2(n_9809),
.Y(n_14751)
);

AND2x2_ASAP7_75t_L g14752 ( 
.A(n_13272),
.B(n_10443),
.Y(n_14752)
);

AND2x2_ASAP7_75t_L g14753 ( 
.A(n_13312),
.B(n_13317),
.Y(n_14753)
);

AO21x1_ASAP7_75t_L g14754 ( 
.A1(n_13584),
.A2(n_10340),
.B(n_11554),
.Y(n_14754)
);

AND2x2_ASAP7_75t_L g14755 ( 
.A(n_13312),
.B(n_10478),
.Y(n_14755)
);

BUFx3_ASAP7_75t_L g14756 ( 
.A(n_13879),
.Y(n_14756)
);

OAI21xp5_ASAP7_75t_L g14757 ( 
.A1(n_12988),
.A2(n_10799),
.B(n_10769),
.Y(n_14757)
);

AND2x2_ASAP7_75t_L g14758 ( 
.A(n_13317),
.B(n_10478),
.Y(n_14758)
);

NOR2x1_ASAP7_75t_SL g14759 ( 
.A(n_13065),
.B(n_9004),
.Y(n_14759)
);

A2O1A1Ixp33_ASAP7_75t_L g14760 ( 
.A1(n_13169),
.A2(n_9350),
.B(n_9297),
.C(n_9845),
.Y(n_14760)
);

INVx2_ASAP7_75t_L g14761 ( 
.A(n_13921),
.Y(n_14761)
);

AOI221xp5_ASAP7_75t_L g14762 ( 
.A1(n_13880),
.A2(n_13878),
.B1(n_13865),
.B2(n_13719),
.C(n_13020),
.Y(n_14762)
);

CKINVDCx20_ASAP7_75t_R g14763 ( 
.A(n_13667),
.Y(n_14763)
);

AOI21xp5_ASAP7_75t_L g14764 ( 
.A1(n_13614),
.A2(n_10707),
.B(n_10657),
.Y(n_14764)
);

AND2x2_ASAP7_75t_L g14765 ( 
.A(n_13319),
.B(n_10478),
.Y(n_14765)
);

A2O1A1Ixp33_ASAP7_75t_L g14766 ( 
.A1(n_13464),
.A2(n_9350),
.B(n_9849),
.C(n_9845),
.Y(n_14766)
);

OR2x2_ASAP7_75t_L g14767 ( 
.A(n_13658),
.B(n_10211),
.Y(n_14767)
);

OR2x2_ASAP7_75t_L g14768 ( 
.A(n_13568),
.B(n_10211),
.Y(n_14768)
);

AND2x4_ASAP7_75t_L g14769 ( 
.A(n_13921),
.B(n_11591),
.Y(n_14769)
);

NOR2xp33_ASAP7_75t_L g14770 ( 
.A(n_13319),
.B(n_10759),
.Y(n_14770)
);

INVxp67_ASAP7_75t_L g14771 ( 
.A(n_13006),
.Y(n_14771)
);

AO32x2_ASAP7_75t_L g14772 ( 
.A1(n_13621),
.A2(n_13488),
.A3(n_13645),
.B1(n_13957),
.B2(n_13719),
.Y(n_14772)
);

AND2x4_ASAP7_75t_L g14773 ( 
.A(n_13949),
.B(n_11623),
.Y(n_14773)
);

NOR2x1_ASAP7_75t_R g14774 ( 
.A(n_13695),
.B(n_13703),
.Y(n_14774)
);

AOI22xp5_ASAP7_75t_L g14775 ( 
.A1(n_13884),
.A2(n_10438),
.B1(n_10451),
.B2(n_11569),
.Y(n_14775)
);

INVx5_ASAP7_75t_L g14776 ( 
.A(n_13949),
.Y(n_14776)
);

INVx2_ASAP7_75t_L g14777 ( 
.A(n_13695),
.Y(n_14777)
);

INVx3_ASAP7_75t_SL g14778 ( 
.A(n_13703),
.Y(n_14778)
);

INVxp67_ASAP7_75t_L g14779 ( 
.A(n_13010),
.Y(n_14779)
);

INVx1_ASAP7_75t_L g14780 ( 
.A(n_12944),
.Y(n_14780)
);

OAI22xp5_ASAP7_75t_L g14781 ( 
.A1(n_13441),
.A2(n_9350),
.B1(n_9035),
.B2(n_9044),
.Y(n_14781)
);

OA21x2_ASAP7_75t_L g14782 ( 
.A1(n_13965),
.A2(n_13980),
.B(n_13975),
.Y(n_14782)
);

AND2x2_ASAP7_75t_L g14783 ( 
.A(n_13674),
.B(n_10478),
.Y(n_14783)
);

OA21x2_ASAP7_75t_L g14784 ( 
.A1(n_13984),
.A2(n_10944),
.B(n_10855),
.Y(n_14784)
);

OR2x6_ASAP7_75t_L g14785 ( 
.A(n_13379),
.B(n_10178),
.Y(n_14785)
);

BUFx3_ASAP7_75t_L g14786 ( 
.A(n_12911),
.Y(n_14786)
);

OAI22xp5_ASAP7_75t_SL g14787 ( 
.A1(n_12919),
.A2(n_9017),
.B1(n_9044),
.B2(n_9035),
.Y(n_14787)
);

AND2x2_ASAP7_75t_L g14788 ( 
.A(n_13697),
.B(n_10478),
.Y(n_14788)
);

AND2x2_ASAP7_75t_L g14789 ( 
.A(n_13749),
.B(n_10480),
.Y(n_14789)
);

O2A1O1Ixp33_ASAP7_75t_L g14790 ( 
.A1(n_13621),
.A2(n_11492),
.B(n_11513),
.C(n_11371),
.Y(n_14790)
);

AND2x4_ASAP7_75t_L g14791 ( 
.A(n_13785),
.B(n_11623),
.Y(n_14791)
);

OAI21x1_ASAP7_75t_L g14792 ( 
.A1(n_13482),
.A2(n_13140),
.B(n_13793),
.Y(n_14792)
);

AND2x4_ASAP7_75t_L g14793 ( 
.A(n_13840),
.B(n_11623),
.Y(n_14793)
);

OAI22xp5_ASAP7_75t_L g14794 ( 
.A1(n_13372),
.A2(n_9035),
.B1(n_9044),
.B2(n_9017),
.Y(n_14794)
);

AND2x2_ASAP7_75t_L g14795 ( 
.A(n_13855),
.B(n_10480),
.Y(n_14795)
);

OAI21xp5_ASAP7_75t_L g14796 ( 
.A1(n_13373),
.A2(n_13418),
.B(n_13408),
.Y(n_14796)
);

AND2x2_ASAP7_75t_L g14797 ( 
.A(n_13872),
.B(n_10480),
.Y(n_14797)
);

AND2x2_ASAP7_75t_L g14798 ( 
.A(n_13877),
.B(n_10480),
.Y(n_14798)
);

INVx1_ASAP7_75t_L g14799 ( 
.A(n_12951),
.Y(n_14799)
);

NOR2xp33_ASAP7_75t_L g14800 ( 
.A(n_13455),
.B(n_10759),
.Y(n_14800)
);

A2O1A1Ixp33_ASAP7_75t_L g14801 ( 
.A1(n_13598),
.A2(n_9849),
.B(n_9865),
.C(n_9845),
.Y(n_14801)
);

NAND2xp5_ASAP7_75t_L g14802 ( 
.A(n_13547),
.B(n_9514),
.Y(n_14802)
);

AND2x2_ASAP7_75t_L g14803 ( 
.A(n_13881),
.B(n_10480),
.Y(n_14803)
);

A2O1A1Ixp33_ASAP7_75t_L g14804 ( 
.A1(n_13982),
.A2(n_9849),
.B(n_9865),
.C(n_9845),
.Y(n_14804)
);

OAI21x1_ASAP7_75t_L g14805 ( 
.A1(n_13907),
.A2(n_12811),
.B(n_12805),
.Y(n_14805)
);

AND2x4_ASAP7_75t_L g14806 ( 
.A(n_13886),
.B(n_11623),
.Y(n_14806)
);

CKINVDCx5p33_ASAP7_75t_R g14807 ( 
.A(n_13379),
.Y(n_14807)
);

O2A1O1Ixp33_ASAP7_75t_L g14808 ( 
.A1(n_13021),
.A2(n_11492),
.B(n_11513),
.C(n_11371),
.Y(n_14808)
);

NOR2xp33_ASAP7_75t_L g14809 ( 
.A(n_13456),
.B(n_10759),
.Y(n_14809)
);

INVx1_ASAP7_75t_L g14810 ( 
.A(n_12953),
.Y(n_14810)
);

AOI221xp5_ASAP7_75t_L g14811 ( 
.A1(n_13022),
.A2(n_11579),
.B1(n_11569),
.B2(n_11513),
.C(n_11550),
.Y(n_14811)
);

AOI22xp5_ASAP7_75t_L g14812 ( 
.A1(n_13890),
.A2(n_10438),
.B1(n_10451),
.B2(n_11579),
.Y(n_14812)
);

INVx2_ASAP7_75t_L g14813 ( 
.A(n_12922),
.Y(n_14813)
);

AND2x2_ASAP7_75t_L g14814 ( 
.A(n_13887),
.B(n_10525),
.Y(n_14814)
);

AND2x2_ASAP7_75t_L g14815 ( 
.A(n_13951),
.B(n_13981),
.Y(n_14815)
);

AND2x2_ASAP7_75t_L g14816 ( 
.A(n_13063),
.B(n_10525),
.Y(n_14816)
);

AOI221xp5_ASAP7_75t_L g14817 ( 
.A1(n_13027),
.A2(n_11550),
.B1(n_11559),
.B2(n_11492),
.C(n_11371),
.Y(n_14817)
);

AND2x2_ASAP7_75t_L g14818 ( 
.A(n_13069),
.B(n_13151),
.Y(n_14818)
);

OR2x2_ASAP7_75t_L g14819 ( 
.A(n_13569),
.B(n_13583),
.Y(n_14819)
);

AND2x2_ASAP7_75t_L g14820 ( 
.A(n_13155),
.B(n_10525),
.Y(n_14820)
);

INVx1_ASAP7_75t_L g14821 ( 
.A(n_12954),
.Y(n_14821)
);

BUFx8_ASAP7_75t_SL g14822 ( 
.A(n_13158),
.Y(n_14822)
);

A2O1A1Ixp33_ASAP7_75t_L g14823 ( 
.A1(n_13360),
.A2(n_9849),
.B(n_9865),
.C(n_9845),
.Y(n_14823)
);

AOI221xp5_ASAP7_75t_L g14824 ( 
.A1(n_13030),
.A2(n_11560),
.B1(n_11559),
.B2(n_11550),
.C(n_10657),
.Y(n_14824)
);

AO21x1_ASAP7_75t_L g14825 ( 
.A1(n_13584),
.A2(n_10340),
.B(n_11554),
.Y(n_14825)
);

OR2x2_ASAP7_75t_L g14826 ( 
.A(n_13619),
.B(n_10217),
.Y(n_14826)
);

INVx1_ASAP7_75t_L g14827 ( 
.A(n_12957),
.Y(n_14827)
);

OA21x2_ASAP7_75t_L g14828 ( 
.A1(n_13987),
.A2(n_10944),
.B(n_10855),
.Y(n_14828)
);

AO32x1_ASAP7_75t_L g14829 ( 
.A1(n_13033),
.A2(n_9787),
.A3(n_9843),
.B1(n_9809),
.B2(n_9796),
.Y(n_14829)
);

OAI21xp5_ASAP7_75t_L g14830 ( 
.A1(n_13368),
.A2(n_10799),
.B(n_10769),
.Y(n_14830)
);

NOR2xp33_ASAP7_75t_L g14831 ( 
.A(n_13465),
.B(n_10907),
.Y(n_14831)
);

INVx3_ASAP7_75t_L g14832 ( 
.A(n_13387),
.Y(n_14832)
);

INVx2_ASAP7_75t_L g14833 ( 
.A(n_12929),
.Y(n_14833)
);

AO22x2_ASAP7_75t_L g14834 ( 
.A1(n_13032),
.A2(n_11559),
.B1(n_11560),
.B2(n_11554),
.Y(n_14834)
);

AND2x4_ASAP7_75t_L g14835 ( 
.A(n_13469),
.B(n_13479),
.Y(n_14835)
);

CKINVDCx5p33_ASAP7_75t_R g14836 ( 
.A(n_13387),
.Y(n_14836)
);

INVx1_ASAP7_75t_L g14837 ( 
.A(n_12959),
.Y(n_14837)
);

OAI21xp5_ASAP7_75t_L g14838 ( 
.A1(n_13957),
.A2(n_12955),
.B(n_13019),
.Y(n_14838)
);

INVx2_ASAP7_75t_L g14839 ( 
.A(n_12930),
.Y(n_14839)
);

AND2x4_ASAP7_75t_L g14840 ( 
.A(n_13480),
.B(n_11623),
.Y(n_14840)
);

AND2x2_ASAP7_75t_L g14841 ( 
.A(n_13159),
.B(n_10525),
.Y(n_14841)
);

INVxp67_ASAP7_75t_L g14842 ( 
.A(n_13034),
.Y(n_14842)
);

INVx1_ASAP7_75t_L g14843 ( 
.A(n_12968),
.Y(n_14843)
);

AOI21xp5_ASAP7_75t_L g14844 ( 
.A1(n_13645),
.A2(n_10710),
.B(n_10657),
.Y(n_14844)
);

A2O1A1Ixp33_ASAP7_75t_L g14845 ( 
.A1(n_13249),
.A2(n_9865),
.B(n_9947),
.C(n_9849),
.Y(n_14845)
);

INVx1_ASAP7_75t_L g14846 ( 
.A(n_12971),
.Y(n_14846)
);

INVx1_ASAP7_75t_L g14847 ( 
.A(n_12973),
.Y(n_14847)
);

OR2x6_ASAP7_75t_L g14848 ( 
.A(n_13709),
.B(n_9005),
.Y(n_14848)
);

OAI21xp5_ASAP7_75t_L g14849 ( 
.A1(n_12955),
.A2(n_10280),
.B(n_10459),
.Y(n_14849)
);

AOI211xp5_ASAP7_75t_L g14850 ( 
.A1(n_13035),
.A2(n_10753),
.B(n_10821),
.C(n_10711),
.Y(n_14850)
);

INVxp33_ASAP7_75t_L g14851 ( 
.A(n_13489),
.Y(n_14851)
);

NAND2x1_ASAP7_75t_L g14852 ( 
.A(n_13710),
.B(n_13986),
.Y(n_14852)
);

INVx1_ASAP7_75t_L g14853 ( 
.A(n_12975),
.Y(n_14853)
);

HB1xp67_ASAP7_75t_L g14854 ( 
.A(n_13044),
.Y(n_14854)
);

AND2x2_ASAP7_75t_L g14855 ( 
.A(n_13163),
.B(n_10525),
.Y(n_14855)
);

INVx3_ASAP7_75t_L g14856 ( 
.A(n_12931),
.Y(n_14856)
);

AND2x2_ASAP7_75t_L g14857 ( 
.A(n_13168),
.B(n_10576),
.Y(n_14857)
);

OR2x2_ASAP7_75t_L g14858 ( 
.A(n_13620),
.B(n_10217),
.Y(n_14858)
);

INVx4_ASAP7_75t_L g14859 ( 
.A(n_12935),
.Y(n_14859)
);

AND2x2_ASAP7_75t_L g14860 ( 
.A(n_13170),
.B(n_10576),
.Y(n_14860)
);

AOI221xp5_ASAP7_75t_L g14861 ( 
.A1(n_13047),
.A2(n_11560),
.B1(n_10710),
.B2(n_11007),
.C(n_10762),
.Y(n_14861)
);

AND2x2_ASAP7_75t_L g14862 ( 
.A(n_13174),
.B(n_10576),
.Y(n_14862)
);

NAND2xp5_ASAP7_75t_L g14863 ( 
.A(n_13178),
.B(n_9514),
.Y(n_14863)
);

AOI22xp33_ASAP7_75t_L g14864 ( 
.A1(n_13895),
.A2(n_9965),
.B1(n_10345),
.B2(n_10810),
.Y(n_14864)
);

CKINVDCx5p33_ASAP7_75t_R g14865 ( 
.A(n_13302),
.Y(n_14865)
);

OR2x2_ASAP7_75t_L g14866 ( 
.A(n_13624),
.B(n_13631),
.Y(n_14866)
);

OA21x2_ASAP7_75t_L g14867 ( 
.A1(n_13814),
.A2(n_10859),
.B(n_10853),
.Y(n_14867)
);

NOR2xp33_ASAP7_75t_L g14868 ( 
.A(n_13490),
.B(n_13513),
.Y(n_14868)
);

INVx1_ASAP7_75t_L g14869 ( 
.A(n_12991),
.Y(n_14869)
);

BUFx3_ASAP7_75t_L g14870 ( 
.A(n_12948),
.Y(n_14870)
);

NOR2x1_ASAP7_75t_L g14871 ( 
.A(n_12952),
.B(n_9017),
.Y(n_14871)
);

OAI21xp5_ASAP7_75t_L g14872 ( 
.A1(n_13019),
.A2(n_10280),
.B(n_10459),
.Y(n_14872)
);

OAI21xp5_ASAP7_75t_L g14873 ( 
.A1(n_13050),
.A2(n_10280),
.B(n_10459),
.Y(n_14873)
);

AND2x2_ASAP7_75t_L g14874 ( 
.A(n_13179),
.B(n_10576),
.Y(n_14874)
);

OR2x2_ASAP7_75t_L g14875 ( 
.A(n_13632),
.B(n_10217),
.Y(n_14875)
);

A2O1A1Ixp33_ASAP7_75t_L g14876 ( 
.A1(n_12983),
.A2(n_9865),
.B(n_9947),
.C(n_9849),
.Y(n_14876)
);

OA21x2_ASAP7_75t_L g14877 ( 
.A1(n_13252),
.A2(n_10860),
.B(n_10859),
.Y(n_14877)
);

OR2x2_ASAP7_75t_L g14878 ( 
.A(n_13634),
.B(n_10217),
.Y(n_14878)
);

NAND2xp5_ASAP7_75t_L g14879 ( 
.A(n_13181),
.B(n_9514),
.Y(n_14879)
);

AND2x2_ASAP7_75t_L g14880 ( 
.A(n_13182),
.B(n_10576),
.Y(n_14880)
);

AOI221xp5_ASAP7_75t_L g14881 ( 
.A1(n_13727),
.A2(n_10710),
.B1(n_11007),
.B2(n_10762),
.C(n_10451),
.Y(n_14881)
);

AND2x2_ASAP7_75t_L g14882 ( 
.A(n_13197),
.B(n_10613),
.Y(n_14882)
);

AOI21xp5_ASAP7_75t_L g14883 ( 
.A1(n_13488),
.A2(n_10710),
.B(n_10808),
.Y(n_14883)
);

A2O1A1Ixp33_ASAP7_75t_L g14884 ( 
.A1(n_13016),
.A2(n_9865),
.B(n_9947),
.C(n_9849),
.Y(n_14884)
);

AND2x2_ASAP7_75t_L g14885 ( 
.A(n_13219),
.B(n_10613),
.Y(n_14885)
);

NOR2x1_ASAP7_75t_SL g14886 ( 
.A(n_12952),
.B(n_9017),
.Y(n_14886)
);

AOI21xp5_ASAP7_75t_L g14887 ( 
.A1(n_13741),
.A2(n_10710),
.B(n_10808),
.Y(n_14887)
);

HB1xp67_ASAP7_75t_L g14888 ( 
.A(n_12997),
.Y(n_14888)
);

INVx1_ASAP7_75t_L g14889 ( 
.A(n_12999),
.Y(n_14889)
);

OAI21x1_ASAP7_75t_SL g14890 ( 
.A1(n_13050),
.A2(n_9662),
.B(n_11660),
.Y(n_14890)
);

BUFx6f_ASAP7_75t_L g14891 ( 
.A(n_12989),
.Y(n_14891)
);

CKINVDCx5p33_ASAP7_75t_R g14892 ( 
.A(n_13314),
.Y(n_14892)
);

NAND3xp33_ASAP7_75t_L g14893 ( 
.A(n_12919),
.B(n_9283),
.C(n_10766),
.Y(n_14893)
);

INVx1_ASAP7_75t_L g14894 ( 
.A(n_13004),
.Y(n_14894)
);

AND2x2_ASAP7_75t_L g14895 ( 
.A(n_13226),
.B(n_10613),
.Y(n_14895)
);

A2O1A1Ixp33_ASAP7_75t_L g14896 ( 
.A1(n_13225),
.A2(n_9865),
.B(n_9947),
.C(n_9849),
.Y(n_14896)
);

INVx1_ASAP7_75t_L g14897 ( 
.A(n_13150),
.Y(n_14897)
);

NOR2x1_ASAP7_75t_SL g14898 ( 
.A(n_13406),
.B(n_13582),
.Y(n_14898)
);

INVxp67_ASAP7_75t_L g14899 ( 
.A(n_12990),
.Y(n_14899)
);

AOI22xp33_ASAP7_75t_L g14900 ( 
.A1(n_13910),
.A2(n_9965),
.B1(n_10345),
.B2(n_10810),
.Y(n_14900)
);

AND2x2_ASAP7_75t_L g14901 ( 
.A(n_13227),
.B(n_10613),
.Y(n_14901)
);

INVx4_ASAP7_75t_L g14902 ( 
.A(n_12994),
.Y(n_14902)
);

A2O1A1Ixp33_ASAP7_75t_L g14903 ( 
.A1(n_13848),
.A2(n_9947),
.B(n_10132),
.C(n_9865),
.Y(n_14903)
);

NAND2xp5_ASAP7_75t_L g14904 ( 
.A(n_13243),
.B(n_13245),
.Y(n_14904)
);

NAND2xp5_ASAP7_75t_L g14905 ( 
.A(n_13251),
.B(n_9523),
.Y(n_14905)
);

OAI22xp5_ASAP7_75t_L g14906 ( 
.A1(n_13848),
.A2(n_9035),
.B1(n_9044),
.B2(n_9017),
.Y(n_14906)
);

NOR2xp33_ASAP7_75t_L g14907 ( 
.A(n_13515),
.B(n_13528),
.Y(n_14907)
);

O2A1O1Ixp33_ASAP7_75t_L g14908 ( 
.A1(n_13485),
.A2(n_10808),
.B(n_10762),
.C(n_10835),
.Y(n_14908)
);

AO32x2_ASAP7_75t_L g14909 ( 
.A1(n_13727),
.A2(n_12446),
.A3(n_12442),
.B1(n_8981),
.B2(n_9084),
.Y(n_14909)
);

NOR2x1_ASAP7_75t_SL g14910 ( 
.A(n_13741),
.B(n_9017),
.Y(n_14910)
);

A2O1A1Ixp33_ASAP7_75t_L g14911 ( 
.A1(n_13866),
.A2(n_10132),
.B(n_10154),
.C(n_9947),
.Y(n_14911)
);

AND2x2_ASAP7_75t_L g14912 ( 
.A(n_13255),
.B(n_10613),
.Y(n_14912)
);

O2A1O1Ixp33_ASAP7_75t_SL g14913 ( 
.A1(n_13252),
.A2(n_11066),
.B(n_11215),
.C(n_11033),
.Y(n_14913)
);

NAND2xp5_ASAP7_75t_L g14914 ( 
.A(n_13388),
.B(n_9523),
.Y(n_14914)
);

AOI221xp5_ASAP7_75t_L g14915 ( 
.A1(n_13774),
.A2(n_11007),
.B1(n_10762),
.B2(n_10451),
.C(n_10438),
.Y(n_14915)
);

OR2x6_ASAP7_75t_L g14916 ( 
.A(n_13534),
.B(n_9005),
.Y(n_14916)
);

OR2x2_ASAP7_75t_L g14917 ( 
.A(n_13638),
.B(n_13641),
.Y(n_14917)
);

O2A1O1Ixp33_ASAP7_75t_SL g14918 ( 
.A1(n_13284),
.A2(n_11215),
.B(n_11261),
.C(n_11066),
.Y(n_14918)
);

AND2x4_ASAP7_75t_L g14919 ( 
.A(n_13535),
.B(n_11357),
.Y(n_14919)
);

AND2x2_ASAP7_75t_L g14920 ( 
.A(n_13913),
.B(n_10777),
.Y(n_14920)
);

INVx3_ASAP7_75t_L g14921 ( 
.A(n_13088),
.Y(n_14921)
);

INVxp67_ASAP7_75t_L g14922 ( 
.A(n_13261),
.Y(n_14922)
);

INVx3_ASAP7_75t_L g14923 ( 
.A(n_13092),
.Y(n_14923)
);

AOI22xp5_ASAP7_75t_L g14924 ( 
.A1(n_13914),
.A2(n_10438),
.B1(n_10451),
.B2(n_10345),
.Y(n_14924)
);

AND2x4_ASAP7_75t_L g14925 ( 
.A(n_13927),
.B(n_11357),
.Y(n_14925)
);

A2O1A1Ixp33_ASAP7_75t_L g14926 ( 
.A1(n_13866),
.A2(n_10132),
.B(n_10154),
.C(n_9947),
.Y(n_14926)
);

NOR2xp33_ASAP7_75t_L g14927 ( 
.A(n_13956),
.B(n_10907),
.Y(n_14927)
);

AND2x2_ASAP7_75t_L g14928 ( 
.A(n_13958),
.B(n_10777),
.Y(n_14928)
);

OAI21xp5_ASAP7_75t_L g14929 ( 
.A1(n_12933),
.A2(n_10873),
.B(n_10872),
.Y(n_14929)
);

AOI21xp5_ASAP7_75t_L g14930 ( 
.A1(n_13774),
.A2(n_10760),
.B(n_10835),
.Y(n_14930)
);

BUFx6f_ASAP7_75t_L g14931 ( 
.A(n_13315),
.Y(n_14931)
);

AO32x2_ASAP7_75t_L g14932 ( 
.A1(n_13817),
.A2(n_8981),
.A3(n_9084),
.B1(n_12226),
.B2(n_12647),
.Y(n_14932)
);

INVx1_ASAP7_75t_L g14933 ( 
.A(n_13161),
.Y(n_14933)
);

AND2x2_ASAP7_75t_L g14934 ( 
.A(n_13717),
.B(n_10777),
.Y(n_14934)
);

AOI21xp5_ASAP7_75t_SL g14935 ( 
.A1(n_13485),
.A2(n_10804),
.B(n_10896),
.Y(n_14935)
);

AND2x4_ASAP7_75t_L g14936 ( 
.A(n_13723),
.B(n_11357),
.Y(n_14936)
);

AND2x2_ASAP7_75t_L g14937 ( 
.A(n_13726),
.B(n_13730),
.Y(n_14937)
);

BUFx4f_ASAP7_75t_L g14938 ( 
.A(n_13316),
.Y(n_14938)
);

AOI21xp5_ASAP7_75t_L g14939 ( 
.A1(n_13817),
.A2(n_10760),
.B(n_10835),
.Y(n_14939)
);

NOR2xp33_ASAP7_75t_SL g14940 ( 
.A(n_13268),
.B(n_10907),
.Y(n_14940)
);

HB1xp67_ASAP7_75t_L g14941 ( 
.A(n_13284),
.Y(n_14941)
);

NOR2xp33_ASAP7_75t_L g14942 ( 
.A(n_13732),
.B(n_10907),
.Y(n_14942)
);

AND2x2_ASAP7_75t_L g14943 ( 
.A(n_13736),
.B(n_10777),
.Y(n_14943)
);

INVx2_ASAP7_75t_L g14944 ( 
.A(n_13318),
.Y(n_14944)
);

OR2x2_ASAP7_75t_L g14945 ( 
.A(n_13649),
.B(n_10217),
.Y(n_14945)
);

AOI21xp5_ASAP7_75t_L g14946 ( 
.A1(n_13514),
.A2(n_10760),
.B(n_10835),
.Y(n_14946)
);

NOR2xp33_ASAP7_75t_L g14947 ( 
.A(n_13755),
.B(n_10986),
.Y(n_14947)
);

HB1xp67_ASAP7_75t_L g14948 ( 
.A(n_13299),
.Y(n_14948)
);

AND2x2_ASAP7_75t_L g14949 ( 
.A(n_13759),
.B(n_10777),
.Y(n_14949)
);

HB1xp67_ASAP7_75t_L g14950 ( 
.A(n_13299),
.Y(n_14950)
);

AND2x4_ASAP7_75t_SL g14951 ( 
.A(n_13772),
.B(n_9608),
.Y(n_14951)
);

AND2x2_ASAP7_75t_L g14952 ( 
.A(n_13776),
.B(n_10794),
.Y(n_14952)
);

NAND2xp5_ASAP7_75t_L g14953 ( 
.A(n_13389),
.B(n_9523),
.Y(n_14953)
);

INVx1_ASAP7_75t_L g14954 ( 
.A(n_13166),
.Y(n_14954)
);

A2O1A1Ixp33_ASAP7_75t_L g14955 ( 
.A1(n_13337),
.A2(n_10132),
.B(n_10154),
.C(n_9947),
.Y(n_14955)
);

INVx2_ASAP7_75t_SL g14956 ( 
.A(n_13714),
.Y(n_14956)
);

AND2x2_ASAP7_75t_L g14957 ( 
.A(n_13778),
.B(n_10794),
.Y(n_14957)
);

BUFx3_ASAP7_75t_L g14958 ( 
.A(n_13279),
.Y(n_14958)
);

OR2x6_ASAP7_75t_L g14959 ( 
.A(n_13322),
.B(n_9005),
.Y(n_14959)
);

OAI22xp5_ASAP7_75t_L g14960 ( 
.A1(n_13626),
.A2(n_9044),
.B1(n_9068),
.B2(n_9035),
.Y(n_14960)
);

INVx1_ASAP7_75t_L g14961 ( 
.A(n_13167),
.Y(n_14961)
);

AND2x2_ASAP7_75t_L g14962 ( 
.A(n_13791),
.B(n_10794),
.Y(n_14962)
);

INVx3_ASAP7_75t_L g14963 ( 
.A(n_13108),
.Y(n_14963)
);

AND2x2_ASAP7_75t_L g14964 ( 
.A(n_13794),
.B(n_10794),
.Y(n_14964)
);

BUFx2_ASAP7_75t_L g14965 ( 
.A(n_13714),
.Y(n_14965)
);

INVx1_ASAP7_75t_L g14966 ( 
.A(n_13171),
.Y(n_14966)
);

AND2x2_ASAP7_75t_L g14967 ( 
.A(n_13795),
.B(n_10794),
.Y(n_14967)
);

AND2x2_ASAP7_75t_L g14968 ( 
.A(n_13803),
.B(n_10829),
.Y(n_14968)
);

AND2x2_ASAP7_75t_L g14969 ( 
.A(n_13808),
.B(n_10829),
.Y(n_14969)
);

A2O1A1Ixp33_ASAP7_75t_L g14970 ( 
.A1(n_12913),
.A2(n_10154),
.B(n_10155),
.C(n_10132),
.Y(n_14970)
);

AND2x2_ASAP7_75t_L g14971 ( 
.A(n_13810),
.B(n_13812),
.Y(n_14971)
);

AOI22xp5_ASAP7_75t_L g14972 ( 
.A1(n_13818),
.A2(n_13820),
.B1(n_13681),
.B2(n_13686),
.Y(n_14972)
);

OAI22xp5_ASAP7_75t_L g14973 ( 
.A1(n_13626),
.A2(n_9044),
.B1(n_9068),
.B2(n_9035),
.Y(n_14973)
);

OAI21x1_ASAP7_75t_L g14974 ( 
.A1(n_13989),
.A2(n_12828),
.B(n_11689),
.Y(n_14974)
);

AO21x2_ASAP7_75t_L g14975 ( 
.A1(n_13185),
.A2(n_13187),
.B(n_13186),
.Y(n_14975)
);

AND2x2_ASAP7_75t_L g14976 ( 
.A(n_13391),
.B(n_10829),
.Y(n_14976)
);

AND2x2_ASAP7_75t_L g14977 ( 
.A(n_13689),
.B(n_10829),
.Y(n_14977)
);

OR2x6_ASAP7_75t_L g14978 ( 
.A(n_13332),
.B(n_9005),
.Y(n_14978)
);

OAI21xp5_ASAP7_75t_L g14979 ( 
.A1(n_12933),
.A2(n_10873),
.B(n_10872),
.Y(n_14979)
);

AND2x2_ASAP7_75t_L g14980 ( 
.A(n_13704),
.B(n_10829),
.Y(n_14980)
);

AOI21xp5_ASAP7_75t_L g14981 ( 
.A1(n_13514),
.A2(n_10760),
.B(n_10835),
.Y(n_14981)
);

INVx3_ASAP7_75t_L g14982 ( 
.A(n_13110),
.Y(n_14982)
);

NAND2xp5_ASAP7_75t_L g14983 ( 
.A(n_13705),
.B(n_9523),
.Y(n_14983)
);

OR2x6_ASAP7_75t_L g14984 ( 
.A(n_13340),
.B(n_9005),
.Y(n_14984)
);

AOI22xp5_ASAP7_75t_L g14985 ( 
.A1(n_13713),
.A2(n_10438),
.B1(n_10345),
.B2(n_11007),
.Y(n_14985)
);

A2O1A1Ixp33_ASAP7_75t_L g14986 ( 
.A1(n_12963),
.A2(n_10154),
.B(n_10155),
.C(n_10132),
.Y(n_14986)
);

AND2x2_ASAP7_75t_L g14987 ( 
.A(n_13654),
.B(n_10833),
.Y(n_14987)
);

OR2x6_ASAP7_75t_L g14988 ( 
.A(n_13341),
.B(n_9005),
.Y(n_14988)
);

OAI22xp5_ASAP7_75t_L g14989 ( 
.A1(n_13357),
.A2(n_9086),
.B1(n_9090),
.B2(n_9068),
.Y(n_14989)
);

BUFx2_ASAP7_75t_L g14990 ( 
.A(n_13714),
.Y(n_14990)
);

INVx1_ASAP7_75t_L g14991 ( 
.A(n_13173),
.Y(n_14991)
);

AND2x2_ASAP7_75t_L g14992 ( 
.A(n_13675),
.B(n_10833),
.Y(n_14992)
);

OR2x2_ASAP7_75t_L g14993 ( 
.A(n_13679),
.B(n_10217),
.Y(n_14993)
);

AND2x6_ASAP7_75t_L g14994 ( 
.A(n_13343),
.B(n_10986),
.Y(n_14994)
);

OAI221xp5_ASAP7_75t_L g14995 ( 
.A1(n_13281),
.A2(n_10345),
.B1(n_13298),
.B2(n_13297),
.C(n_10831),
.Y(n_14995)
);

BUFx3_ASAP7_75t_L g14996 ( 
.A(n_13346),
.Y(n_14996)
);

CKINVDCx5p33_ASAP7_75t_R g14997 ( 
.A(n_13347),
.Y(n_14997)
);

AO22x2_ASAP7_75t_L g14998 ( 
.A1(n_13348),
.A2(n_11614),
.B1(n_11578),
.B2(n_11303),
.Y(n_14998)
);

NAND2xp5_ASAP7_75t_L g14999 ( 
.A(n_13176),
.B(n_9523),
.Y(n_14999)
);

OR2x2_ASAP7_75t_L g15000 ( 
.A(n_13357),
.B(n_10217),
.Y(n_15000)
);

AND2x2_ASAP7_75t_L g15001 ( 
.A(n_13398),
.B(n_10833),
.Y(n_15001)
);

O2A1O1Ixp33_ASAP7_75t_SL g15002 ( 
.A1(n_13310),
.A2(n_11303),
.B(n_11261),
.C(n_10307),
.Y(n_15002)
);

INVx2_ASAP7_75t_L g15003 ( 
.A(n_14072),
.Y(n_15003)
);

INVx2_ASAP7_75t_L g15004 ( 
.A(n_14249),
.Y(n_15004)
);

BUFx12f_ASAP7_75t_L g15005 ( 
.A(n_13996),
.Y(n_15005)
);

OR2x2_ASAP7_75t_L g15006 ( 
.A(n_14079),
.B(n_13900),
.Y(n_15006)
);

NAND2x1_ASAP7_75t_L g15007 ( 
.A(n_14481),
.B(n_13353),
.Y(n_15007)
);

NOR2xp33_ASAP7_75t_L g15008 ( 
.A(n_14032),
.B(n_13415),
.Y(n_15008)
);

OR2x2_ASAP7_75t_L g15009 ( 
.A(n_14020),
.B(n_13900),
.Y(n_15009)
);

AND2x2_ASAP7_75t_L g15010 ( 
.A(n_14039),
.B(n_13416),
.Y(n_15010)
);

INVx2_ASAP7_75t_L g15011 ( 
.A(n_14776),
.Y(n_15011)
);

AND2x2_ASAP7_75t_L g15012 ( 
.A(n_14364),
.B(n_14194),
.Y(n_15012)
);

INVx3_ASAP7_75t_L g15013 ( 
.A(n_14502),
.Y(n_15013)
);

AND2x2_ASAP7_75t_L g15014 ( 
.A(n_14022),
.B(n_13419),
.Y(n_15014)
);

INVx1_ASAP7_75t_L g15015 ( 
.A(n_14181),
.Y(n_15015)
);

OR2x2_ASAP7_75t_L g15016 ( 
.A(n_14012),
.B(n_13906),
.Y(n_15016)
);

AND2x2_ASAP7_75t_L g15017 ( 
.A(n_14036),
.B(n_13421),
.Y(n_15017)
);

HB1xp67_ASAP7_75t_L g15018 ( 
.A(n_14374),
.Y(n_15018)
);

INVx1_ASAP7_75t_L g15019 ( 
.A(n_14246),
.Y(n_15019)
);

INVx2_ASAP7_75t_L g15020 ( 
.A(n_14776),
.Y(n_15020)
);

HB1xp67_ASAP7_75t_L g15021 ( 
.A(n_14113),
.Y(n_15021)
);

INVx1_ASAP7_75t_L g15022 ( 
.A(n_14941),
.Y(n_15022)
);

AND2x4_ASAP7_75t_SL g15023 ( 
.A(n_14108),
.B(n_14068),
.Y(n_15023)
);

OR2x2_ASAP7_75t_L g15024 ( 
.A(n_14088),
.B(n_13906),
.Y(n_15024)
);

INVx1_ASAP7_75t_L g15025 ( 
.A(n_14948),
.Y(n_15025)
);

INVx2_ASAP7_75t_L g15026 ( 
.A(n_14776),
.Y(n_15026)
);

OAI22xp5_ASAP7_75t_L g15027 ( 
.A1(n_14017),
.A2(n_13572),
.B1(n_13554),
.B2(n_9872),
.Y(n_15027)
);

BUFx2_ASAP7_75t_L g15028 ( 
.A(n_14975),
.Y(n_15028)
);

INVx2_ASAP7_75t_L g15029 ( 
.A(n_14026),
.Y(n_15029)
);

AND2x2_ASAP7_75t_L g15030 ( 
.A(n_14031),
.B(n_13424),
.Y(n_15030)
);

INVx2_ASAP7_75t_L g15031 ( 
.A(n_14026),
.Y(n_15031)
);

AND2x2_ASAP7_75t_L g15032 ( 
.A(n_14134),
.B(n_14179),
.Y(n_15032)
);

AND2x4_ASAP7_75t_L g15033 ( 
.A(n_14492),
.B(n_13371),
.Y(n_15033)
);

INVx1_ASAP7_75t_L g15034 ( 
.A(n_14950),
.Y(n_15034)
);

NAND2xp5_ASAP7_75t_L g15035 ( 
.A(n_14267),
.B(n_13376),
.Y(n_15035)
);

AND2x2_ASAP7_75t_L g15036 ( 
.A(n_14179),
.B(n_13425),
.Y(n_15036)
);

INVx2_ASAP7_75t_L g15037 ( 
.A(n_14033),
.Y(n_15037)
);

INVx1_ASAP7_75t_L g15038 ( 
.A(n_14129),
.Y(n_15038)
);

HB1xp67_ASAP7_75t_L g15039 ( 
.A(n_14400),
.Y(n_15039)
);

INVxp67_ASAP7_75t_SL g15040 ( 
.A(n_14541),
.Y(n_15040)
);

AND2x2_ASAP7_75t_L g15041 ( 
.A(n_14202),
.B(n_13432),
.Y(n_15041)
);

INVx2_ASAP7_75t_L g15042 ( 
.A(n_14033),
.Y(n_15042)
);

AO21x2_ASAP7_75t_L g15043 ( 
.A1(n_14604),
.A2(n_13186),
.B(n_13185),
.Y(n_15043)
);

AND2x2_ASAP7_75t_L g15044 ( 
.A(n_14119),
.B(n_13434),
.Y(n_15044)
);

INVx2_ASAP7_75t_L g15045 ( 
.A(n_14146),
.Y(n_15045)
);

AND2x4_ASAP7_75t_L g15046 ( 
.A(n_14740),
.B(n_13381),
.Y(n_15046)
);

OAI221xp5_ASAP7_75t_L g15047 ( 
.A1(n_14002),
.A2(n_10831),
.B1(n_10893),
.B2(n_10892),
.C(n_10846),
.Y(n_15047)
);

INVx2_ASAP7_75t_L g15048 ( 
.A(n_14146),
.Y(n_15048)
);

OA21x2_ASAP7_75t_L g15049 ( 
.A1(n_14207),
.A2(n_13325),
.B(n_13310),
.Y(n_15049)
);

NAND2xp5_ASAP7_75t_L g15050 ( 
.A(n_14077),
.B(n_13386),
.Y(n_15050)
);

INVx2_ASAP7_75t_L g15051 ( 
.A(n_14345),
.Y(n_15051)
);

INVx4_ASAP7_75t_SL g15052 ( 
.A(n_14082),
.Y(n_15052)
);

AOI22xp33_ASAP7_75t_SL g15053 ( 
.A1(n_14038),
.A2(n_9872),
.B1(n_9892),
.B2(n_9838),
.Y(n_15053)
);

AND2x4_ASAP7_75t_L g15054 ( 
.A(n_14756),
.B(n_13439),
.Y(n_15054)
);

INVx1_ASAP7_75t_L g15055 ( 
.A(n_14420),
.Y(n_15055)
);

OA21x2_ASAP7_75t_L g15056 ( 
.A1(n_14207),
.A2(n_13330),
.B(n_13325),
.Y(n_15056)
);

INVx2_ASAP7_75t_L g15057 ( 
.A(n_14345),
.Y(n_15057)
);

INVx2_ASAP7_75t_L g15058 ( 
.A(n_14304),
.Y(n_15058)
);

INVx2_ASAP7_75t_SL g15059 ( 
.A(n_14431),
.Y(n_15059)
);

INVx1_ASAP7_75t_L g15060 ( 
.A(n_14473),
.Y(n_15060)
);

INVx1_ASAP7_75t_L g15061 ( 
.A(n_14477),
.Y(n_15061)
);

INVx2_ASAP7_75t_L g15062 ( 
.A(n_14119),
.Y(n_15062)
);

INVx2_ASAP7_75t_L g15063 ( 
.A(n_14303),
.Y(n_15063)
);

INVx1_ASAP7_75t_L g15064 ( 
.A(n_14557),
.Y(n_15064)
);

INVx1_ASAP7_75t_L g15065 ( 
.A(n_14564),
.Y(n_15065)
);

AND2x4_ASAP7_75t_L g15066 ( 
.A(n_14049),
.B(n_14092),
.Y(n_15066)
);

AND2x4_ASAP7_75t_L g15067 ( 
.A(n_14035),
.B(n_14401),
.Y(n_15067)
);

INVx1_ASAP7_75t_L g15068 ( 
.A(n_14172),
.Y(n_15068)
);

AND2x4_ASAP7_75t_L g15069 ( 
.A(n_14006),
.B(n_13443),
.Y(n_15069)
);

INVx1_ASAP7_75t_L g15070 ( 
.A(n_14197),
.Y(n_15070)
);

HB1xp67_ASAP7_75t_L g15071 ( 
.A(n_14212),
.Y(n_15071)
);

INVxp67_ASAP7_75t_SL g15072 ( 
.A(n_14544),
.Y(n_15072)
);

OA21x2_ASAP7_75t_L g15073 ( 
.A1(n_14260),
.A2(n_14838),
.B(n_14227),
.Y(n_15073)
);

INVx1_ASAP7_75t_L g15074 ( 
.A(n_14226),
.Y(n_15074)
);

AND2x2_ASAP7_75t_L g15075 ( 
.A(n_14281),
.B(n_14423),
.Y(n_15075)
);

INVx1_ASAP7_75t_L g15076 ( 
.A(n_14235),
.Y(n_15076)
);

INVx1_ASAP7_75t_L g15077 ( 
.A(n_14243),
.Y(n_15077)
);

BUFx2_ASAP7_75t_L g15078 ( 
.A(n_14278),
.Y(n_15078)
);

AND2x2_ASAP7_75t_L g15079 ( 
.A(n_14281),
.B(n_13446),
.Y(n_15079)
);

OR2x2_ASAP7_75t_L g15080 ( 
.A(n_14101),
.B(n_13554),
.Y(n_15080)
);

INVx1_ASAP7_75t_L g15081 ( 
.A(n_14245),
.Y(n_15081)
);

AND2x2_ASAP7_75t_L g15082 ( 
.A(n_14063),
.B(n_14064),
.Y(n_15082)
);

INVx2_ASAP7_75t_L g15083 ( 
.A(n_14303),
.Y(n_15083)
);

AND2x2_ASAP7_75t_L g15084 ( 
.A(n_14107),
.B(n_13453),
.Y(n_15084)
);

AOI22xp33_ASAP7_75t_L g15085 ( 
.A1(n_14047),
.A2(n_10345),
.B1(n_10760),
.B2(n_13486),
.Y(n_15085)
);

INVx1_ASAP7_75t_L g15086 ( 
.A(n_14253),
.Y(n_15086)
);

OR2x2_ASAP7_75t_L g15087 ( 
.A(n_14110),
.B(n_13572),
.Y(n_15087)
);

INVx2_ASAP7_75t_L g15088 ( 
.A(n_14373),
.Y(n_15088)
);

AND2x4_ASAP7_75t_SL g15089 ( 
.A(n_14213),
.B(n_9608),
.Y(n_15089)
);

INVx1_ASAP7_75t_L g15090 ( 
.A(n_14263),
.Y(n_15090)
);

INVx2_ASAP7_75t_L g15091 ( 
.A(n_14407),
.Y(n_15091)
);

AND2x2_ASAP7_75t_SL g15092 ( 
.A(n_14147),
.B(n_13076),
.Y(n_15092)
);

INVx2_ASAP7_75t_L g15093 ( 
.A(n_14448),
.Y(n_15093)
);

NAND2xp5_ASAP7_75t_L g15094 ( 
.A(n_14331),
.B(n_13180),
.Y(n_15094)
);

INVx3_ASAP7_75t_L g15095 ( 
.A(n_14183),
.Y(n_15095)
);

AND2x4_ASAP7_75t_L g15096 ( 
.A(n_14391),
.B(n_13454),
.Y(n_15096)
);

NAND2xp5_ASAP7_75t_L g15097 ( 
.A(n_14251),
.B(n_13192),
.Y(n_15097)
);

AND2x2_ASAP7_75t_L g15098 ( 
.A(n_14111),
.B(n_13194),
.Y(n_15098)
);

INVx3_ASAP7_75t_L g15099 ( 
.A(n_14402),
.Y(n_15099)
);

INVx1_ASAP7_75t_L g15100 ( 
.A(n_14264),
.Y(n_15100)
);

INVx3_ASAP7_75t_L g15101 ( 
.A(n_14254),
.Y(n_15101)
);

NOR2xp33_ASAP7_75t_L g15102 ( 
.A(n_14008),
.B(n_10986),
.Y(n_15102)
);

INVx1_ASAP7_75t_L g15103 ( 
.A(n_14282),
.Y(n_15103)
);

AND2x2_ASAP7_75t_L g15104 ( 
.A(n_14231),
.B(n_13196),
.Y(n_15104)
);

INVx2_ASAP7_75t_L g15105 ( 
.A(n_14306),
.Y(n_15105)
);

NAND2xp5_ASAP7_75t_L g15106 ( 
.A(n_14132),
.B(n_13199),
.Y(n_15106)
);

NAND2xp5_ASAP7_75t_L g15107 ( 
.A(n_14149),
.B(n_13202),
.Y(n_15107)
);

NAND2xp5_ASAP7_75t_L g15108 ( 
.A(n_14176),
.B(n_13203),
.Y(n_15108)
);

OR2x2_ASAP7_75t_L g15109 ( 
.A(n_14045),
.B(n_12982),
.Y(n_15109)
);

NOR2x1_ASAP7_75t_SL g15110 ( 
.A(n_14154),
.B(n_13698),
.Y(n_15110)
);

AND2x2_ASAP7_75t_L g15111 ( 
.A(n_14233),
.B(n_14238),
.Y(n_15111)
);

OR2x2_ASAP7_75t_L g15112 ( 
.A(n_14084),
.B(n_13623),
.Y(n_15112)
);

INVx2_ASAP7_75t_L g15113 ( 
.A(n_14306),
.Y(n_15113)
);

AND2x2_ASAP7_75t_L g15114 ( 
.A(n_14159),
.B(n_13205),
.Y(n_15114)
);

AND2x4_ASAP7_75t_L g15115 ( 
.A(n_14018),
.B(n_13207),
.Y(n_15115)
);

INVx2_ASAP7_75t_L g15116 ( 
.A(n_14291),
.Y(n_15116)
);

INVx2_ASAP7_75t_L g15117 ( 
.A(n_14483),
.Y(n_15117)
);

AND2x2_ASAP7_75t_L g15118 ( 
.A(n_14160),
.B(n_13208),
.Y(n_15118)
);

INVx1_ASAP7_75t_L g15119 ( 
.A(n_14314),
.Y(n_15119)
);

AND2x2_ASAP7_75t_L g15120 ( 
.A(n_14164),
.B(n_14171),
.Y(n_15120)
);

AND2x2_ASAP7_75t_L g15121 ( 
.A(n_14485),
.B(n_13209),
.Y(n_15121)
);

HB1xp67_ASAP7_75t_L g15122 ( 
.A(n_14255),
.Y(n_15122)
);

AND2x2_ASAP7_75t_L g15123 ( 
.A(n_14007),
.B(n_14177),
.Y(n_15123)
);

HB1xp67_ASAP7_75t_L g15124 ( 
.A(n_14255),
.Y(n_15124)
);

INVx2_ASAP7_75t_L g15125 ( 
.A(n_14483),
.Y(n_15125)
);

INVx1_ASAP7_75t_L g15126 ( 
.A(n_14335),
.Y(n_15126)
);

INVx1_ASAP7_75t_L g15127 ( 
.A(n_14337),
.Y(n_15127)
);

OR2x2_ASAP7_75t_L g15128 ( 
.A(n_14819),
.B(n_13628),
.Y(n_15128)
);

AND2x2_ASAP7_75t_L g15129 ( 
.A(n_14778),
.B(n_13213),
.Y(n_15129)
);

AND2x2_ASAP7_75t_SL g15130 ( 
.A(n_14266),
.B(n_13076),
.Y(n_15130)
);

AND2x2_ASAP7_75t_L g15131 ( 
.A(n_14166),
.B(n_13214),
.Y(n_15131)
);

AND2x2_ASAP7_75t_L g15132 ( 
.A(n_13994),
.B(n_13216),
.Y(n_15132)
);

INVx1_ASAP7_75t_L g15133 ( 
.A(n_14343),
.Y(n_15133)
);

AND2x2_ASAP7_75t_L g15134 ( 
.A(n_14178),
.B(n_13217),
.Y(n_15134)
);

NAND2xp5_ASAP7_75t_L g15135 ( 
.A(n_14004),
.B(n_13220),
.Y(n_15135)
);

INVx1_ASAP7_75t_L g15136 ( 
.A(n_14348),
.Y(n_15136)
);

AND2x2_ASAP7_75t_L g15137 ( 
.A(n_14095),
.B(n_13229),
.Y(n_15137)
);

INVx6_ASAP7_75t_L g15138 ( 
.A(n_14713),
.Y(n_15138)
);

INVx1_ASAP7_75t_L g15139 ( 
.A(n_14013),
.Y(n_15139)
);

BUFx3_ASAP7_75t_L g15140 ( 
.A(n_14617),
.Y(n_15140)
);

OR2x2_ASAP7_75t_L g15141 ( 
.A(n_14866),
.B(n_13629),
.Y(n_15141)
);

AND2x4_ASAP7_75t_L g15142 ( 
.A(n_14097),
.B(n_13231),
.Y(n_15142)
);

NAND2xp5_ASAP7_75t_L g15143 ( 
.A(n_14015),
.B(n_13233),
.Y(n_15143)
);

NAND2xp5_ASAP7_75t_L g15144 ( 
.A(n_14027),
.B(n_13239),
.Y(n_15144)
);

INVx1_ASAP7_75t_L g15145 ( 
.A(n_14023),
.Y(n_15145)
);

NOR2xp33_ASAP7_75t_R g15146 ( 
.A(n_14366),
.B(n_10986),
.Y(n_15146)
);

NAND2xp5_ASAP7_75t_L g15147 ( 
.A(n_14028),
.B(n_13240),
.Y(n_15147)
);

INVx2_ASAP7_75t_L g15148 ( 
.A(n_14532),
.Y(n_15148)
);

INVx1_ASAP7_75t_L g15149 ( 
.A(n_14046),
.Y(n_15149)
);

INVx5_ASAP7_75t_L g15150 ( 
.A(n_14675),
.Y(n_15150)
);

HB1xp67_ASAP7_75t_L g15151 ( 
.A(n_14714),
.Y(n_15151)
);

BUFx3_ASAP7_75t_L g15152 ( 
.A(n_14519),
.Y(n_15152)
);

INVx2_ASAP7_75t_L g15153 ( 
.A(n_14532),
.Y(n_15153)
);

INVx1_ASAP7_75t_L g15154 ( 
.A(n_14048),
.Y(n_15154)
);

INVx2_ASAP7_75t_L g15155 ( 
.A(n_14580),
.Y(n_15155)
);

INVx2_ASAP7_75t_L g15156 ( 
.A(n_14607),
.Y(n_15156)
);

NAND2xp5_ASAP7_75t_L g15157 ( 
.A(n_14044),
.B(n_13241),
.Y(n_15157)
);

INVx2_ASAP7_75t_L g15158 ( 
.A(n_14456),
.Y(n_15158)
);

AND2x2_ASAP7_75t_L g15159 ( 
.A(n_14098),
.B(n_13247),
.Y(n_15159)
);

AND2x2_ASAP7_75t_L g15160 ( 
.A(n_14742),
.B(n_13248),
.Y(n_15160)
);

BUFx3_ASAP7_75t_L g15161 ( 
.A(n_14519),
.Y(n_15161)
);

BUFx3_ASAP7_75t_L g15162 ( 
.A(n_14519),
.Y(n_15162)
);

AND2x2_ASAP7_75t_L g15163 ( 
.A(n_14173),
.B(n_13257),
.Y(n_15163)
);

AND2x2_ASAP7_75t_L g15164 ( 
.A(n_14126),
.B(n_13262),
.Y(n_15164)
);

OR2x2_ASAP7_75t_L g15165 ( 
.A(n_14917),
.B(n_13633),
.Y(n_15165)
);

INVx1_ASAP7_75t_L g15166 ( 
.A(n_14062),
.Y(n_15166)
);

AND2x2_ASAP7_75t_L g15167 ( 
.A(n_14128),
.B(n_13263),
.Y(n_15167)
);

INVx2_ASAP7_75t_L g15168 ( 
.A(n_14753),
.Y(n_15168)
);

NOR2x1p5_ASAP7_75t_L g15169 ( 
.A(n_13995),
.B(n_10135),
.Y(n_15169)
);

BUFx3_ASAP7_75t_L g15170 ( 
.A(n_14094),
.Y(n_15170)
);

CKINVDCx5p33_ASAP7_75t_R g15171 ( 
.A(n_14310),
.Y(n_15171)
);

NAND2xp5_ASAP7_75t_L g15172 ( 
.A(n_14078),
.B(n_13264),
.Y(n_15172)
);

OR2x2_ASAP7_75t_L g15173 ( 
.A(n_14131),
.B(n_14144),
.Y(n_15173)
);

INVx2_ASAP7_75t_L g15174 ( 
.A(n_14886),
.Y(n_15174)
);

AND2x2_ASAP7_75t_L g15175 ( 
.A(n_14570),
.B(n_13266),
.Y(n_15175)
);

AND2x2_ASAP7_75t_L g15176 ( 
.A(n_14439),
.B(n_13270),
.Y(n_15176)
);

NOR2xp33_ASAP7_75t_L g15177 ( 
.A(n_14297),
.B(n_11144),
.Y(n_15177)
);

INVx1_ASAP7_75t_L g15178 ( 
.A(n_14066),
.Y(n_15178)
);

HB1xp67_ASAP7_75t_L g15179 ( 
.A(n_14661),
.Y(n_15179)
);

AND2x2_ASAP7_75t_L g15180 ( 
.A(n_14042),
.B(n_13275),
.Y(n_15180)
);

INVx2_ASAP7_75t_L g15181 ( 
.A(n_14106),
.Y(n_15181)
);

BUFx3_ASAP7_75t_L g15182 ( 
.A(n_14822),
.Y(n_15182)
);

NAND2xp5_ASAP7_75t_L g15183 ( 
.A(n_14186),
.B(n_13277),
.Y(n_15183)
);

AND2x2_ASAP7_75t_L g15184 ( 
.A(n_14058),
.B(n_13280),
.Y(n_15184)
);

INVx2_ASAP7_75t_L g15185 ( 
.A(n_14618),
.Y(n_15185)
);

INVx1_ASAP7_75t_L g15186 ( 
.A(n_14067),
.Y(n_15186)
);

NAND2xp5_ASAP7_75t_L g15187 ( 
.A(n_14225),
.B(n_13285),
.Y(n_15187)
);

INVx2_ASAP7_75t_SL g15188 ( 
.A(n_14651),
.Y(n_15188)
);

INVx2_ASAP7_75t_L g15189 ( 
.A(n_14632),
.Y(n_15189)
);

INVx2_ASAP7_75t_L g15190 ( 
.A(n_14130),
.Y(n_15190)
);

NAND2xp5_ASAP7_75t_L g15191 ( 
.A(n_14232),
.B(n_13286),
.Y(n_15191)
);

INVx1_ASAP7_75t_L g15192 ( 
.A(n_14074),
.Y(n_15192)
);

OR2x2_ASAP7_75t_SL g15193 ( 
.A(n_13991),
.B(n_13417),
.Y(n_15193)
);

INVx2_ASAP7_75t_L g15194 ( 
.A(n_14311),
.Y(n_15194)
);

OR2x2_ASAP7_75t_L g15195 ( 
.A(n_14354),
.B(n_13635),
.Y(n_15195)
);

HB1xp67_ASAP7_75t_L g15196 ( 
.A(n_14852),
.Y(n_15196)
);

OAI22xp33_ASAP7_75t_L g15197 ( 
.A1(n_14375),
.A2(n_9872),
.B1(n_9892),
.B2(n_9838),
.Y(n_15197)
);

INVx2_ASAP7_75t_L g15198 ( 
.A(n_14100),
.Y(n_15198)
);

AND2x2_ASAP7_75t_L g15199 ( 
.A(n_14059),
.B(n_13287),
.Y(n_15199)
);

AND2x2_ASAP7_75t_L g15200 ( 
.A(n_14025),
.B(n_13289),
.Y(n_15200)
);

INVx1_ASAP7_75t_L g15201 ( 
.A(n_14081),
.Y(n_15201)
);

INVx5_ASAP7_75t_L g15202 ( 
.A(n_14675),
.Y(n_15202)
);

INVx1_ASAP7_75t_L g15203 ( 
.A(n_14083),
.Y(n_15203)
);

INVx3_ASAP7_75t_L g15204 ( 
.A(n_14548),
.Y(n_15204)
);

AOI22xp33_ASAP7_75t_L g15205 ( 
.A1(n_14209),
.A2(n_13486),
.B1(n_11007),
.B2(n_9283),
.Y(n_15205)
);

BUFx6f_ASAP7_75t_L g15206 ( 
.A(n_14309),
.Y(n_15206)
);

HB1xp67_ASAP7_75t_L g15207 ( 
.A(n_14362),
.Y(n_15207)
);

INVx1_ASAP7_75t_L g15208 ( 
.A(n_14089),
.Y(n_15208)
);

HB1xp67_ASAP7_75t_L g15209 ( 
.A(n_14379),
.Y(n_15209)
);

INVx4_ASAP7_75t_L g15210 ( 
.A(n_14284),
.Y(n_15210)
);

INVx1_ASAP7_75t_L g15211 ( 
.A(n_14093),
.Y(n_15211)
);

OR2x2_ASAP7_75t_L g15212 ( 
.A(n_14157),
.B(n_13636),
.Y(n_15212)
);

BUFx2_ASAP7_75t_L g15213 ( 
.A(n_14278),
.Y(n_15213)
);

BUFx3_ASAP7_75t_L g15214 ( 
.A(n_14104),
.Y(n_15214)
);

NOR2x1_ASAP7_75t_SL g15215 ( 
.A(n_14154),
.B(n_13698),
.Y(n_15215)
);

AND2x2_ASAP7_75t_L g15216 ( 
.A(n_14040),
.B(n_13290),
.Y(n_15216)
);

INVx1_ASAP7_75t_L g15217 ( 
.A(n_14140),
.Y(n_15217)
);

AND2x4_ASAP7_75t_L g15218 ( 
.A(n_14514),
.B(n_13291),
.Y(n_15218)
);

AND2x2_ASAP7_75t_L g15219 ( 
.A(n_14041),
.B(n_14135),
.Y(n_15219)
);

INVx2_ASAP7_75t_L g15220 ( 
.A(n_14763),
.Y(n_15220)
);

OA21x2_ASAP7_75t_L g15221 ( 
.A1(n_14260),
.A2(n_13414),
.B(n_13330),
.Y(n_15221)
);

INVxp67_ASAP7_75t_L g15222 ( 
.A(n_14009),
.Y(n_15222)
);

HB1xp67_ASAP7_75t_L g15223 ( 
.A(n_14395),
.Y(n_15223)
);

INVx3_ASAP7_75t_SL g15224 ( 
.A(n_14284),
.Y(n_15224)
);

AND2x4_ASAP7_75t_L g15225 ( 
.A(n_14417),
.B(n_13292),
.Y(n_15225)
);

AND2x2_ASAP7_75t_L g15226 ( 
.A(n_14141),
.B(n_13295),
.Y(n_15226)
);

BUFx3_ASAP7_75t_L g15227 ( 
.A(n_14675),
.Y(n_15227)
);

INVx2_ASAP7_75t_L g15228 ( 
.A(n_14517),
.Y(n_15228)
);

INVx2_ASAP7_75t_L g15229 ( 
.A(n_14528),
.Y(n_15229)
);

OAI332xp33_ASAP7_75t_L g15230 ( 
.A1(n_14174),
.A2(n_13104),
.A3(n_13760),
.B1(n_13751),
.B2(n_13765),
.B3(n_13767),
.C1(n_13758),
.C2(n_13757),
.Y(n_15230)
);

BUFx3_ASAP7_75t_L g15231 ( 
.A(n_14125),
.Y(n_15231)
);

NAND2xp5_ASAP7_75t_L g15232 ( 
.A(n_14247),
.B(n_13300),
.Y(n_15232)
);

AO21x2_ASAP7_75t_L g15233 ( 
.A1(n_14222),
.A2(n_13195),
.B(n_13187),
.Y(n_15233)
);

INVx1_ASAP7_75t_L g15234 ( 
.A(n_14145),
.Y(n_15234)
);

NAND2xp5_ASAP7_75t_L g15235 ( 
.A(n_14295),
.B(n_13305),
.Y(n_15235)
);

AND2x2_ASAP7_75t_L g15236 ( 
.A(n_14412),
.B(n_13306),
.Y(n_15236)
);

INVx2_ASAP7_75t_L g15237 ( 
.A(n_14711),
.Y(n_15237)
);

INVx2_ASAP7_75t_L g15238 ( 
.A(n_14732),
.Y(n_15238)
);

AOI22xp33_ASAP7_75t_L g15239 ( 
.A1(n_13998),
.A2(n_9283),
.B1(n_13824),
.B2(n_10124),
.Y(n_15239)
);

INVx2_ASAP7_75t_L g15240 ( 
.A(n_14737),
.Y(n_15240)
);

AND2x2_ASAP7_75t_L g15241 ( 
.A(n_14087),
.B(n_13311),
.Y(n_15241)
);

INVx1_ASAP7_75t_L g15242 ( 
.A(n_14153),
.Y(n_15242)
);

AND2x2_ASAP7_75t_L g15243 ( 
.A(n_14091),
.B(n_13313),
.Y(n_15243)
);

OR2x2_ASAP7_75t_L g15244 ( 
.A(n_14112),
.B(n_14175),
.Y(n_15244)
);

INVx2_ASAP7_75t_L g15245 ( 
.A(n_14752),
.Y(n_15245)
);

AND2x2_ASAP7_75t_L g15246 ( 
.A(n_14003),
.B(n_13320),
.Y(n_15246)
);

NAND2xp5_ASAP7_75t_L g15247 ( 
.A(n_14057),
.B(n_13323),
.Y(n_15247)
);

INVx1_ASAP7_75t_L g15248 ( 
.A(n_14158),
.Y(n_15248)
);

AND2x2_ASAP7_75t_L g15249 ( 
.A(n_14499),
.B(n_13324),
.Y(n_15249)
);

AND2x2_ASAP7_75t_L g15250 ( 
.A(n_14815),
.B(n_13329),
.Y(n_15250)
);

NOR2x1_ASAP7_75t_L g15251 ( 
.A(n_14525),
.B(n_13896),
.Y(n_15251)
);

INVxp67_ASAP7_75t_L g15252 ( 
.A(n_14774),
.Y(n_15252)
);

INVx2_ASAP7_75t_L g15253 ( 
.A(n_14411),
.Y(n_15253)
);

AND2x4_ASAP7_75t_L g15254 ( 
.A(n_14612),
.B(n_13331),
.Y(n_15254)
);

AND2x2_ASAP7_75t_L g15255 ( 
.A(n_14185),
.B(n_13333),
.Y(n_15255)
);

INVx1_ASAP7_75t_L g15256 ( 
.A(n_14605),
.Y(n_15256)
);

BUFx3_ASAP7_75t_L g15257 ( 
.A(n_14630),
.Y(n_15257)
);

HB1xp67_ASAP7_75t_L g15258 ( 
.A(n_14965),
.Y(n_15258)
);

INVx1_ASAP7_75t_L g15259 ( 
.A(n_14854),
.Y(n_15259)
);

INVx1_ASAP7_75t_L g15260 ( 
.A(n_14888),
.Y(n_15260)
);

INVx3_ASAP7_75t_L g15261 ( 
.A(n_14052),
.Y(n_15261)
);

NAND2xp5_ASAP7_75t_L g15262 ( 
.A(n_14593),
.B(n_13338),
.Y(n_15262)
);

INVx1_ASAP7_75t_L g15263 ( 
.A(n_14406),
.Y(n_15263)
);

AND2x2_ASAP7_75t_L g15264 ( 
.A(n_14188),
.B(n_14369),
.Y(n_15264)
);

INVx2_ASAP7_75t_SL g15265 ( 
.A(n_14938),
.Y(n_15265)
);

INVx3_ASAP7_75t_L g15266 ( 
.A(n_14229),
.Y(n_15266)
);

INVxp67_ASAP7_75t_L g15267 ( 
.A(n_14530),
.Y(n_15267)
);

AOI22xp33_ASAP7_75t_L g15268 ( 
.A1(n_14117),
.A2(n_9283),
.B1(n_13824),
.B2(n_10124),
.Y(n_15268)
);

INVx1_ASAP7_75t_L g15269 ( 
.A(n_14782),
.Y(n_15269)
);

AND2x4_ASAP7_75t_L g15270 ( 
.A(n_14777),
.B(n_13344),
.Y(n_15270)
);

INVx2_ASAP7_75t_L g15271 ( 
.A(n_14422),
.Y(n_15271)
);

AND2x2_ASAP7_75t_L g15272 ( 
.A(n_14076),
.B(n_13345),
.Y(n_15272)
);

OAI22xp5_ASAP7_75t_L g15273 ( 
.A1(n_14024),
.A2(n_14029),
.B1(n_14103),
.B2(n_14118),
.Y(n_15273)
);

INVx1_ASAP7_75t_L g15274 ( 
.A(n_14782),
.Y(n_15274)
);

OR2x2_ASAP7_75t_L g15275 ( 
.A(n_14162),
.B(n_13351),
.Y(n_15275)
);

INVx1_ASAP7_75t_L g15276 ( 
.A(n_14408),
.Y(n_15276)
);

AND2x2_ASAP7_75t_L g15277 ( 
.A(n_14221),
.B(n_13359),
.Y(n_15277)
);

NAND2xp5_ASAP7_75t_L g15278 ( 
.A(n_14721),
.B(n_13369),
.Y(n_15278)
);

NOR2xp33_ASAP7_75t_L g15279 ( 
.A(n_14500),
.B(n_11144),
.Y(n_15279)
);

INVx1_ASAP7_75t_L g15280 ( 
.A(n_14416),
.Y(n_15280)
);

AOI22xp33_ASAP7_75t_L g15281 ( 
.A1(n_14211),
.A2(n_9283),
.B1(n_10124),
.B2(n_9590),
.Y(n_15281)
);

INVx2_ASAP7_75t_L g15282 ( 
.A(n_14438),
.Y(n_15282)
);

OAI211xp5_ASAP7_75t_L g15283 ( 
.A1(n_14250),
.A2(n_13079),
.B(n_13336),
.C(n_13326),
.Y(n_15283)
);

HB1xp67_ASAP7_75t_L g15284 ( 
.A(n_14965),
.Y(n_15284)
);

INVx2_ASAP7_75t_L g15285 ( 
.A(n_14440),
.Y(n_15285)
);

INVx1_ASAP7_75t_L g15286 ( 
.A(n_14462),
.Y(n_15286)
);

HB1xp67_ASAP7_75t_L g15287 ( 
.A(n_14990),
.Y(n_15287)
);

INVx3_ASAP7_75t_L g15288 ( 
.A(n_14230),
.Y(n_15288)
);

AND2x4_ASAP7_75t_L g15289 ( 
.A(n_14494),
.B(n_13374),
.Y(n_15289)
);

OR2x2_ASAP7_75t_L g15290 ( 
.A(n_14220),
.B(n_14455),
.Y(n_15290)
);

INVx1_ASAP7_75t_L g15291 ( 
.A(n_14472),
.Y(n_15291)
);

AND2x2_ASAP7_75t_L g15292 ( 
.A(n_14228),
.B(n_13375),
.Y(n_15292)
);

INVx2_ASAP7_75t_L g15293 ( 
.A(n_14527),
.Y(n_15293)
);

INVx1_ASAP7_75t_L g15294 ( 
.A(n_14488),
.Y(n_15294)
);

AND2x2_ASAP7_75t_L g15295 ( 
.A(n_14204),
.B(n_13394),
.Y(n_15295)
);

INVx2_ASAP7_75t_L g15296 ( 
.A(n_14571),
.Y(n_15296)
);

AOI22xp33_ASAP7_75t_SL g15297 ( 
.A1(n_14122),
.A2(n_9872),
.B1(n_9892),
.B2(n_9838),
.Y(n_15297)
);

AND2x4_ASAP7_75t_L g15298 ( 
.A(n_14576),
.B(n_13395),
.Y(n_15298)
);

INVx1_ASAP7_75t_L g15299 ( 
.A(n_14503),
.Y(n_15299)
);

HB1xp67_ASAP7_75t_L g15300 ( 
.A(n_14990),
.Y(n_15300)
);

HB1xp67_ASAP7_75t_L g15301 ( 
.A(n_14424),
.Y(n_15301)
);

BUFx3_ASAP7_75t_L g15302 ( 
.A(n_14706),
.Y(n_15302)
);

INVx2_ASAP7_75t_L g15303 ( 
.A(n_14594),
.Y(n_15303)
);

BUFx2_ASAP7_75t_L g15304 ( 
.A(n_14871),
.Y(n_15304)
);

AND2x2_ASAP7_75t_L g15305 ( 
.A(n_14371),
.B(n_13399),
.Y(n_15305)
);

INVx1_ASAP7_75t_SL g15306 ( 
.A(n_14071),
.Y(n_15306)
);

AND2x2_ASAP7_75t_L g15307 ( 
.A(n_14377),
.B(n_13403),
.Y(n_15307)
);

INVx2_ASAP7_75t_L g15308 ( 
.A(n_14628),
.Y(n_15308)
);

BUFx2_ASAP7_75t_L g15309 ( 
.A(n_14525),
.Y(n_15309)
);

INVxp67_ASAP7_75t_SL g15310 ( 
.A(n_14644),
.Y(n_15310)
);

INVx2_ASAP7_75t_L g15311 ( 
.A(n_14657),
.Y(n_15311)
);

INVx2_ASAP7_75t_L g15312 ( 
.A(n_14755),
.Y(n_15312)
);

AOI221xp5_ASAP7_75t_L g15313 ( 
.A1(n_13992),
.A2(n_13896),
.B1(n_11603),
.B2(n_11627),
.C(n_10762),
.Y(n_15313)
);

AND2x2_ASAP7_75t_L g15314 ( 
.A(n_14403),
.B(n_13411),
.Y(n_15314)
);

AND2x2_ASAP7_75t_L g15315 ( 
.A(n_14409),
.B(n_13412),
.Y(n_15315)
);

OR2x2_ASAP7_75t_L g15316 ( 
.A(n_14478),
.B(n_13423),
.Y(n_15316)
);

INVx1_ASAP7_75t_L g15317 ( 
.A(n_14509),
.Y(n_15317)
);

AND2x2_ASAP7_75t_L g15318 ( 
.A(n_14139),
.B(n_13426),
.Y(n_15318)
);

AND2x2_ASAP7_75t_L g15319 ( 
.A(n_14136),
.B(n_14200),
.Y(n_15319)
);

BUFx2_ASAP7_75t_L g15320 ( 
.A(n_14638),
.Y(n_15320)
);

INVx1_ASAP7_75t_L g15321 ( 
.A(n_14526),
.Y(n_15321)
);

OR2x2_ASAP7_75t_L g15322 ( 
.A(n_14486),
.B(n_13428),
.Y(n_15322)
);

OAI21x1_ASAP7_75t_L g15323 ( 
.A1(n_14747),
.A2(n_13779),
.B(n_13771),
.Y(n_15323)
);

AND2x2_ASAP7_75t_L g15324 ( 
.A(n_14326),
.B(n_14328),
.Y(n_15324)
);

AND2x4_ASAP7_75t_L g15325 ( 
.A(n_14669),
.B(n_13429),
.Y(n_15325)
);

NOR2xp33_ASAP7_75t_L g15326 ( 
.A(n_14109),
.B(n_11144),
.Y(n_15326)
);

INVx1_ASAP7_75t_L g15327 ( 
.A(n_14542),
.Y(n_15327)
);

AND2x2_ASAP7_75t_L g15328 ( 
.A(n_14332),
.B(n_13431),
.Y(n_15328)
);

INVx1_ASAP7_75t_L g15329 ( 
.A(n_14545),
.Y(n_15329)
);

INVx1_ASAP7_75t_L g15330 ( 
.A(n_14547),
.Y(n_15330)
);

AND2x4_ASAP7_75t_L g15331 ( 
.A(n_14696),
.B(n_13437),
.Y(n_15331)
);

INVx1_ASAP7_75t_L g15332 ( 
.A(n_14549),
.Y(n_15332)
);

INVx3_ASAP7_75t_L g15333 ( 
.A(n_14234),
.Y(n_15333)
);

AO31x2_ASAP7_75t_L g15334 ( 
.A1(n_14638),
.A2(n_13444),
.A3(n_13461),
.B(n_13440),
.Y(n_15334)
);

INVx1_ASAP7_75t_L g15335 ( 
.A(n_14559),
.Y(n_15335)
);

AND2x2_ASAP7_75t_L g15336 ( 
.A(n_14336),
.B(n_13473),
.Y(n_15336)
);

AND2x2_ASAP7_75t_L g15337 ( 
.A(n_14363),
.B(n_13475),
.Y(n_15337)
);

INVx1_ASAP7_75t_SL g15338 ( 
.A(n_14070),
.Y(n_15338)
);

AND2x2_ASAP7_75t_L g15339 ( 
.A(n_13997),
.B(n_13477),
.Y(n_15339)
);

OAI21xp5_ASAP7_75t_SL g15340 ( 
.A1(n_14152),
.A2(n_10846),
.B(n_10831),
.Y(n_15340)
);

BUFx2_ASAP7_75t_L g15341 ( 
.A(n_14673),
.Y(n_15341)
);

INVx1_ASAP7_75t_L g15342 ( 
.A(n_14566),
.Y(n_15342)
);

INVx2_ASAP7_75t_SL g15343 ( 
.A(n_14723),
.Y(n_15343)
);

BUFx6f_ASAP7_75t_L g15344 ( 
.A(n_14321),
.Y(n_15344)
);

INVx1_ASAP7_75t_L g15345 ( 
.A(n_14636),
.Y(n_15345)
);

CKINVDCx5p33_ASAP7_75t_R g15346 ( 
.A(n_14321),
.Y(n_15346)
);

AND2x2_ASAP7_75t_L g15347 ( 
.A(n_14050),
.B(n_13478),
.Y(n_15347)
);

INVx1_ASAP7_75t_L g15348 ( 
.A(n_14637),
.Y(n_15348)
);

AND2x2_ASAP7_75t_L g15349 ( 
.A(n_14708),
.B(n_13491),
.Y(n_15349)
);

AND2x2_ASAP7_75t_L g15350 ( 
.A(n_14283),
.B(n_13493),
.Y(n_15350)
);

AND2x2_ASAP7_75t_L g15351 ( 
.A(n_14299),
.B(n_13497),
.Y(n_15351)
);

INVx4_ASAP7_75t_L g15352 ( 
.A(n_14599),
.Y(n_15352)
);

BUFx2_ASAP7_75t_L g15353 ( 
.A(n_14673),
.Y(n_15353)
);

BUFx2_ASAP7_75t_L g15354 ( 
.A(n_14069),
.Y(n_15354)
);

OR2x2_ASAP7_75t_L g15355 ( 
.A(n_14201),
.B(n_13498),
.Y(n_15355)
);

AND2x2_ASAP7_75t_L g15356 ( 
.A(n_14317),
.B(n_13500),
.Y(n_15356)
);

INVx1_ASAP7_75t_L g15357 ( 
.A(n_14654),
.Y(n_15357)
);

HB1xp67_ASAP7_75t_L g15358 ( 
.A(n_14725),
.Y(n_15358)
);

BUFx12f_ASAP7_75t_L g15359 ( 
.A(n_14555),
.Y(n_15359)
);

INVx2_ASAP7_75t_L g15360 ( 
.A(n_14758),
.Y(n_15360)
);

AND2x2_ASAP7_75t_L g15361 ( 
.A(n_14116),
.B(n_13501),
.Y(n_15361)
);

AND2x2_ASAP7_75t_L g15362 ( 
.A(n_14156),
.B(n_13504),
.Y(n_15362)
);

HB1xp67_ASAP7_75t_L g15363 ( 
.A(n_14761),
.Y(n_15363)
);

NAND2xp5_ASAP7_75t_L g15364 ( 
.A(n_14193),
.B(n_13507),
.Y(n_15364)
);

INVx4_ASAP7_75t_L g15365 ( 
.A(n_14457),
.Y(n_15365)
);

INVxp67_ASAP7_75t_L g15366 ( 
.A(n_14010),
.Y(n_15366)
);

INVx1_ASAP7_75t_L g15367 ( 
.A(n_14666),
.Y(n_15367)
);

OR2x2_ASAP7_75t_L g15368 ( 
.A(n_14203),
.B(n_13509),
.Y(n_15368)
);

AO21x2_ASAP7_75t_L g15369 ( 
.A1(n_14214),
.A2(n_13230),
.B(n_13195),
.Y(n_15369)
);

INVx2_ASAP7_75t_L g15370 ( 
.A(n_14765),
.Y(n_15370)
);

INVx2_ASAP7_75t_L g15371 ( 
.A(n_14735),
.Y(n_15371)
);

BUFx6f_ASAP7_75t_L g15372 ( 
.A(n_14700),
.Y(n_15372)
);

INVx2_ASAP7_75t_L g15373 ( 
.A(n_14738),
.Y(n_15373)
);

AND2x4_ASAP7_75t_L g15374 ( 
.A(n_14114),
.B(n_13512),
.Y(n_15374)
);

HB1xp67_ASAP7_75t_L g15375 ( 
.A(n_14956),
.Y(n_15375)
);

INVx2_ASAP7_75t_L g15376 ( 
.A(n_14748),
.Y(n_15376)
);

INVx1_ASAP7_75t_L g15377 ( 
.A(n_14897),
.Y(n_15377)
);

BUFx6f_ASAP7_75t_L g15378 ( 
.A(n_14700),
.Y(n_15378)
);

HB1xp67_ASAP7_75t_L g15379 ( 
.A(n_14958),
.Y(n_15379)
);

INVx2_ASAP7_75t_L g15380 ( 
.A(n_14769),
.Y(n_15380)
);

INVx1_ASAP7_75t_L g15381 ( 
.A(n_14933),
.Y(n_15381)
);

AOI21xp5_ASAP7_75t_SL g15382 ( 
.A1(n_14127),
.A2(n_13079),
.B(n_13326),
.Y(n_15382)
);

AND2x2_ASAP7_75t_L g15383 ( 
.A(n_14239),
.B(n_14248),
.Y(n_15383)
);

INVx1_ASAP7_75t_L g15384 ( 
.A(n_14954),
.Y(n_15384)
);

INVx2_ASAP7_75t_L g15385 ( 
.A(n_14773),
.Y(n_15385)
);

INVx2_ASAP7_75t_L g15386 ( 
.A(n_14910),
.Y(n_15386)
);

AOI22xp33_ASAP7_75t_L g15387 ( 
.A1(n_13999),
.A2(n_9283),
.B1(n_10124),
.B2(n_9590),
.Y(n_15387)
);

INVx1_ASAP7_75t_L g15388 ( 
.A(n_14961),
.Y(n_15388)
);

INVx1_ASAP7_75t_L g15389 ( 
.A(n_14966),
.Y(n_15389)
);

INVxp67_ASAP7_75t_SL g15390 ( 
.A(n_14759),
.Y(n_15390)
);

AO21x2_ASAP7_75t_L g15391 ( 
.A1(n_14001),
.A2(n_13236),
.B(n_13230),
.Y(n_15391)
);

INVx1_ASAP7_75t_L g15392 ( 
.A(n_14991),
.Y(n_15392)
);

AND2x2_ASAP7_75t_L g15393 ( 
.A(n_14271),
.B(n_13517),
.Y(n_15393)
);

INVx2_ASAP7_75t_L g15394 ( 
.A(n_14578),
.Y(n_15394)
);

BUFx3_ASAP7_75t_L g15395 ( 
.A(n_14807),
.Y(n_15395)
);

BUFx3_ASAP7_75t_L g15396 ( 
.A(n_14836),
.Y(n_15396)
);

INVx1_ASAP7_75t_L g15397 ( 
.A(n_14667),
.Y(n_15397)
);

AO31x2_ASAP7_75t_L g15398 ( 
.A1(n_14664),
.A2(n_13521),
.A3(n_13536),
.B(n_13531),
.Y(n_15398)
);

OR2x2_ASAP7_75t_L g15399 ( 
.A(n_14904),
.B(n_13548),
.Y(n_15399)
);

NAND2xp5_ASAP7_75t_L g15400 ( 
.A(n_14734),
.B(n_13550),
.Y(n_15400)
);

BUFx2_ASAP7_75t_L g15401 ( 
.A(n_14772),
.Y(n_15401)
);

AND2x4_ASAP7_75t_L g15402 ( 
.A(n_14619),
.B(n_13559),
.Y(n_15402)
);

AND2x2_ASAP7_75t_L g15403 ( 
.A(n_14279),
.B(n_13561),
.Y(n_15403)
);

INVx1_ASAP7_75t_SL g15404 ( 
.A(n_14697),
.Y(n_15404)
);

INVx1_ASAP7_75t_L g15405 ( 
.A(n_14687),
.Y(n_15405)
);

INVx1_ASAP7_75t_L g15406 ( 
.A(n_14720),
.Y(n_15406)
);

INVx2_ASAP7_75t_L g15407 ( 
.A(n_14588),
.Y(n_15407)
);

INVx1_ASAP7_75t_L g15408 ( 
.A(n_14736),
.Y(n_15408)
);

INVx2_ASAP7_75t_L g15409 ( 
.A(n_14606),
.Y(n_15409)
);

INVx2_ASAP7_75t_L g15410 ( 
.A(n_14608),
.Y(n_15410)
);

INVx1_ASAP7_75t_L g15411 ( 
.A(n_14744),
.Y(n_15411)
);

INVx3_ASAP7_75t_L g15412 ( 
.A(n_14252),
.Y(n_15412)
);

BUFx2_ASAP7_75t_L g15413 ( 
.A(n_14772),
.Y(n_15413)
);

INVxp67_ASAP7_75t_SL g15414 ( 
.A(n_14446),
.Y(n_15414)
);

INVx1_ASAP7_75t_L g15415 ( 
.A(n_14750),
.Y(n_15415)
);

INVx4_ASAP7_75t_L g15416 ( 
.A(n_14457),
.Y(n_15416)
);

AND2x4_ASAP7_75t_L g15417 ( 
.A(n_14581),
.B(n_13562),
.Y(n_15417)
);

AOI22xp33_ASAP7_75t_L g15418 ( 
.A1(n_14000),
.A2(n_9283),
.B1(n_10124),
.B2(n_9590),
.Y(n_15418)
);

NAND2xp5_ASAP7_75t_L g15419 ( 
.A(n_14899),
.B(n_13563),
.Y(n_15419)
);

INVx1_ASAP7_75t_L g15420 ( 
.A(n_14780),
.Y(n_15420)
);

NAND2xp5_ASAP7_75t_L g15421 ( 
.A(n_14726),
.B(n_13566),
.Y(n_15421)
);

AND2x2_ASAP7_75t_L g15422 ( 
.A(n_14280),
.B(n_13570),
.Y(n_15422)
);

INVx1_ASAP7_75t_L g15423 ( 
.A(n_14799),
.Y(n_15423)
);

NAND2xp5_ASAP7_75t_L g15424 ( 
.A(n_14922),
.B(n_13577),
.Y(n_15424)
);

OR2x2_ASAP7_75t_L g15425 ( 
.A(n_14394),
.B(n_14376),
.Y(n_15425)
);

AND2x2_ASAP7_75t_L g15426 ( 
.A(n_14722),
.B(n_13578),
.Y(n_15426)
);

OR2x6_ASAP7_75t_L g15427 ( 
.A(n_14484),
.B(n_9756),
.Y(n_15427)
);

INVx2_ASAP7_75t_L g15428 ( 
.A(n_14609),
.Y(n_15428)
);

INVx4_ASAP7_75t_L g15429 ( 
.A(n_14484),
.Y(n_15429)
);

INVx2_ASAP7_75t_L g15430 ( 
.A(n_14611),
.Y(n_15430)
);

NAND2xp5_ASAP7_75t_L g15431 ( 
.A(n_14859),
.B(n_13585),
.Y(n_15431)
);

AND2x2_ASAP7_75t_L g15432 ( 
.A(n_14120),
.B(n_14121),
.Y(n_15432)
);

NAND2xp5_ASAP7_75t_L g15433 ( 
.A(n_14902),
.B(n_13587),
.Y(n_15433)
);

INVx1_ASAP7_75t_L g15434 ( 
.A(n_14810),
.Y(n_15434)
);

AND2x2_ASAP7_75t_L g15435 ( 
.A(n_14123),
.B(n_13590),
.Y(n_15435)
);

INVx1_ASAP7_75t_L g15436 ( 
.A(n_14821),
.Y(n_15436)
);

BUFx2_ASAP7_75t_L g15437 ( 
.A(n_14085),
.Y(n_15437)
);

AND2x2_ASAP7_75t_L g15438 ( 
.A(n_14265),
.B(n_13591),
.Y(n_15438)
);

INVx2_ASAP7_75t_L g15439 ( 
.A(n_14639),
.Y(n_15439)
);

AND2x2_ASAP7_75t_L g15440 ( 
.A(n_14296),
.B(n_13593),
.Y(n_15440)
);

AND2x2_ASAP7_75t_L g15441 ( 
.A(n_14308),
.B(n_13595),
.Y(n_15441)
);

INVx2_ASAP7_75t_L g15442 ( 
.A(n_14138),
.Y(n_15442)
);

INVxp67_ASAP7_75t_SL g15443 ( 
.A(n_14898),
.Y(n_15443)
);

INVx2_ASAP7_75t_L g15444 ( 
.A(n_14187),
.Y(n_15444)
);

NOR2xp33_ASAP7_75t_L g15445 ( 
.A(n_14405),
.B(n_11144),
.Y(n_15445)
);

AND2x2_ASAP7_75t_L g15446 ( 
.A(n_14189),
.B(n_13597),
.Y(n_15446)
);

INVx1_ASAP7_75t_L g15447 ( 
.A(n_14827),
.Y(n_15447)
);

AND2x2_ASAP7_75t_L g15448 ( 
.A(n_14192),
.B(n_10833),
.Y(n_15448)
);

AND2x2_ASAP7_75t_L g15449 ( 
.A(n_14151),
.B(n_10833),
.Y(n_15449)
);

HB1xp67_ASAP7_75t_L g15450 ( 
.A(n_14620),
.Y(n_15450)
);

OAI22xp33_ASAP7_75t_L g15451 ( 
.A1(n_14090),
.A2(n_9872),
.B1(n_9892),
.B2(n_9838),
.Y(n_15451)
);

AND2x2_ASAP7_75t_L g15452 ( 
.A(n_14629),
.B(n_10838),
.Y(n_15452)
);

INVx1_ASAP7_75t_L g15453 ( 
.A(n_14837),
.Y(n_15453)
);

AND2x2_ASAP7_75t_L g15454 ( 
.A(n_14474),
.B(n_10838),
.Y(n_15454)
);

INVx2_ASAP7_75t_L g15455 ( 
.A(n_14206),
.Y(n_15455)
);

OR2x2_ASAP7_75t_L g15456 ( 
.A(n_14427),
.B(n_13673),
.Y(n_15456)
);

AND2x2_ASAP7_75t_L g15457 ( 
.A(n_14490),
.B(n_10838),
.Y(n_15457)
);

AOI22xp33_ASAP7_75t_L g15458 ( 
.A1(n_14150),
.A2(n_9283),
.B1(n_10124),
.B2(n_9590),
.Y(n_15458)
);

INVx1_ASAP7_75t_L g15459 ( 
.A(n_14843),
.Y(n_15459)
);

INVx2_ASAP7_75t_L g15460 ( 
.A(n_14210),
.Y(n_15460)
);

AND2x2_ASAP7_75t_L g15461 ( 
.A(n_14413),
.B(n_10838),
.Y(n_15461)
);

INVx2_ASAP7_75t_L g15462 ( 
.A(n_14218),
.Y(n_15462)
);

BUFx2_ASAP7_75t_L g15463 ( 
.A(n_14085),
.Y(n_15463)
);

OR2x2_ASAP7_75t_L g15464 ( 
.A(n_14921),
.B(n_13673),
.Y(n_15464)
);

INVx1_ASAP7_75t_L g15465 ( 
.A(n_14846),
.Y(n_15465)
);

INVx2_ASAP7_75t_L g15466 ( 
.A(n_14680),
.Y(n_15466)
);

AND2x2_ASAP7_75t_L g15467 ( 
.A(n_14425),
.B(n_10838),
.Y(n_15467)
);

OR2x2_ASAP7_75t_L g15468 ( 
.A(n_14923),
.B(n_13141),
.Y(n_15468)
);

BUFx6f_ASAP7_75t_L g15469 ( 
.A(n_14891),
.Y(n_15469)
);

NAND2xp5_ASAP7_75t_L g15470 ( 
.A(n_14865),
.B(n_13599),
.Y(n_15470)
);

OR2x6_ASAP7_75t_L g15471 ( 
.A(n_14389),
.B(n_9756),
.Y(n_15471)
);

INVx2_ASAP7_75t_L g15472 ( 
.A(n_14682),
.Y(n_15472)
);

BUFx2_ASAP7_75t_L g15473 ( 
.A(n_14298),
.Y(n_15473)
);

HB1xp67_ASAP7_75t_L g15474 ( 
.A(n_14620),
.Y(n_15474)
);

INVx2_ASAP7_75t_L g15475 ( 
.A(n_14690),
.Y(n_15475)
);

AND2x4_ASAP7_75t_L g15476 ( 
.A(n_14786),
.B(n_11357),
.Y(n_15476)
);

INVx4_ASAP7_75t_R g15477 ( 
.A(n_14692),
.Y(n_15477)
);

NAND2xp5_ASAP7_75t_L g15478 ( 
.A(n_14892),
.B(n_13600),
.Y(n_15478)
);

AND2x2_ASAP7_75t_L g15479 ( 
.A(n_14436),
.B(n_14461),
.Y(n_15479)
);

INVx2_ASAP7_75t_L g15480 ( 
.A(n_14691),
.Y(n_15480)
);

NOR2x1_ASAP7_75t_L g15481 ( 
.A(n_14198),
.B(n_13712),
.Y(n_15481)
);

INVx1_ASAP7_75t_L g15482 ( 
.A(n_14847),
.Y(n_15482)
);

AND2x2_ASAP7_75t_SL g15483 ( 
.A(n_14014),
.B(n_9792),
.Y(n_15483)
);

NOR2x1_ASAP7_75t_L g15484 ( 
.A(n_14011),
.B(n_13712),
.Y(n_15484)
);

NAND2xp5_ASAP7_75t_L g15485 ( 
.A(n_14997),
.B(n_13601),
.Y(n_15485)
);

INVx2_ASAP7_75t_L g15486 ( 
.A(n_14693),
.Y(n_15486)
);

HB1xp67_ASAP7_75t_L g15487 ( 
.A(n_14870),
.Y(n_15487)
);

BUFx3_ASAP7_75t_L g15488 ( 
.A(n_14994),
.Y(n_15488)
);

INVx2_ASAP7_75t_L g15489 ( 
.A(n_14710),
.Y(n_15489)
);

BUFx3_ASAP7_75t_L g15490 ( 
.A(n_14994),
.Y(n_15490)
);

INVx1_ASAP7_75t_L g15491 ( 
.A(n_14853),
.Y(n_15491)
);

INVx1_ASAP7_75t_L g15492 ( 
.A(n_14869),
.Y(n_15492)
);

INVx2_ASAP7_75t_L g15493 ( 
.A(n_14891),
.Y(n_15493)
);

AND2x2_ASAP7_75t_L g15494 ( 
.A(n_14634),
.B(n_14196),
.Y(n_15494)
);

AND2x2_ASAP7_75t_L g15495 ( 
.A(n_14572),
.B(n_10870),
.Y(n_15495)
);

INVxp67_ASAP7_75t_SL g15496 ( 
.A(n_14357),
.Y(n_15496)
);

HB1xp67_ASAP7_75t_L g15497 ( 
.A(n_14996),
.Y(n_15497)
);

OR2x2_ASAP7_75t_L g15498 ( 
.A(n_14963),
.B(n_13160),
.Y(n_15498)
);

OR2x2_ASAP7_75t_L g15499 ( 
.A(n_14982),
.B(n_12910),
.Y(n_15499)
);

NAND2xp5_ASAP7_75t_L g15500 ( 
.A(n_14294),
.B(n_13604),
.Y(n_15500)
);

OR2x2_ASAP7_75t_L g15501 ( 
.A(n_14447),
.B(n_13849),
.Y(n_15501)
);

INVx2_ASAP7_75t_L g15502 ( 
.A(n_14645),
.Y(n_15502)
);

AND2x2_ASAP7_75t_L g15503 ( 
.A(n_14575),
.B(n_10870),
.Y(n_15503)
);

INVx1_ASAP7_75t_L g15504 ( 
.A(n_14889),
.Y(n_15504)
);

INVx1_ASAP7_75t_L g15505 ( 
.A(n_14894),
.Y(n_15505)
);

OR2x2_ASAP7_75t_L g15506 ( 
.A(n_14099),
.B(n_13862),
.Y(n_15506)
);

AOI21xp33_ASAP7_75t_L g15507 ( 
.A1(n_14142),
.A2(n_13783),
.B(n_13781),
.Y(n_15507)
);

AND2x2_ASAP7_75t_L g15508 ( 
.A(n_14437),
.B(n_14443),
.Y(n_15508)
);

AND2x2_ASAP7_75t_L g15509 ( 
.A(n_14463),
.B(n_10870),
.Y(n_15509)
);

AND2x4_ASAP7_75t_SL g15510 ( 
.A(n_14433),
.B(n_10135),
.Y(n_15510)
);

INVx1_ASAP7_75t_L g15511 ( 
.A(n_14633),
.Y(n_15511)
);

AND2x2_ASAP7_75t_L g15512 ( 
.A(n_14468),
.B(n_10870),
.Y(n_15512)
);

NAND2xp5_ASAP7_75t_L g15513 ( 
.A(n_14771),
.B(n_13605),
.Y(n_15513)
);

INVx2_ASAP7_75t_L g15514 ( 
.A(n_14649),
.Y(n_15514)
);

AND2x2_ASAP7_75t_L g15515 ( 
.A(n_14469),
.B(n_10870),
.Y(n_15515)
);

AND2x4_ASAP7_75t_L g15516 ( 
.A(n_14161),
.B(n_11357),
.Y(n_15516)
);

AND2x2_ASAP7_75t_L g15517 ( 
.A(n_14563),
.B(n_11009),
.Y(n_15517)
);

BUFx2_ASAP7_75t_L g15518 ( 
.A(n_14298),
.Y(n_15518)
);

INVx2_ASAP7_75t_L g15519 ( 
.A(n_14650),
.Y(n_15519)
);

INVx1_ASAP7_75t_L g15520 ( 
.A(n_14779),
.Y(n_15520)
);

BUFx3_ASAP7_75t_L g15521 ( 
.A(n_14994),
.Y(n_15521)
);

OR2x2_ASAP7_75t_L g15522 ( 
.A(n_14813),
.B(n_13920),
.Y(n_15522)
);

OR2x2_ASAP7_75t_L g15523 ( 
.A(n_14833),
.B(n_13936),
.Y(n_15523)
);

AND2x2_ASAP7_75t_L g15524 ( 
.A(n_14951),
.B(n_11009),
.Y(n_15524)
);

AND2x2_ASAP7_75t_L g15525 ( 
.A(n_14388),
.B(n_11009),
.Y(n_15525)
);

AND2x2_ASAP7_75t_L g15526 ( 
.A(n_14180),
.B(n_11009),
.Y(n_15526)
);

AND2x2_ASAP7_75t_L g15527 ( 
.A(n_14182),
.B(n_11009),
.Y(n_15527)
);

OR2x2_ASAP7_75t_L g15528 ( 
.A(n_14839),
.B(n_13606),
.Y(n_15528)
);

AO21x2_ASAP7_75t_L g15529 ( 
.A1(n_14168),
.A2(n_14272),
.B(n_14034),
.Y(n_15529)
);

NAND2xp5_ASAP7_75t_L g15530 ( 
.A(n_14842),
.B(n_13610),
.Y(n_15530)
);

BUFx2_ASAP7_75t_L g15531 ( 
.A(n_14016),
.Y(n_15531)
);

INVxp67_ASAP7_75t_SL g15532 ( 
.A(n_14333),
.Y(n_15532)
);

AND2x4_ASAP7_75t_SL g15533 ( 
.A(n_14533),
.B(n_10135),
.Y(n_15533)
);

AOI222xp33_ASAP7_75t_L g15534 ( 
.A1(n_14021),
.A2(n_9911),
.B1(n_9872),
.B2(n_9941),
.C1(n_9892),
.C2(n_9838),
.Y(n_15534)
);

INVxp67_ASAP7_75t_SL g15535 ( 
.A(n_14381),
.Y(n_15535)
);

INVx2_ASAP7_75t_L g15536 ( 
.A(n_14663),
.Y(n_15536)
);

BUFx3_ASAP7_75t_L g15537 ( 
.A(n_14573),
.Y(n_15537)
);

INVx1_ASAP7_75t_L g15538 ( 
.A(n_14867),
.Y(n_15538)
);

INVx1_ASAP7_75t_L g15539 ( 
.A(n_14867),
.Y(n_15539)
);

INVx2_ASAP7_75t_L g15540 ( 
.A(n_14671),
.Y(n_15540)
);

AOI221xp5_ASAP7_75t_L g15541 ( 
.A1(n_14170),
.A2(n_11627),
.B1(n_11603),
.B2(n_10879),
.C(n_9892),
.Y(n_15541)
);

AOI22xp33_ASAP7_75t_L g15542 ( 
.A1(n_14167),
.A2(n_9283),
.B1(n_10124),
.B2(n_9590),
.Y(n_15542)
);

INVxp67_ASAP7_75t_L g15543 ( 
.A(n_14148),
.Y(n_15543)
);

OR2x2_ASAP7_75t_L g15544 ( 
.A(n_14501),
.B(n_13612),
.Y(n_15544)
);

INVx2_ASAP7_75t_L g15545 ( 
.A(n_14783),
.Y(n_15545)
);

INVx8_ASAP7_75t_L g15546 ( 
.A(n_14642),
.Y(n_15546)
);

INVx2_ASAP7_75t_L g15547 ( 
.A(n_14788),
.Y(n_15547)
);

INVx1_ASAP7_75t_L g15548 ( 
.A(n_14877),
.Y(n_15548)
);

INVx1_ASAP7_75t_L g15549 ( 
.A(n_14877),
.Y(n_15549)
);

INVx1_ASAP7_75t_L g15550 ( 
.A(n_14944),
.Y(n_15550)
);

AND2x2_ASAP7_75t_L g15551 ( 
.A(n_14818),
.B(n_10244),
.Y(n_15551)
);

INVx3_ASAP7_75t_L g15552 ( 
.A(n_14459),
.Y(n_15552)
);

NAND2xp5_ASAP7_75t_L g15553 ( 
.A(n_14868),
.B(n_13613),
.Y(n_15553)
);

OR2x2_ASAP7_75t_L g15554 ( 
.A(n_14531),
.B(n_13615),
.Y(n_15554)
);

INVx2_ASAP7_75t_L g15555 ( 
.A(n_14789),
.Y(n_15555)
);

INVx3_ASAP7_75t_L g15556 ( 
.A(n_14511),
.Y(n_15556)
);

BUFx6f_ASAP7_75t_L g15557 ( 
.A(n_14931),
.Y(n_15557)
);

INVx1_ASAP7_75t_L g15558 ( 
.A(n_14937),
.Y(n_15558)
);

INVx1_ASAP7_75t_L g15559 ( 
.A(n_14971),
.Y(n_15559)
);

INVxp67_ASAP7_75t_L g15560 ( 
.A(n_14370),
.Y(n_15560)
);

INVx2_ASAP7_75t_L g15561 ( 
.A(n_14795),
.Y(n_15561)
);

OA21x2_ASAP7_75t_L g15562 ( 
.A1(n_14883),
.A2(n_13436),
.B(n_13414),
.Y(n_15562)
);

AND2x2_ASAP7_75t_L g15563 ( 
.A(n_14624),
.B(n_10244),
.Y(n_15563)
);

INVx1_ASAP7_75t_L g15564 ( 
.A(n_14835),
.Y(n_15564)
);

INVxp67_ASAP7_75t_SL g15565 ( 
.A(n_14080),
.Y(n_15565)
);

AND2x4_ASAP7_75t_L g15566 ( 
.A(n_14313),
.B(n_11359),
.Y(n_15566)
);

CKINVDCx8_ASAP7_75t_R g15567 ( 
.A(n_14496),
.Y(n_15567)
);

AND2x2_ASAP7_75t_L g15568 ( 
.A(n_14770),
.B(n_10244),
.Y(n_15568)
);

INVx1_ASAP7_75t_L g15569 ( 
.A(n_14215),
.Y(n_15569)
);

INVx3_ASAP7_75t_L g15570 ( 
.A(n_14516),
.Y(n_15570)
);

INVx1_ASAP7_75t_L g15571 ( 
.A(n_14215),
.Y(n_15571)
);

BUFx2_ASAP7_75t_L g15572 ( 
.A(n_14016),
.Y(n_15572)
);

NAND2xp5_ASAP7_75t_L g15573 ( 
.A(n_14907),
.B(n_13786),
.Y(n_15573)
);

INVx1_ASAP7_75t_L g15574 ( 
.A(n_14287),
.Y(n_15574)
);

INVx2_ASAP7_75t_L g15575 ( 
.A(n_14797),
.Y(n_15575)
);

INVx2_ASAP7_75t_L g15576 ( 
.A(n_14798),
.Y(n_15576)
);

INVx2_ASAP7_75t_L g15577 ( 
.A(n_14803),
.Y(n_15577)
);

AND2x2_ASAP7_75t_L g15578 ( 
.A(n_14398),
.B(n_10408),
.Y(n_15578)
);

BUFx6f_ASAP7_75t_L g15579 ( 
.A(n_14931),
.Y(n_15579)
);

INVx1_ASAP7_75t_L g15580 ( 
.A(n_14287),
.Y(n_15580)
);

AND2x2_ASAP7_75t_L g15581 ( 
.A(n_14410),
.B(n_10408),
.Y(n_15581)
);

INVx2_ASAP7_75t_L g15582 ( 
.A(n_14814),
.Y(n_15582)
);

INVx2_ASAP7_75t_L g15583 ( 
.A(n_14418),
.Y(n_15583)
);

INVx2_ASAP7_75t_L g15584 ( 
.A(n_14832),
.Y(n_15584)
);

AND2x2_ASAP7_75t_L g15585 ( 
.A(n_14414),
.B(n_10408),
.Y(n_15585)
);

INVx1_ASAP7_75t_L g15586 ( 
.A(n_14307),
.Y(n_15586)
);

OR2x2_ASAP7_75t_L g15587 ( 
.A(n_14574),
.B(n_13787),
.Y(n_15587)
);

NAND2xp5_ASAP7_75t_SL g15588 ( 
.A(n_14276),
.B(n_11144),
.Y(n_15588)
);

OR2x2_ASAP7_75t_L g15589 ( 
.A(n_14585),
.B(n_13788),
.Y(n_15589)
);

AND2x2_ASAP7_75t_L g15590 ( 
.A(n_14430),
.B(n_10427),
.Y(n_15590)
);

AND2x2_ASAP7_75t_L g15591 ( 
.A(n_14432),
.B(n_10427),
.Y(n_15591)
);

BUFx2_ASAP7_75t_L g15592 ( 
.A(n_14273),
.Y(n_15592)
);

AND2x2_ASAP7_75t_L g15593 ( 
.A(n_14553),
.B(n_10427),
.Y(n_15593)
);

AOI21xp5_ASAP7_75t_L g15594 ( 
.A1(n_14065),
.A2(n_13370),
.B(n_13190),
.Y(n_15594)
);

BUFx2_ASAP7_75t_L g15595 ( 
.A(n_14054),
.Y(n_15595)
);

AO21x2_ASAP7_75t_L g15596 ( 
.A1(n_14055),
.A2(n_14124),
.B(n_14334),
.Y(n_15596)
);

INVx1_ASAP7_75t_L g15597 ( 
.A(n_14307),
.Y(n_15597)
);

INVx1_ASAP7_75t_L g15598 ( 
.A(n_14856),
.Y(n_15598)
);

AND2x2_ASAP7_75t_L g15599 ( 
.A(n_14558),
.B(n_10437),
.Y(n_15599)
);

NAND2xp5_ASAP7_75t_L g15600 ( 
.A(n_14429),
.B(n_13790),
.Y(n_15600)
);

OR2x2_ASAP7_75t_L g15601 ( 
.A(n_14602),
.B(n_13792),
.Y(n_15601)
);

AOI21xp33_ASAP7_75t_SL g15602 ( 
.A1(n_14056),
.A2(n_13336),
.B(n_10846),
.Y(n_15602)
);

INVx1_ASAP7_75t_L g15603 ( 
.A(n_14275),
.Y(n_15603)
);

INVx1_ASAP7_75t_L g15604 ( 
.A(n_14359),
.Y(n_15604)
);

INVx2_ASAP7_75t_L g15605 ( 
.A(n_14346),
.Y(n_15605)
);

OAI21xp5_ASAP7_75t_L g15606 ( 
.A1(n_14060),
.A2(n_13190),
.B(n_13121),
.Y(n_15606)
);

BUFx3_ASAP7_75t_L g15607 ( 
.A(n_14640),
.Y(n_15607)
);

AND2x2_ASAP7_75t_L g15608 ( 
.A(n_14560),
.B(n_10437),
.Y(n_15608)
);

INVx2_ASAP7_75t_SL g15609 ( 
.A(n_14916),
.Y(n_15609)
);

AND2x2_ASAP7_75t_L g15610 ( 
.A(n_14561),
.B(n_10437),
.Y(n_15610)
);

BUFx12f_ASAP7_75t_L g15611 ( 
.A(n_14848),
.Y(n_15611)
);

INVx3_ASAP7_75t_L g15612 ( 
.A(n_14791),
.Y(n_15612)
);

INVx2_ASAP7_75t_L g15613 ( 
.A(n_14349),
.Y(n_15613)
);

INVx1_ASAP7_75t_L g15614 ( 
.A(n_14359),
.Y(n_15614)
);

BUFx3_ASAP7_75t_L g15615 ( 
.A(n_14647),
.Y(n_15615)
);

INVx1_ASAP7_75t_L g15616 ( 
.A(n_14368),
.Y(n_15616)
);

AOI31xp33_ASAP7_75t_SL g15617 ( 
.A1(n_14274),
.A2(n_11303),
.A3(n_11261),
.B(n_11340),
.Y(n_15617)
);

INVx1_ASAP7_75t_L g15618 ( 
.A(n_14368),
.Y(n_15618)
);

AO21x2_ASAP7_75t_L g15619 ( 
.A1(n_14191),
.A2(n_13236),
.B(n_13796),
.Y(n_15619)
);

INVx2_ASAP7_75t_L g15620 ( 
.A(n_14353),
.Y(n_15620)
);

NAND2xp5_ASAP7_75t_L g15621 ( 
.A(n_14851),
.B(n_13815),
.Y(n_15621)
);

INVx2_ASAP7_75t_SL g15622 ( 
.A(n_14916),
.Y(n_15622)
);

AND2x4_ASAP7_75t_L g15623 ( 
.A(n_14318),
.B(n_11359),
.Y(n_15623)
);

NAND2xp5_ASAP7_75t_L g15624 ( 
.A(n_14258),
.B(n_13816),
.Y(n_15624)
);

INVx2_ASAP7_75t_L g15625 ( 
.A(n_14793),
.Y(n_15625)
);

INVx1_ASAP7_75t_L g15626 ( 
.A(n_14390),
.Y(n_15626)
);

INVx1_ASAP7_75t_L g15627 ( 
.A(n_14390),
.Y(n_15627)
);

AND2x2_ASAP7_75t_L g15628 ( 
.A(n_14491),
.B(n_10492),
.Y(n_15628)
);

INVxp67_ASAP7_75t_SL g15629 ( 
.A(n_14404),
.Y(n_15629)
);

INVx1_ASAP7_75t_L g15630 ( 
.A(n_14396),
.Y(n_15630)
);

AND2x2_ASAP7_75t_L g15631 ( 
.A(n_14498),
.B(n_10492),
.Y(n_15631)
);

INVx2_ASAP7_75t_L g15632 ( 
.A(n_14806),
.Y(n_15632)
);

CKINVDCx20_ASAP7_75t_R g15633 ( 
.A(n_14662),
.Y(n_15633)
);

INVx1_ASAP7_75t_SL g15634 ( 
.A(n_14216),
.Y(n_15634)
);

INVx1_ASAP7_75t_L g15635 ( 
.A(n_14396),
.Y(n_15635)
);

AND2x2_ASAP7_75t_L g15636 ( 
.A(n_14512),
.B(n_10492),
.Y(n_15636)
);

INVx1_ASAP7_75t_L g15637 ( 
.A(n_14972),
.Y(n_15637)
);

INVx2_ASAP7_75t_L g15638 ( 
.A(n_14195),
.Y(n_15638)
);

INVx2_ASAP7_75t_L g15639 ( 
.A(n_14674),
.Y(n_15639)
);

AOI33xp33_ASAP7_75t_L g15640 ( 
.A1(n_14393),
.A2(n_13827),
.A3(n_13825),
.B1(n_13829),
.B2(n_13826),
.B3(n_13821),
.Y(n_15640)
);

INVx2_ASAP7_75t_L g15641 ( 
.A(n_14676),
.Y(n_15641)
);

NAND2x1_ASAP7_75t_L g15642 ( 
.A(n_14338),
.B(n_13445),
.Y(n_15642)
);

AND2x2_ASAP7_75t_L g15643 ( 
.A(n_14518),
.B(n_10553),
.Y(n_15643)
);

AOI22xp33_ASAP7_75t_L g15644 ( 
.A1(n_14051),
.A2(n_10124),
.B1(n_9590),
.B2(n_9965),
.Y(n_15644)
);

INVx3_ASAP7_75t_SL g15645 ( 
.A(n_14848),
.Y(n_15645)
);

AOI33xp33_ASAP7_75t_L g15646 ( 
.A1(n_14257),
.A2(n_14019),
.A3(n_14190),
.B1(n_14762),
.B2(n_14292),
.B3(n_14325),
.Y(n_15646)
);

AND2x4_ASAP7_75t_L g15647 ( 
.A(n_14073),
.B(n_11359),
.Y(n_15647)
);

INVx1_ASAP7_75t_L g15648 ( 
.A(n_14435),
.Y(n_15648)
);

NAND2xp5_ASAP7_75t_L g15649 ( 
.A(n_14277),
.B(n_13831),
.Y(n_15649)
);

INVx1_ASAP7_75t_L g15650 ( 
.A(n_14442),
.Y(n_15650)
);

INVx1_ASAP7_75t_L g15651 ( 
.A(n_14444),
.Y(n_15651)
);

OR2x2_ASAP7_75t_L g15652 ( 
.A(n_14616),
.B(n_13833),
.Y(n_15652)
);

HB1xp67_ASAP7_75t_L g15653 ( 
.A(n_14505),
.Y(n_15653)
);

NOR2xp33_ASAP7_75t_SL g15654 ( 
.A(n_14268),
.B(n_14199),
.Y(n_15654)
);

AOI22xp33_ASAP7_75t_SL g15655 ( 
.A1(n_14115),
.A2(n_9872),
.B1(n_9892),
.B2(n_9838),
.Y(n_15655)
);

AND2x2_ASAP7_75t_L g15656 ( 
.A(n_14523),
.B(n_10553),
.Y(n_15656)
);

NOR2x1_ASAP7_75t_L g15657 ( 
.A(n_14288),
.B(n_13837),
.Y(n_15657)
);

AND2x4_ASAP7_75t_L g15658 ( 
.A(n_14466),
.B(n_11359),
.Y(n_15658)
);

INVx1_ASAP7_75t_L g15659 ( 
.A(n_14450),
.Y(n_15659)
);

AND2x2_ASAP7_75t_L g15660 ( 
.A(n_14534),
.B(n_10553),
.Y(n_15660)
);

BUFx3_ASAP7_75t_L g15661 ( 
.A(n_14731),
.Y(n_15661)
);

AOI21x1_ASAP7_75t_L g15662 ( 
.A1(n_14505),
.A2(n_13452),
.B(n_13436),
.Y(n_15662)
);

INVx2_ASAP7_75t_L g15663 ( 
.A(n_14677),
.Y(n_15663)
);

BUFx6f_ASAP7_75t_L g15664 ( 
.A(n_14582),
.Y(n_15664)
);

INVx1_ASAP7_75t_L g15665 ( 
.A(n_14497),
.Y(n_15665)
);

NAND2xp5_ASAP7_75t_L g15666 ( 
.A(n_14508),
.B(n_13839),
.Y(n_15666)
);

AND2x2_ASAP7_75t_L g15667 ( 
.A(n_14536),
.B(n_10555),
.Y(n_15667)
);

INVx2_ASAP7_75t_L g15668 ( 
.A(n_14678),
.Y(n_15668)
);

INVx1_ASAP7_75t_L g15669 ( 
.A(n_14567),
.Y(n_15669)
);

INVx2_ASAP7_75t_L g15670 ( 
.A(n_14543),
.Y(n_15670)
);

NAND2xp5_ASAP7_75t_L g15671 ( 
.A(n_14707),
.B(n_13844),
.Y(n_15671)
);

INVx2_ASAP7_75t_SL g15672 ( 
.A(n_14959),
.Y(n_15672)
);

INVx1_ASAP7_75t_L g15673 ( 
.A(n_14487),
.Y(n_15673)
);

INVx1_ASAP7_75t_L g15674 ( 
.A(n_14365),
.Y(n_15674)
);

INVx1_ASAP7_75t_L g15675 ( 
.A(n_14372),
.Y(n_15675)
);

INVx2_ASAP7_75t_L g15676 ( 
.A(n_14550),
.Y(n_15676)
);

BUFx3_ASAP7_75t_L g15677 ( 
.A(n_14927),
.Y(n_15677)
);

INVx2_ASAP7_75t_L g15678 ( 
.A(n_14552),
.Y(n_15678)
);

AND2x2_ASAP7_75t_L g15679 ( 
.A(n_14242),
.B(n_10555),
.Y(n_15679)
);

OR2x2_ASAP7_75t_L g15680 ( 
.A(n_14237),
.B(n_13847),
.Y(n_15680)
);

AND2x4_ASAP7_75t_L g15681 ( 
.A(n_14479),
.B(n_11359),
.Y(n_15681)
);

INVxp67_ASAP7_75t_L g15682 ( 
.A(n_14940),
.Y(n_15682)
);

INVx1_ASAP7_75t_L g15683 ( 
.A(n_14569),
.Y(n_15683)
);

INVx1_ASAP7_75t_L g15684 ( 
.A(n_14569),
.Y(n_15684)
);

INVx2_ASAP7_75t_L g15685 ( 
.A(n_14290),
.Y(n_15685)
);

INVxp67_ASAP7_75t_L g15686 ( 
.A(n_14568),
.Y(n_15686)
);

AND2x2_ASAP7_75t_L g15687 ( 
.A(n_14471),
.B(n_14670),
.Y(n_15687)
);

INVx1_ASAP7_75t_L g15688 ( 
.A(n_14597),
.Y(n_15688)
);

OR2x2_ASAP7_75t_L g15689 ( 
.A(n_14244),
.B(n_10217),
.Y(n_15689)
);

AND2x2_ASAP7_75t_L g15690 ( 
.A(n_14694),
.B(n_10555),
.Y(n_15690)
);

INVx3_ASAP7_75t_L g15691 ( 
.A(n_14626),
.Y(n_15691)
);

OR2x2_ASAP7_75t_L g15692 ( 
.A(n_14169),
.B(n_14302),
.Y(n_15692)
);

NAND2xp5_ASAP7_75t_L g15693 ( 
.A(n_14489),
.B(n_13902),
.Y(n_15693)
);

AND2x4_ASAP7_75t_L g15694 ( 
.A(n_14495),
.B(n_11455),
.Y(n_15694)
);

AND2x2_ASAP7_75t_L g15695 ( 
.A(n_14358),
.B(n_10592),
.Y(n_15695)
);

AO31x2_ASAP7_75t_L g15696 ( 
.A1(n_14754),
.A2(n_13908),
.A3(n_13909),
.B(n_13905),
.Y(n_15696)
);

NOR2x1p5_ASAP7_75t_L g15697 ( 
.A(n_14105),
.B(n_10135),
.Y(n_15697)
);

AND2x2_ASAP7_75t_L g15698 ( 
.A(n_14360),
.B(n_10592),
.Y(n_15698)
);

AOI22xp33_ASAP7_75t_L g15699 ( 
.A1(n_14217),
.A2(n_9590),
.B1(n_9965),
.B2(n_11603),
.Y(n_15699)
);

INVx2_ASAP7_75t_L g15700 ( 
.A(n_14293),
.Y(n_15700)
);

AND2x4_ASAP7_75t_L g15701 ( 
.A(n_14658),
.B(n_11455),
.Y(n_15701)
);

AND2x4_ASAP7_75t_L g15702 ( 
.A(n_14590),
.B(n_11455),
.Y(n_15702)
);

INVx1_ASAP7_75t_L g15703 ( 
.A(n_14597),
.Y(n_15703)
);

OR2x2_ASAP7_75t_L g15704 ( 
.A(n_14312),
.B(n_10965),
.Y(n_15704)
);

AND2x2_ASAP7_75t_L g15705 ( 
.A(n_14367),
.B(n_10592),
.Y(n_15705)
);

INVx1_ASAP7_75t_L g15706 ( 
.A(n_14452),
.Y(n_15706)
);

INVx2_ASAP7_75t_L g15707 ( 
.A(n_14301),
.Y(n_15707)
);

INVx2_ASAP7_75t_L g15708 ( 
.A(n_14315),
.Y(n_15708)
);

HB1xp67_ASAP7_75t_L g15709 ( 
.A(n_14825),
.Y(n_15709)
);

INVxp67_ASAP7_75t_SL g15710 ( 
.A(n_14053),
.Y(n_15710)
);

INVx2_ASAP7_75t_L g15711 ( 
.A(n_14323),
.Y(n_15711)
);

INVx1_ASAP7_75t_L g15712 ( 
.A(n_14513),
.Y(n_15712)
);

INVx1_ASAP7_75t_L g15713 ( 
.A(n_14236),
.Y(n_15713)
);

INVx1_ASAP7_75t_L g15714 ( 
.A(n_14240),
.Y(n_15714)
);

INVx2_ASAP7_75t_L g15715 ( 
.A(n_14339),
.Y(n_15715)
);

INVxp67_ASAP7_75t_SL g15716 ( 
.A(n_14043),
.Y(n_15716)
);

INVx1_ASAP7_75t_L g15717 ( 
.A(n_14733),
.Y(n_15717)
);

INVx1_ASAP7_75t_L g15718 ( 
.A(n_14745),
.Y(n_15718)
);

INVx2_ASAP7_75t_L g15719 ( 
.A(n_14840),
.Y(n_15719)
);

AND2x2_ASAP7_75t_L g15720 ( 
.A(n_14959),
.B(n_14978),
.Y(n_15720)
);

INVx2_ASAP7_75t_L g15721 ( 
.A(n_14475),
.Y(n_15721)
);

BUFx3_ASAP7_75t_L g15722 ( 
.A(n_14800),
.Y(n_15722)
);

INVx1_ASAP7_75t_L g15723 ( 
.A(n_14223),
.Y(n_15723)
);

INVx2_ASAP7_75t_L g15724 ( 
.A(n_14920),
.Y(n_15724)
);

INVx1_ASAP7_75t_L g15725 ( 
.A(n_14464),
.Y(n_15725)
);

HB1xp67_ASAP7_75t_L g15726 ( 
.A(n_14329),
.Y(n_15726)
);

INVx2_ASAP7_75t_L g15727 ( 
.A(n_14928),
.Y(n_15727)
);

BUFx2_ASAP7_75t_L g15728 ( 
.A(n_14054),
.Y(n_15728)
);

AND2x4_ASAP7_75t_L g15729 ( 
.A(n_14978),
.B(n_11455),
.Y(n_15729)
);

BUFx2_ASAP7_75t_L g15730 ( 
.A(n_14352),
.Y(n_15730)
);

INVx1_ASAP7_75t_L g15731 ( 
.A(n_14464),
.Y(n_15731)
);

AND2x2_ASAP7_75t_L g15732 ( 
.A(n_14984),
.B(n_10623),
.Y(n_15732)
);

OR2x2_ASAP7_75t_L g15733 ( 
.A(n_14163),
.B(n_10974),
.Y(n_15733)
);

INVx3_ASAP7_75t_L g15734 ( 
.A(n_14919),
.Y(n_15734)
);

INVx2_ASAP7_75t_L g15735 ( 
.A(n_14816),
.Y(n_15735)
);

INVx2_ASAP7_75t_SL g15736 ( 
.A(n_14984),
.Y(n_15736)
);

INVx1_ASAP7_75t_L g15737 ( 
.A(n_14305),
.Y(n_15737)
);

BUFx2_ASAP7_75t_L g15738 ( 
.A(n_14352),
.Y(n_15738)
);

NAND2xp5_ASAP7_75t_L g15739 ( 
.A(n_14724),
.B(n_13912),
.Y(n_15739)
);

AND2x2_ASAP7_75t_L g15740 ( 
.A(n_14988),
.B(n_10623),
.Y(n_15740)
);

NOR2xp33_ASAP7_75t_L g15741 ( 
.A(n_14809),
.B(n_11463),
.Y(n_15741)
);

BUFx2_ASAP7_75t_L g15742 ( 
.A(n_14086),
.Y(n_15742)
);

AND2x2_ASAP7_75t_L g15743 ( 
.A(n_14988),
.B(n_10623),
.Y(n_15743)
);

INVx5_ASAP7_75t_SL g15744 ( 
.A(n_14587),
.Y(n_15744)
);

BUFx3_ASAP7_75t_L g15745 ( 
.A(n_14831),
.Y(n_15745)
);

INVxp67_ASAP7_75t_L g15746 ( 
.A(n_14942),
.Y(n_15746)
);

BUFx6f_ASAP7_75t_L g15747 ( 
.A(n_14592),
.Y(n_15747)
);

AND2x2_ASAP7_75t_L g15748 ( 
.A(n_14947),
.B(n_11455),
.Y(n_15748)
);

INVx2_ASAP7_75t_L g15749 ( 
.A(n_14976),
.Y(n_15749)
);

INVx2_ASAP7_75t_L g15750 ( 
.A(n_14977),
.Y(n_15750)
);

OAI222xp33_ASAP7_75t_L g15751 ( 
.A1(n_14300),
.A2(n_10461),
.B1(n_10846),
.B2(n_10893),
.C1(n_10892),
.C2(n_10831),
.Y(n_15751)
);

AOI22xp33_ASAP7_75t_SL g15752 ( 
.A1(n_14005),
.A2(n_9872),
.B1(n_9892),
.B2(n_9838),
.Y(n_15752)
);

INVxp67_ASAP7_75t_SL g15753 ( 
.A(n_14137),
.Y(n_15753)
);

INVx2_ASAP7_75t_L g15754 ( 
.A(n_14980),
.Y(n_15754)
);

AND2x4_ASAP7_75t_L g15755 ( 
.A(n_14925),
.B(n_11509),
.Y(n_15755)
);

AND2x2_ASAP7_75t_L g15756 ( 
.A(n_14587),
.B(n_11509),
.Y(n_15756)
);

INVx1_ASAP7_75t_L g15757 ( 
.A(n_14330),
.Y(n_15757)
);

AND2x2_ASAP7_75t_L g15758 ( 
.A(n_14591),
.B(n_11509),
.Y(n_15758)
);

INVx1_ASAP7_75t_L g15759 ( 
.A(n_14347),
.Y(n_15759)
);

NAND2xp5_ASAP7_75t_L g15760 ( 
.A(n_14705),
.B(n_13915),
.Y(n_15760)
);

INVx1_ASAP7_75t_L g15761 ( 
.A(n_14767),
.Y(n_15761)
);

AND2x4_ASAP7_75t_L g15762 ( 
.A(n_14936),
.B(n_11509),
.Y(n_15762)
);

INVx4_ASAP7_75t_L g15763 ( 
.A(n_14591),
.Y(n_15763)
);

AND2x4_ASAP7_75t_L g15764 ( 
.A(n_14641),
.B(n_11509),
.Y(n_15764)
);

INVx2_ASAP7_75t_L g15765 ( 
.A(n_14987),
.Y(n_15765)
);

AND2x2_ASAP7_75t_L g15766 ( 
.A(n_14641),
.B(n_11113),
.Y(n_15766)
);

AND2x2_ASAP7_75t_L g15767 ( 
.A(n_14992),
.B(n_11113),
.Y(n_15767)
);

INVx2_ASAP7_75t_L g15768 ( 
.A(n_14820),
.Y(n_15768)
);

INVx1_ASAP7_75t_L g15769 ( 
.A(n_14361),
.Y(n_15769)
);

INVx2_ASAP7_75t_SL g15770 ( 
.A(n_14785),
.Y(n_15770)
);

AND2x2_ASAP7_75t_L g15771 ( 
.A(n_14934),
.B(n_11113),
.Y(n_15771)
);

INVx2_ASAP7_75t_L g15772 ( 
.A(n_14841),
.Y(n_15772)
);

AND2x4_ASAP7_75t_L g15773 ( 
.A(n_14855),
.B(n_11624),
.Y(n_15773)
);

INVx1_ASAP7_75t_L g15774 ( 
.A(n_14826),
.Y(n_15774)
);

OR2x2_ASAP7_75t_L g15775 ( 
.A(n_14165),
.B(n_10974),
.Y(n_15775)
);

INVx1_ASAP7_75t_L g15776 ( 
.A(n_14858),
.Y(n_15776)
);

AND2x4_ASAP7_75t_L g15777 ( 
.A(n_14943),
.B(n_11624),
.Y(n_15777)
);

OR2x2_ASAP7_75t_L g15778 ( 
.A(n_14426),
.B(n_10975),
.Y(n_15778)
);

AND2x2_ASAP7_75t_L g15779 ( 
.A(n_14949),
.B(n_11116),
.Y(n_15779)
);

OR2x2_ASAP7_75t_L g15780 ( 
.A(n_14261),
.B(n_10975),
.Y(n_15780)
);

INVx1_ASAP7_75t_L g15781 ( 
.A(n_14875),
.Y(n_15781)
);

AND2x2_ASAP7_75t_L g15782 ( 
.A(n_14952),
.B(n_11116),
.Y(n_15782)
);

AND2x2_ASAP7_75t_L g15783 ( 
.A(n_14957),
.B(n_11116),
.Y(n_15783)
);

INVx1_ASAP7_75t_L g15784 ( 
.A(n_14878),
.Y(n_15784)
);

AND2x2_ASAP7_75t_L g15785 ( 
.A(n_14962),
.B(n_11151),
.Y(n_15785)
);

AOI22xp33_ASAP7_75t_L g15786 ( 
.A1(n_14269),
.A2(n_9590),
.B1(n_9965),
.B2(n_11603),
.Y(n_15786)
);

NAND2xp5_ASAP7_75t_L g15787 ( 
.A(n_14537),
.B(n_13916),
.Y(n_15787)
);

INVx2_ASAP7_75t_L g15788 ( 
.A(n_14857),
.Y(n_15788)
);

INVx3_ASAP7_75t_L g15789 ( 
.A(n_14785),
.Y(n_15789)
);

AO21x2_ASAP7_75t_L g15790 ( 
.A1(n_14133),
.A2(n_13798),
.B(n_13796),
.Y(n_15790)
);

BUFx2_ASAP7_75t_L g15791 ( 
.A(n_14086),
.Y(n_15791)
);

AND2x4_ASAP7_75t_L g15792 ( 
.A(n_14860),
.B(n_11624),
.Y(n_15792)
);

OR2x2_ASAP7_75t_L g15793 ( 
.A(n_14672),
.B(n_10987),
.Y(n_15793)
);

NAND2xp5_ASAP7_75t_L g15794 ( 
.A(n_14344),
.B(n_13917),
.Y(n_15794)
);

OAI22xp5_ASAP7_75t_L g15795 ( 
.A1(n_14205),
.A2(n_9872),
.B1(n_9892),
.B2(n_9838),
.Y(n_15795)
);

AND2x2_ASAP7_75t_L g15796 ( 
.A(n_14964),
.B(n_11151),
.Y(n_15796)
);

INVx4_ASAP7_75t_L g15797 ( 
.A(n_14862),
.Y(n_15797)
);

INVx1_ASAP7_75t_L g15798 ( 
.A(n_14945),
.Y(n_15798)
);

INVx3_ASAP7_75t_L g15799 ( 
.A(n_14874),
.Y(n_15799)
);

INVx1_ASAP7_75t_L g15800 ( 
.A(n_14993),
.Y(n_15800)
);

AND2x2_ASAP7_75t_L g15801 ( 
.A(n_14967),
.B(n_11151),
.Y(n_15801)
);

AND2x2_ASAP7_75t_L g15802 ( 
.A(n_14968),
.B(n_11153),
.Y(n_15802)
);

INVx2_ASAP7_75t_L g15803 ( 
.A(n_14880),
.Y(n_15803)
);

INVx1_ASAP7_75t_L g15804 ( 
.A(n_14703),
.Y(n_15804)
);

INVx1_ASAP7_75t_L g15805 ( 
.A(n_14712),
.Y(n_15805)
);

BUFx2_ASAP7_75t_L g15806 ( 
.A(n_13993),
.Y(n_15806)
);

INVx1_ASAP7_75t_L g15807 ( 
.A(n_14715),
.Y(n_15807)
);

INVxp67_ASAP7_75t_L g15808 ( 
.A(n_14718),
.Y(n_15808)
);

INVx2_ASAP7_75t_L g15809 ( 
.A(n_14882),
.Y(n_15809)
);

INVxp67_ASAP7_75t_SL g15810 ( 
.A(n_14355),
.Y(n_15810)
);

INVx1_ASAP7_75t_L g15811 ( 
.A(n_14719),
.Y(n_15811)
);

AND2x2_ASAP7_75t_L g15812 ( 
.A(n_14969),
.B(n_11153),
.Y(n_15812)
);

AND2x2_ASAP7_75t_L g15813 ( 
.A(n_14885),
.B(n_11153),
.Y(n_15813)
);

HB1xp67_ASAP7_75t_L g15814 ( 
.A(n_14380),
.Y(n_15814)
);

INVx2_ASAP7_75t_L g15815 ( 
.A(n_14895),
.Y(n_15815)
);

NAND3xp33_ASAP7_75t_L g15816 ( 
.A(n_14184),
.B(n_13472),
.C(n_13452),
.Y(n_15816)
);

INVx1_ASAP7_75t_L g15817 ( 
.A(n_14768),
.Y(n_15817)
);

NAND2x1p5_ASAP7_75t_L g15818 ( 
.A(n_14075),
.B(n_8151),
.Y(n_15818)
);

AOI22xp33_ASAP7_75t_L g15819 ( 
.A1(n_14061),
.A2(n_14316),
.B1(n_14208),
.B2(n_14102),
.Y(n_15819)
);

OR2x2_ASAP7_75t_L g15820 ( 
.A(n_14689),
.B(n_10987),
.Y(n_15820)
);

AND2x2_ASAP7_75t_L g15821 ( 
.A(n_14901),
.B(n_11182),
.Y(n_15821)
);

INVx2_ASAP7_75t_L g15822 ( 
.A(n_14912),
.Y(n_15822)
);

AND2x2_ASAP7_75t_L g15823 ( 
.A(n_15001),
.B(n_11182),
.Y(n_15823)
);

INVx2_ASAP7_75t_L g15824 ( 
.A(n_14434),
.Y(n_15824)
);

INVx1_ASAP7_75t_L g15825 ( 
.A(n_14324),
.Y(n_15825)
);

INVx3_ASAP7_75t_L g15826 ( 
.A(n_14286),
.Y(n_15826)
);

INVx1_ASAP7_75t_L g15827 ( 
.A(n_14324),
.Y(n_15827)
);

INVx1_ASAP7_75t_L g15828 ( 
.A(n_14834),
.Y(n_15828)
);

OR2x2_ASAP7_75t_L g15829 ( 
.A(n_14143),
.B(n_10988),
.Y(n_15829)
);

INVx2_ASAP7_75t_L g15830 ( 
.A(n_14434),
.Y(n_15830)
);

HB1xp67_ASAP7_75t_L g15831 ( 
.A(n_14743),
.Y(n_15831)
);

AND2x2_ASAP7_75t_L g15832 ( 
.A(n_14327),
.B(n_11182),
.Y(n_15832)
);

INVx2_ASAP7_75t_L g15833 ( 
.A(n_14465),
.Y(n_15833)
);

HB1xp67_ASAP7_75t_L g15834 ( 
.A(n_14743),
.Y(n_15834)
);

BUFx2_ASAP7_75t_L g15835 ( 
.A(n_13993),
.Y(n_15835)
);

BUFx2_ASAP7_75t_L g15836 ( 
.A(n_14037),
.Y(n_15836)
);

AOI22xp33_ASAP7_75t_L g15837 ( 
.A1(n_14037),
.A2(n_9965),
.B1(n_11627),
.B2(n_11603),
.Y(n_15837)
);

AND2x4_ASAP7_75t_L g15838 ( 
.A(n_14804),
.B(n_11624),
.Y(n_15838)
);

HB1xp67_ASAP7_75t_L g15839 ( 
.A(n_14787),
.Y(n_15839)
);

NAND2xp5_ASAP7_75t_L g15840 ( 
.A(n_14289),
.B(n_13923),
.Y(n_15840)
);

INVx1_ASAP7_75t_L g15841 ( 
.A(n_14834),
.Y(n_15841)
);

AND2x2_ASAP7_75t_L g15842 ( 
.A(n_14342),
.B(n_14350),
.Y(n_15842)
);

AND2x4_ASAP7_75t_L g15843 ( 
.A(n_14583),
.B(n_11624),
.Y(n_15843)
);

HB1xp67_ASAP7_75t_L g15844 ( 
.A(n_14974),
.Y(n_15844)
);

AO21x2_ASAP7_75t_L g15845 ( 
.A1(n_14451),
.A2(n_13798),
.B(n_13472),
.Y(n_15845)
);

HB1xp67_ASAP7_75t_L g15846 ( 
.A(n_14241),
.Y(n_15846)
);

AND2x2_ASAP7_75t_L g15847 ( 
.A(n_14340),
.B(n_11221),
.Y(n_15847)
);

BUFx2_ASAP7_75t_L g15848 ( 
.A(n_14224),
.Y(n_15848)
);

INVx1_ASAP7_75t_L g15849 ( 
.A(n_14584),
.Y(n_15849)
);

HB1xp67_ASAP7_75t_L g15850 ( 
.A(n_14322),
.Y(n_15850)
);

INVx2_ASAP7_75t_L g15851 ( 
.A(n_14465),
.Y(n_15851)
);

AND2x2_ASAP7_75t_L g15852 ( 
.A(n_14378),
.B(n_11221),
.Y(n_15852)
);

INVx1_ASAP7_75t_L g15853 ( 
.A(n_14586),
.Y(n_15853)
);

INVx1_ASAP7_75t_L g15854 ( 
.A(n_14683),
.Y(n_15854)
);

INVx1_ASAP7_75t_L g15855 ( 
.A(n_14686),
.Y(n_15855)
);

AND2x2_ASAP7_75t_L g15856 ( 
.A(n_14224),
.B(n_11221),
.Y(n_15856)
);

INVxp67_ASAP7_75t_L g15857 ( 
.A(n_14504),
.Y(n_15857)
);

INVx2_ASAP7_75t_L g15858 ( 
.A(n_14467),
.Y(n_15858)
);

AND2x2_ASAP7_75t_L g15859 ( 
.A(n_14285),
.B(n_9068),
.Y(n_15859)
);

OR2x2_ASAP7_75t_L g15860 ( 
.A(n_14802),
.B(n_10988),
.Y(n_15860)
);

INVx2_ASAP7_75t_L g15861 ( 
.A(n_14467),
.Y(n_15861)
);

AND2x2_ASAP7_75t_L g15862 ( 
.A(n_14096),
.B(n_9068),
.Y(n_15862)
);

NAND2xp5_ASAP7_75t_L g15863 ( 
.A(n_14351),
.B(n_13928),
.Y(n_15863)
);

INVx1_ASAP7_75t_L g15864 ( 
.A(n_14688),
.Y(n_15864)
);

NOR2x1_ASAP7_75t_L g15865 ( 
.A(n_14935),
.B(n_13121),
.Y(n_15865)
);

NAND2xp5_ASAP7_75t_L g15866 ( 
.A(n_14876),
.B(n_14884),
.Y(n_15866)
);

INVx1_ASAP7_75t_L g15867 ( 
.A(n_14699),
.Y(n_15867)
);

AND2x2_ASAP7_75t_L g15868 ( 
.A(n_14096),
.B(n_9068),
.Y(n_15868)
);

AND2x2_ASAP7_75t_L g15869 ( 
.A(n_15075),
.B(n_14341),
.Y(n_15869)
);

NAND4xp25_ASAP7_75t_L g15870 ( 
.A(n_15273),
.B(n_14262),
.C(n_14256),
.D(n_14219),
.Y(n_15870)
);

AOI221xp5_ASAP7_75t_L g15871 ( 
.A1(n_15848),
.A2(n_14387),
.B1(n_14320),
.B2(n_14319),
.C(n_14623),
.Y(n_15871)
);

NAND2xp5_ASAP7_75t_L g15872 ( 
.A(n_15437),
.B(n_14796),
.Y(n_15872)
);

AOI22xp33_ASAP7_75t_L g15873 ( 
.A1(n_15529),
.A2(n_14155),
.B1(n_14421),
.B2(n_14635),
.Y(n_15873)
);

NAND2xp5_ASAP7_75t_L g15874 ( 
.A(n_15437),
.B(n_14970),
.Y(n_15874)
);

NAND3xp33_ASAP7_75t_L g15875 ( 
.A(n_15484),
.B(n_14470),
.C(n_14515),
.Y(n_15875)
);

AOI221xp5_ASAP7_75t_L g15876 ( 
.A1(n_15848),
.A2(n_14652),
.B1(n_14861),
.B2(n_14270),
.C(n_14913),
.Y(n_15876)
);

NOR2xp33_ASAP7_75t_L g15877 ( 
.A(n_15013),
.B(n_14995),
.Y(n_15877)
);

NAND2xp5_ASAP7_75t_L g15878 ( 
.A(n_15463),
.B(n_14986),
.Y(n_15878)
);

NAND2xp5_ASAP7_75t_L g15879 ( 
.A(n_15463),
.B(n_14845),
.Y(n_15879)
);

AND2x2_ASAP7_75t_L g15880 ( 
.A(n_15023),
.B(n_14030),
.Y(n_15880)
);

AOI22xp33_ASAP7_75t_SL g15881 ( 
.A1(n_15531),
.A2(n_14065),
.B1(n_14030),
.B2(n_14259),
.Y(n_15881)
);

AND2x2_ASAP7_75t_L g15882 ( 
.A(n_15032),
.B(n_14655),
.Y(n_15882)
);

AOI22xp33_ASAP7_75t_L g15883 ( 
.A1(n_15531),
.A2(n_14546),
.B1(n_14356),
.B2(n_14716),
.Y(n_15883)
);

AND2x2_ASAP7_75t_L g15884 ( 
.A(n_15182),
.B(n_14610),
.Y(n_15884)
);

AND2x2_ASAP7_75t_L g15885 ( 
.A(n_15012),
.B(n_14601),
.Y(n_15885)
);

NAND4xp25_ASAP7_75t_L g15886 ( 
.A(n_15819),
.B(n_14419),
.C(n_14384),
.D(n_14493),
.Y(n_15886)
);

NOR2xp33_ASAP7_75t_SL g15887 ( 
.A(n_15306),
.B(n_11463),
.Y(n_15887)
);

AND2x2_ASAP7_75t_L g15888 ( 
.A(n_15003),
.B(n_14259),
.Y(n_15888)
);

NAND3xp33_ASAP7_75t_L g15889 ( 
.A(n_15473),
.B(n_14881),
.C(n_14520),
.Y(n_15889)
);

OAI22xp5_ASAP7_75t_L g15890 ( 
.A1(n_15572),
.A2(n_14684),
.B1(n_14460),
.B2(n_14556),
.Y(n_15890)
);

AND2x2_ASAP7_75t_SL g15891 ( 
.A(n_15572),
.B(n_14554),
.Y(n_15891)
);

AOI221xp5_ASAP7_75t_L g15892 ( 
.A1(n_15473),
.A2(n_14918),
.B1(n_15002),
.B2(n_14908),
.C(n_14811),
.Y(n_15892)
);

NAND3xp33_ASAP7_75t_L g15893 ( 
.A(n_15518),
.B(n_14562),
.C(n_14915),
.Y(n_15893)
);

AND2x2_ASAP7_75t_L g15894 ( 
.A(n_15123),
.B(n_14695),
.Y(n_15894)
);

AND2x2_ASAP7_75t_L g15895 ( 
.A(n_15067),
.B(n_14698),
.Y(n_15895)
);

NAND2xp5_ASAP7_75t_L g15896 ( 
.A(n_15518),
.B(n_15078),
.Y(n_15896)
);

AOI22xp33_ASAP7_75t_L g15897 ( 
.A1(n_15842),
.A2(n_14397),
.B1(n_14382),
.B2(n_14648),
.Y(n_15897)
);

AND2x2_ASAP7_75t_L g15898 ( 
.A(n_15067),
.B(n_14805),
.Y(n_15898)
);

NAND2xp5_ASAP7_75t_L g15899 ( 
.A(n_15078),
.B(n_14896),
.Y(n_15899)
);

AND2x2_ASAP7_75t_L g15900 ( 
.A(n_15443),
.B(n_14903),
.Y(n_15900)
);

NOR3xp33_ASAP7_75t_SL g15901 ( 
.A(n_15346),
.B(n_14458),
.C(n_14729),
.Y(n_15901)
);

NOR3xp33_ASAP7_75t_L g15902 ( 
.A(n_15352),
.B(n_14596),
.C(n_14415),
.Y(n_15902)
);

NAND2xp5_ASAP7_75t_L g15903 ( 
.A(n_15213),
.B(n_14823),
.Y(n_15903)
);

OAI221xp5_ASAP7_75t_L g15904 ( 
.A1(n_15810),
.A2(n_14524),
.B1(n_14577),
.B2(n_14985),
.C(n_14924),
.Y(n_15904)
);

NAND3xp33_ASAP7_75t_L g15905 ( 
.A(n_15709),
.B(n_14887),
.C(n_14844),
.Y(n_15905)
);

AND2x2_ASAP7_75t_L g15906 ( 
.A(n_15120),
.B(n_14911),
.Y(n_15906)
);

OAI221xp5_ASAP7_75t_L g15907 ( 
.A1(n_15213),
.A2(n_14730),
.B1(n_14900),
.B2(n_14864),
.C(n_14660),
.Y(n_15907)
);

AND2x2_ASAP7_75t_L g15908 ( 
.A(n_15082),
.B(n_14926),
.Y(n_15908)
);

INVx1_ASAP7_75t_L g15909 ( 
.A(n_15122),
.Y(n_15909)
);

NAND2xp5_ASAP7_75t_L g15910 ( 
.A(n_15379),
.B(n_14955),
.Y(n_15910)
);

OAI221xp5_ASAP7_75t_SL g15911 ( 
.A1(n_15646),
.A2(n_14627),
.B1(n_14646),
.B2(n_14449),
.C(n_14824),
.Y(n_15911)
);

NAND3xp33_ASAP7_75t_L g15912 ( 
.A(n_15816),
.B(n_14764),
.C(n_14930),
.Y(n_15912)
);

OA211x2_ASAP7_75t_L g15913 ( 
.A1(n_15654),
.A2(n_14603),
.B(n_14598),
.C(n_14746),
.Y(n_15913)
);

AOI22xp33_ASAP7_75t_L g15914 ( 
.A1(n_15619),
.A2(n_14428),
.B1(n_11627),
.B2(n_14453),
.Y(n_15914)
);

NAND3xp33_ASAP7_75t_L g15915 ( 
.A(n_15073),
.B(n_14939),
.C(n_14946),
.Y(n_15915)
);

NAND2xp5_ASAP7_75t_L g15916 ( 
.A(n_15487),
.B(n_14701),
.Y(n_15916)
);

NAND2xp5_ASAP7_75t_SL g15917 ( 
.A(n_15197),
.B(n_14766),
.Y(n_15917)
);

OAI22xp5_ASAP7_75t_L g15918 ( 
.A1(n_15730),
.A2(n_14760),
.B1(n_14741),
.B2(n_9838),
.Y(n_15918)
);

AND2x2_ASAP7_75t_L g15919 ( 
.A(n_15066),
.B(n_14739),
.Y(n_15919)
);

NOR2xp33_ASAP7_75t_L g15920 ( 
.A(n_15005),
.B(n_14595),
.Y(n_15920)
);

NAND4xp25_ASAP7_75t_L g15921 ( 
.A(n_15008),
.B(n_14850),
.C(n_14631),
.D(n_14625),
.Y(n_15921)
);

NAND2xp5_ASAP7_75t_L g15922 ( 
.A(n_15497),
.B(n_14614),
.Y(n_15922)
);

NAND2xp33_ASAP7_75t_SL g15923 ( 
.A(n_15730),
.B(n_10711),
.Y(n_15923)
);

NAND3xp33_ASAP7_75t_L g15924 ( 
.A(n_15073),
.B(n_14981),
.C(n_14812),
.Y(n_15924)
);

AND2x2_ASAP7_75t_L g15925 ( 
.A(n_15066),
.B(n_14727),
.Y(n_15925)
);

AND2x2_ASAP7_75t_L g15926 ( 
.A(n_15059),
.B(n_14749),
.Y(n_15926)
);

AND2x2_ASAP7_75t_L g15927 ( 
.A(n_15140),
.B(n_15219),
.Y(n_15927)
);

AOI22xp33_ASAP7_75t_SL g15928 ( 
.A1(n_15738),
.A2(n_14600),
.B1(n_14989),
.B2(n_14665),
.Y(n_15928)
);

NAND3xp33_ASAP7_75t_L g15929 ( 
.A(n_15382),
.B(n_14775),
.C(n_14893),
.Y(n_15929)
);

NAND2xp5_ASAP7_75t_L g15930 ( 
.A(n_15071),
.B(n_14906),
.Y(n_15930)
);

NOR2xp33_ASAP7_75t_R g15931 ( 
.A(n_15171),
.B(n_15138),
.Y(n_15931)
);

NAND3xp33_ASAP7_75t_L g15932 ( 
.A(n_15738),
.B(n_14480),
.C(n_14476),
.Y(n_15932)
);

NAND2xp5_ASAP7_75t_L g15933 ( 
.A(n_15004),
.B(n_14781),
.Y(n_15933)
);

NAND3xp33_ASAP7_75t_L g15934 ( 
.A(n_15846),
.B(n_14551),
.C(n_14656),
.Y(n_15934)
);

NAND2xp5_ASAP7_75t_SL g15935 ( 
.A(n_15701),
.B(n_14709),
.Y(n_15935)
);

INVx1_ASAP7_75t_L g15936 ( 
.A(n_15124),
.Y(n_15936)
);

AND2x2_ASAP7_75t_L g15937 ( 
.A(n_15265),
.B(n_15079),
.Y(n_15937)
);

NAND2xp5_ASAP7_75t_L g15938 ( 
.A(n_15222),
.B(n_14960),
.Y(n_15938)
);

AOI22xp33_ASAP7_75t_SL g15939 ( 
.A1(n_15862),
.A2(n_14973),
.B1(n_14794),
.B2(n_14890),
.Y(n_15939)
);

OAI22xp5_ASAP7_75t_L g15940 ( 
.A1(n_15193),
.A2(n_9838),
.B1(n_9892),
.B2(n_9872),
.Y(n_15940)
);

AOI221xp5_ASAP7_75t_L g15941 ( 
.A1(n_15068),
.A2(n_14622),
.B1(n_14615),
.B2(n_14538),
.C(n_14510),
.Y(n_15941)
);

NAND3xp33_ASAP7_75t_L g15942 ( 
.A(n_15481),
.B(n_14685),
.C(n_14656),
.Y(n_15942)
);

OAI22xp5_ASAP7_75t_L g15943 ( 
.A1(n_15560),
.A2(n_9872),
.B1(n_9941),
.B2(n_9911),
.Y(n_15943)
);

OAI221xp5_ASAP7_75t_L g15944 ( 
.A1(n_15085),
.A2(n_14399),
.B1(n_14445),
.B2(n_14392),
.C(n_14385),
.Y(n_15944)
);

INVx2_ASAP7_75t_L g15945 ( 
.A(n_15150),
.Y(n_15945)
);

AND2x2_ASAP7_75t_L g15946 ( 
.A(n_15220),
.B(n_14749),
.Y(n_15946)
);

OA211x2_ASAP7_75t_L g15947 ( 
.A1(n_15007),
.A2(n_14757),
.B(n_14830),
.C(n_14540),
.Y(n_15947)
);

AND2x2_ASAP7_75t_L g15948 ( 
.A(n_15252),
.B(n_14539),
.Y(n_15948)
);

NAND2xp5_ASAP7_75t_L g15949 ( 
.A(n_15058),
.B(n_15000),
.Y(n_15949)
);

NAND2xp5_ASAP7_75t_L g15950 ( 
.A(n_15188),
.B(n_14999),
.Y(n_15950)
);

AND2x2_ASAP7_75t_SL g15951 ( 
.A(n_15374),
.B(n_11463),
.Y(n_15951)
);

INVx1_ASAP7_75t_L g15952 ( 
.A(n_15028),
.Y(n_15952)
);

AND2x2_ASAP7_75t_L g15953 ( 
.A(n_15432),
.B(n_14539),
.Y(n_15953)
);

NAND2xp5_ASAP7_75t_L g15954 ( 
.A(n_15168),
.B(n_14653),
.Y(n_15954)
);

OAI21xp33_ASAP7_75t_SL g15955 ( 
.A1(n_15092),
.A2(n_14792),
.B(n_14929),
.Y(n_15955)
);

NAND2xp5_ASAP7_75t_L g15956 ( 
.A(n_15185),
.B(n_14704),
.Y(n_15956)
);

AND2x2_ASAP7_75t_L g15957 ( 
.A(n_15095),
.B(n_14386),
.Y(n_15957)
);

NAND2xp5_ASAP7_75t_SL g15958 ( 
.A(n_15701),
.B(n_14801),
.Y(n_15958)
);

NAND3xp33_ASAP7_75t_L g15959 ( 
.A(n_15806),
.B(n_14702),
.C(n_14685),
.Y(n_15959)
);

NAND2xp5_ASAP7_75t_L g15960 ( 
.A(n_15189),
.B(n_15030),
.Y(n_15960)
);

OR2x2_ASAP7_75t_L g15961 ( 
.A(n_15006),
.B(n_14914),
.Y(n_15961)
);

AOI221xp5_ASAP7_75t_L g15962 ( 
.A1(n_15753),
.A2(n_14535),
.B1(n_14589),
.B2(n_14717),
.C(n_14979),
.Y(n_15962)
);

NAND2xp5_ASAP7_75t_L g15963 ( 
.A(n_15254),
.B(n_14953),
.Y(n_15963)
);

NAND2xp5_ASAP7_75t_L g15964 ( 
.A(n_15254),
.B(n_14983),
.Y(n_15964)
);

NAND2xp5_ASAP7_75t_L g15965 ( 
.A(n_15010),
.B(n_14863),
.Y(n_15965)
);

NAND2xp5_ASAP7_75t_L g15966 ( 
.A(n_15115),
.B(n_14879),
.Y(n_15966)
);

AND2x2_ASAP7_75t_L g15967 ( 
.A(n_15302),
.B(n_14386),
.Y(n_15967)
);

AND2x2_ASAP7_75t_L g15968 ( 
.A(n_15257),
.B(n_14905),
.Y(n_15968)
);

AND2x2_ASAP7_75t_L g15969 ( 
.A(n_15105),
.B(n_14728),
.Y(n_15969)
);

AND2x2_ASAP7_75t_L g15970 ( 
.A(n_15113),
.B(n_14728),
.Y(n_15970)
);

NAND2xp5_ASAP7_75t_L g15971 ( 
.A(n_15115),
.B(n_13931),
.Y(n_15971)
);

AND2x2_ASAP7_75t_L g15972 ( 
.A(n_15261),
.B(n_14621),
.Y(n_15972)
);

NAND2xp5_ASAP7_75t_L g15973 ( 
.A(n_15036),
.B(n_13932),
.Y(n_15973)
);

NAND2xp5_ASAP7_75t_L g15974 ( 
.A(n_15051),
.B(n_13935),
.Y(n_15974)
);

NAND2xp5_ASAP7_75t_L g15975 ( 
.A(n_15057),
.B(n_13939),
.Y(n_15975)
);

NAND2xp5_ASAP7_75t_L g15976 ( 
.A(n_15564),
.B(n_13945),
.Y(n_15976)
);

NAND4xp25_ASAP7_75t_L g15977 ( 
.A(n_15170),
.B(n_14579),
.C(n_14482),
.D(n_14659),
.Y(n_15977)
);

AND2x2_ASAP7_75t_L g15978 ( 
.A(n_15089),
.B(n_14621),
.Y(n_15978)
);

NAND2xp5_ASAP7_75t_L g15979 ( 
.A(n_15018),
.B(n_15039),
.Y(n_15979)
);

OAI221xp5_ASAP7_75t_SL g15980 ( 
.A1(n_15458),
.A2(n_14790),
.B1(n_14817),
.B2(n_14808),
.C(n_14679),
.Y(n_15980)
);

AND2x2_ASAP7_75t_L g15981 ( 
.A(n_15204),
.B(n_14679),
.Y(n_15981)
);

OAI221xp5_ASAP7_75t_L g15982 ( 
.A1(n_15752),
.A2(n_14521),
.B1(n_14681),
.B2(n_14849),
.C(n_14522),
.Y(n_15982)
);

NAND2xp5_ASAP7_75t_L g15983 ( 
.A(n_15091),
.B(n_13946),
.Y(n_15983)
);

AOI21xp5_ASAP7_75t_L g15984 ( 
.A1(n_15594),
.A2(n_14751),
.B(n_14441),
.Y(n_15984)
);

NAND2xp5_ASAP7_75t_L g15985 ( 
.A(n_15093),
.B(n_13950),
.Y(n_15985)
);

NAND2xp5_ASAP7_75t_L g15986 ( 
.A(n_15417),
.B(n_13954),
.Y(n_15986)
);

AND2x2_ASAP7_75t_L g15987 ( 
.A(n_15111),
.B(n_10547),
.Y(n_15987)
);

NAND2x1_ASAP7_75t_L g15988 ( 
.A(n_15477),
.B(n_14507),
.Y(n_15988)
);

AND2x2_ASAP7_75t_L g15989 ( 
.A(n_15264),
.B(n_10547),
.Y(n_15989)
);

NAND2xp5_ASAP7_75t_L g15990 ( 
.A(n_15417),
.B(n_13955),
.Y(n_15990)
);

AOI21xp33_ASAP7_75t_L g15991 ( 
.A1(n_15596),
.A2(n_14702),
.B(n_11520),
.Y(n_15991)
);

OAI221xp5_ASAP7_75t_SL g15992 ( 
.A1(n_15414),
.A2(n_15239),
.B1(n_15354),
.B2(n_15644),
.C(n_15283),
.Y(n_15992)
);

AND2x2_ASAP7_75t_L g15993 ( 
.A(n_15052),
.B(n_15041),
.Y(n_15993)
);

NAND2xp5_ASAP7_75t_SL g15994 ( 
.A(n_15374),
.B(n_15206),
.Y(n_15994)
);

NAND2xp5_ASAP7_75t_L g15995 ( 
.A(n_15206),
.B(n_13960),
.Y(n_15995)
);

NAND2xp5_ASAP7_75t_L g15996 ( 
.A(n_15117),
.B(n_9086),
.Y(n_15996)
);

NAND2xp5_ASAP7_75t_SL g15997 ( 
.A(n_15868),
.B(n_10711),
.Y(n_15997)
);

BUFx3_ASAP7_75t_L g15998 ( 
.A(n_15138),
.Y(n_15998)
);

AND2x2_ASAP7_75t_L g15999 ( 
.A(n_15052),
.B(n_10547),
.Y(n_15999)
);

NAND2xp5_ASAP7_75t_L g16000 ( 
.A(n_15125),
.B(n_15148),
.Y(n_16000)
);

OAI22xp5_ASAP7_75t_L g16001 ( 
.A1(n_15657),
.A2(n_9911),
.B1(n_9954),
.B2(n_9941),
.Y(n_16001)
);

NAND3xp33_ASAP7_75t_L g16002 ( 
.A(n_15806),
.B(n_14873),
.C(n_14872),
.Y(n_16002)
);

AND2x2_ASAP7_75t_L g16003 ( 
.A(n_15045),
.B(n_15048),
.Y(n_16003)
);

NAND2xp5_ASAP7_75t_L g16004 ( 
.A(n_15153),
.B(n_9086),
.Y(n_16004)
);

NAND3xp33_ASAP7_75t_L g16005 ( 
.A(n_15835),
.B(n_13282),
.C(n_13232),
.Y(n_16005)
);

AND2x2_ASAP7_75t_L g16006 ( 
.A(n_15395),
.B(n_14529),
.Y(n_16006)
);

HB1xp67_ASAP7_75t_L g16007 ( 
.A(n_15742),
.Y(n_16007)
);

NAND2xp5_ASAP7_75t_L g16008 ( 
.A(n_15158),
.B(n_9086),
.Y(n_16008)
);

NAND2xp5_ASAP7_75t_L g16009 ( 
.A(n_15358),
.B(n_15363),
.Y(n_16009)
);

INVxp67_ASAP7_75t_L g16010 ( 
.A(n_15021),
.Y(n_16010)
);

AND2x2_ASAP7_75t_SL g16011 ( 
.A(n_15835),
.B(n_11463),
.Y(n_16011)
);

NAND3xp33_ASAP7_75t_L g16012 ( 
.A(n_15836),
.B(n_13282),
.C(n_13232),
.Y(n_16012)
);

NAND2xp5_ASAP7_75t_L g16013 ( 
.A(n_15246),
.B(n_9086),
.Y(n_16013)
);

NAND3xp33_ASAP7_75t_L g16014 ( 
.A(n_15836),
.B(n_15151),
.C(n_15595),
.Y(n_16014)
);

NAND2xp5_ASAP7_75t_L g16015 ( 
.A(n_15029),
.B(n_15031),
.Y(n_16015)
);

NAND3xp33_ASAP7_75t_L g16016 ( 
.A(n_15595),
.B(n_13370),
.C(n_13650),
.Y(n_16016)
);

NAND2xp5_ASAP7_75t_L g16017 ( 
.A(n_15037),
.B(n_9086),
.Y(n_16017)
);

OAI21xp33_ASAP7_75t_L g16018 ( 
.A1(n_15565),
.A2(n_10461),
.B(n_11130),
.Y(n_16018)
);

AOI22xp33_ASAP7_75t_L g16019 ( 
.A1(n_15856),
.A2(n_11627),
.B1(n_10766),
.B2(n_10879),
.Y(n_16019)
);

NAND3xp33_ASAP7_75t_L g16020 ( 
.A(n_15728),
.B(n_13672),
.C(n_13650),
.Y(n_16020)
);

NAND2xp5_ASAP7_75t_L g16021 ( 
.A(n_15042),
.B(n_9090),
.Y(n_16021)
);

NAND2xp5_ASAP7_75t_L g16022 ( 
.A(n_15402),
.B(n_9090),
.Y(n_16022)
);

NAND2xp5_ASAP7_75t_L g16023 ( 
.A(n_15402),
.B(n_9090),
.Y(n_16023)
);

INVx2_ASAP7_75t_L g16024 ( 
.A(n_15150),
.Y(n_16024)
);

NAND3xp33_ASAP7_75t_L g16025 ( 
.A(n_15728),
.B(n_13690),
.C(n_13672),
.Y(n_16025)
);

AND2x2_ASAP7_75t_L g16026 ( 
.A(n_15396),
.B(n_14529),
.Y(n_16026)
);

OA21x2_ASAP7_75t_L g16027 ( 
.A1(n_15028),
.A2(n_14383),
.B(n_13711),
.Y(n_16027)
);

OAI21xp33_ASAP7_75t_L g16028 ( 
.A1(n_15062),
.A2(n_10461),
.B(n_11130),
.Y(n_16028)
);

NAND2xp5_ASAP7_75t_L g16029 ( 
.A(n_15466),
.B(n_9090),
.Y(n_16029)
);

AOI221xp5_ASAP7_75t_L g16030 ( 
.A1(n_15742),
.A2(n_14998),
.B1(n_14668),
.B2(n_14613),
.C(n_14506),
.Y(n_16030)
);

NAND3xp33_ASAP7_75t_L g16031 ( 
.A(n_15354),
.B(n_13711),
.C(n_13690),
.Y(n_16031)
);

NAND2xp5_ASAP7_75t_SL g16032 ( 
.A(n_15372),
.B(n_10711),
.Y(n_16032)
);

AND2x2_ASAP7_75t_L g16033 ( 
.A(n_15214),
.B(n_11336),
.Y(n_16033)
);

OA21x2_ASAP7_75t_L g16034 ( 
.A1(n_15791),
.A2(n_13744),
.B(n_13738),
.Y(n_16034)
);

AOI22xp33_ASAP7_75t_L g16035 ( 
.A1(n_15359),
.A2(n_10766),
.B1(n_10879),
.B2(n_10896),
.Y(n_16035)
);

NOR2xp33_ASAP7_75t_L g16036 ( 
.A(n_15099),
.B(n_11463),
.Y(n_16036)
);

AND2x2_ASAP7_75t_L g16037 ( 
.A(n_15101),
.B(n_11336),
.Y(n_16037)
);

AOI21xp5_ASAP7_75t_SL g16038 ( 
.A1(n_15110),
.A2(n_13952),
.B(n_13990),
.Y(n_16038)
);

NAND3xp33_ASAP7_75t_L g16039 ( 
.A(n_15301),
.B(n_13744),
.C(n_13738),
.Y(n_16039)
);

AND2x2_ASAP7_75t_L g16040 ( 
.A(n_15063),
.B(n_11336),
.Y(n_16040)
);

OAI221xp5_ASAP7_75t_SL g16041 ( 
.A1(n_15366),
.A2(n_10461),
.B1(n_14643),
.B2(n_9397),
.C(n_9308),
.Y(n_16041)
);

NAND3xp33_ASAP7_75t_L g16042 ( 
.A(n_15791),
.B(n_13753),
.C(n_10766),
.Y(n_16042)
);

AND2x2_ASAP7_75t_L g16043 ( 
.A(n_15083),
.B(n_15088),
.Y(n_16043)
);

NAND3xp33_ASAP7_75t_L g16044 ( 
.A(n_15606),
.B(n_13753),
.C(n_10766),
.Y(n_16044)
);

AND2x2_ASAP7_75t_L g16045 ( 
.A(n_15687),
.B(n_15014),
.Y(n_16045)
);

NAND2xp5_ASAP7_75t_L g16046 ( 
.A(n_15472),
.B(n_9090),
.Y(n_16046)
);

OAI21xp5_ASAP7_75t_SL g16047 ( 
.A1(n_15338),
.A2(n_10893),
.B(n_10892),
.Y(n_16047)
);

NOR3xp33_ASAP7_75t_L g16048 ( 
.A(n_15365),
.B(n_14454),
.C(n_13969),
.Y(n_16048)
);

AOI22xp33_ASAP7_75t_L g16049 ( 
.A1(n_15369),
.A2(n_10766),
.B1(n_10879),
.B2(n_10896),
.Y(n_16049)
);

NAND2xp5_ASAP7_75t_L g16050 ( 
.A(n_15475),
.B(n_15480),
.Y(n_16050)
);

AND2x2_ASAP7_75t_L g16051 ( 
.A(n_15096),
.B(n_11342),
.Y(n_16051)
);

NAND2xp5_ASAP7_75t_L g16052 ( 
.A(n_15486),
.B(n_9097),
.Y(n_16052)
);

NAND3xp33_ASAP7_75t_L g16053 ( 
.A(n_15313),
.B(n_15179),
.C(n_15706),
.Y(n_16053)
);

OAI21xp5_ASAP7_75t_L g16054 ( 
.A1(n_15865),
.A2(n_15602),
.B(n_15863),
.Y(n_16054)
);

NAND2xp5_ASAP7_75t_L g16055 ( 
.A(n_15489),
.B(n_9097),
.Y(n_16055)
);

NAND2xp5_ASAP7_75t_L g16056 ( 
.A(n_15502),
.B(n_9097),
.Y(n_16056)
);

NOR3xp33_ASAP7_75t_L g16057 ( 
.A(n_15416),
.B(n_13969),
.C(n_13964),
.Y(n_16057)
);

OAI221xp5_ASAP7_75t_SL g16058 ( 
.A1(n_15418),
.A2(n_10461),
.B1(n_14643),
.B2(n_9308),
.C(n_9397),
.Y(n_16058)
);

NAND3xp33_ASAP7_75t_L g16059 ( 
.A(n_15592),
.B(n_10896),
.C(n_10874),
.Y(n_16059)
);

NAND2xp5_ASAP7_75t_L g16060 ( 
.A(n_15514),
.B(n_9097),
.Y(n_16060)
);

OAI22xp5_ASAP7_75t_L g16061 ( 
.A1(n_15053),
.A2(n_9941),
.B1(n_9954),
.B2(n_9911),
.Y(n_16061)
);

AND2x2_ASAP7_75t_L g16062 ( 
.A(n_15096),
.B(n_11342),
.Y(n_16062)
);

NAND2xp5_ASAP7_75t_L g16063 ( 
.A(n_15519),
.B(n_9097),
.Y(n_16063)
);

OAI22xp5_ASAP7_75t_L g16064 ( 
.A1(n_15297),
.A2(n_9941),
.B1(n_9954),
.B2(n_9911),
.Y(n_16064)
);

OA21x2_ASAP7_75t_L g16065 ( 
.A1(n_15401),
.A2(n_13979),
.B(n_13964),
.Y(n_16065)
);

AND2x2_ASAP7_75t_L g16066 ( 
.A(n_15017),
.B(n_15198),
.Y(n_16066)
);

NAND2xp5_ASAP7_75t_L g16067 ( 
.A(n_15536),
.B(n_9097),
.Y(n_16067)
);

AND2x2_ASAP7_75t_L g16068 ( 
.A(n_15044),
.B(n_11342),
.Y(n_16068)
);

NAND2xp5_ASAP7_75t_L g16069 ( 
.A(n_15540),
.B(n_9125),
.Y(n_16069)
);

NAND2xp5_ASAP7_75t_L g16070 ( 
.A(n_15218),
.B(n_9125),
.Y(n_16070)
);

NAND2xp5_ASAP7_75t_SL g16071 ( 
.A(n_15372),
.B(n_10711),
.Y(n_16071)
);

OAI21xp5_ASAP7_75t_L g16072 ( 
.A1(n_15247),
.A2(n_10781),
.B(n_13952),
.Y(n_16072)
);

NAND2xp5_ASAP7_75t_L g16073 ( 
.A(n_15218),
.B(n_9125),
.Y(n_16073)
);

AND2x2_ASAP7_75t_L g16074 ( 
.A(n_15231),
.B(n_11374),
.Y(n_16074)
);

NAND2xp5_ASAP7_75t_SL g16075 ( 
.A(n_15378),
.B(n_10711),
.Y(n_16075)
);

INVx1_ASAP7_75t_L g16076 ( 
.A(n_15309),
.Y(n_16076)
);

NOR2xp33_ASAP7_75t_L g16077 ( 
.A(n_15378),
.B(n_15404),
.Y(n_16077)
);

NAND2xp5_ASAP7_75t_L g16078 ( 
.A(n_15055),
.B(n_9125),
.Y(n_16078)
);

AND2x2_ASAP7_75t_L g16079 ( 
.A(n_15069),
.B(n_11374),
.Y(n_16079)
);

OAI22xp5_ASAP7_75t_L g16080 ( 
.A1(n_15655),
.A2(n_9911),
.B1(n_9954),
.B2(n_9941),
.Y(n_16080)
);

AOI22xp33_ASAP7_75t_L g16081 ( 
.A1(n_15795),
.A2(n_10879),
.B1(n_10896),
.B2(n_10874),
.Y(n_16081)
);

OA21x2_ASAP7_75t_L g16082 ( 
.A1(n_15401),
.A2(n_13988),
.B(n_13979),
.Y(n_16082)
);

NAND2xp5_ASAP7_75t_L g16083 ( 
.A(n_15060),
.B(n_9125),
.Y(n_16083)
);

NAND4xp25_ASAP7_75t_L g16084 ( 
.A(n_15279),
.B(n_10063),
.C(n_9448),
.D(n_9677),
.Y(n_16084)
);

NAND3xp33_ASAP7_75t_L g16085 ( 
.A(n_15592),
.B(n_10896),
.C(n_10874),
.Y(n_16085)
);

OAI22xp5_ASAP7_75t_L g16086 ( 
.A1(n_15268),
.A2(n_9911),
.B1(n_9954),
.B2(n_9941),
.Y(n_16086)
);

NOR3xp33_ASAP7_75t_L g16087 ( 
.A(n_15210),
.B(n_13988),
.C(n_10381),
.Y(n_16087)
);

OAI21xp33_ASAP7_75t_L g16088 ( 
.A1(n_15840),
.A2(n_10461),
.B(n_11130),
.Y(n_16088)
);

NAND2xp5_ASAP7_75t_L g16089 ( 
.A(n_15061),
.B(n_9125),
.Y(n_16089)
);

OA211x2_ASAP7_75t_L g16090 ( 
.A1(n_15102),
.A2(n_9335),
.B(n_9249),
.C(n_9870),
.Y(n_16090)
);

NOR3xp33_ASAP7_75t_SL g16091 ( 
.A(n_15588),
.B(n_9697),
.C(n_11520),
.Y(n_16091)
);

NAND2xp5_ASAP7_75t_L g16092 ( 
.A(n_15064),
.B(n_11130),
.Y(n_16092)
);

NAND4xp25_ASAP7_75t_L g16093 ( 
.A(n_15537),
.B(n_10063),
.C(n_9351),
.D(n_9677),
.Y(n_16093)
);

OAI221xp5_ASAP7_75t_SL g16094 ( 
.A1(n_15857),
.A2(n_10461),
.B1(n_9397),
.B2(n_9308),
.C(n_9231),
.Y(n_16094)
);

INVxp67_ASAP7_75t_L g16095 ( 
.A(n_15839),
.Y(n_16095)
);

AOI22xp33_ASAP7_75t_L g16096 ( 
.A1(n_15697),
.A2(n_15850),
.B1(n_15852),
.B2(n_15637),
.Y(n_16096)
);

NAND2xp5_ASAP7_75t_L g16097 ( 
.A(n_15065),
.B(n_11130),
.Y(n_16097)
);

NAND3xp33_ASAP7_75t_L g16098 ( 
.A(n_15172),
.B(n_10874),
.C(n_10804),
.Y(n_16098)
);

AOI22xp33_ASAP7_75t_SL g16099 ( 
.A1(n_15233),
.A2(n_9941),
.B1(n_9954),
.B2(n_9911),
.Y(n_16099)
);

NAND3xp33_ASAP7_75t_L g16100 ( 
.A(n_15653),
.B(n_15826),
.C(n_15413),
.Y(n_16100)
);

NAND4xp25_ASAP7_75t_L g16101 ( 
.A(n_15607),
.B(n_10063),
.C(n_9351),
.D(n_9677),
.Y(n_16101)
);

NOR2xp33_ASAP7_75t_L g16102 ( 
.A(n_15224),
.B(n_15429),
.Y(n_16102)
);

OAI21xp5_ASAP7_75t_SL g16103 ( 
.A1(n_15177),
.A2(n_15682),
.B(n_15686),
.Y(n_16103)
);

NAND2xp5_ASAP7_75t_SL g16104 ( 
.A(n_15647),
.B(n_10753),
.Y(n_16104)
);

INVx2_ASAP7_75t_L g16105 ( 
.A(n_15150),
.Y(n_16105)
);

NOR3xp33_ASAP7_75t_L g16106 ( 
.A(n_15543),
.B(n_10381),
.C(n_10314),
.Y(n_16106)
);

NOR2xp33_ASAP7_75t_SL g16107 ( 
.A(n_15567),
.B(n_11520),
.Y(n_16107)
);

NAND2xp5_ASAP7_75t_L g16108 ( 
.A(n_15430),
.B(n_11130),
.Y(n_16108)
);

NAND2xp5_ASAP7_75t_L g16109 ( 
.A(n_15439),
.B(n_10643),
.Y(n_16109)
);

NAND3xp33_ASAP7_75t_L g16110 ( 
.A(n_15413),
.B(n_10874),
.C(n_10804),
.Y(n_16110)
);

NAND2xp5_ASAP7_75t_L g16111 ( 
.A(n_15131),
.B(n_10643),
.Y(n_16111)
);

AND2x2_ASAP7_75t_L g16112 ( 
.A(n_15319),
.B(n_11374),
.Y(n_16112)
);

OAI22xp5_ASAP7_75t_L g16113 ( 
.A1(n_15500),
.A2(n_9911),
.B1(n_9954),
.B2(n_9941),
.Y(n_16113)
);

NOR2xp33_ASAP7_75t_L g16114 ( 
.A(n_15546),
.B(n_11520),
.Y(n_16114)
);

AND2x2_ASAP7_75t_L g16115 ( 
.A(n_15033),
.B(n_11386),
.Y(n_16115)
);

OAI221xp5_ASAP7_75t_SL g16116 ( 
.A1(n_15786),
.A2(n_9397),
.B1(n_9308),
.B2(n_10307),
.C(n_10304),
.Y(n_16116)
);

AND2x2_ASAP7_75t_L g16117 ( 
.A(n_15033),
.B(n_11386),
.Y(n_16117)
);

NAND3xp33_ASAP7_75t_L g16118 ( 
.A(n_15600),
.B(n_10874),
.C(n_10804),
.Y(n_16118)
);

AND2x2_ASAP7_75t_L g16119 ( 
.A(n_15129),
.B(n_11386),
.Y(n_16119)
);

OAI221xp5_ASAP7_75t_L g16120 ( 
.A1(n_15617),
.A2(n_10972),
.B1(n_11028),
.B2(n_10893),
.C(n_10892),
.Y(n_16120)
);

AND2x2_ASAP7_75t_L g16121 ( 
.A(n_15324),
.B(n_11389),
.Y(n_16121)
);

NAND4xp25_ASAP7_75t_L g16122 ( 
.A(n_15615),
.B(n_10063),
.C(n_9351),
.D(n_9677),
.Y(n_16122)
);

OAI22xp5_ASAP7_75t_L g16123 ( 
.A1(n_15808),
.A2(n_15304),
.B1(n_15251),
.B2(n_15483),
.Y(n_16123)
);

OAI21xp33_ASAP7_75t_SL g16124 ( 
.A1(n_15130),
.A2(n_14909),
.B(n_14932),
.Y(n_16124)
);

NOR2x1_ASAP7_75t_L g16125 ( 
.A(n_15043),
.B(n_14784),
.Y(n_16125)
);

AND2x2_ASAP7_75t_L g16126 ( 
.A(n_15583),
.B(n_11389),
.Y(n_16126)
);

NAND2xp5_ASAP7_75t_L g16127 ( 
.A(n_15639),
.B(n_10643),
.Y(n_16127)
);

AND2x2_ASAP7_75t_L g16128 ( 
.A(n_15155),
.B(n_11389),
.Y(n_16128)
);

NAND3xp33_ASAP7_75t_L g16129 ( 
.A(n_15364),
.B(n_10804),
.C(n_10791),
.Y(n_16129)
);

OAI21xp5_ASAP7_75t_L g16130 ( 
.A1(n_15649),
.A2(n_10781),
.B(n_10804),
.Y(n_16130)
);

AOI22xp33_ASAP7_75t_SL g16131 ( 
.A1(n_15790),
.A2(n_9941),
.B1(n_9954),
.B2(n_9911),
.Y(n_16131)
);

AND2x2_ASAP7_75t_L g16132 ( 
.A(n_15156),
.B(n_11400),
.Y(n_16132)
);

AND2x2_ASAP7_75t_L g16133 ( 
.A(n_15612),
.B(n_11400),
.Y(n_16133)
);

OAI22xp5_ASAP7_75t_L g16134 ( 
.A1(n_15304),
.A2(n_9911),
.B1(n_9954),
.B2(n_9941),
.Y(n_16134)
);

AND2x2_ASAP7_75t_L g16135 ( 
.A(n_15116),
.B(n_11400),
.Y(n_16135)
);

AND2x2_ASAP7_75t_L g16136 ( 
.A(n_15190),
.B(n_11404),
.Y(n_16136)
);

AOI22xp33_ASAP7_75t_L g16137 ( 
.A1(n_15546),
.A2(n_10791),
.B1(n_10513),
.B2(n_10718),
.Y(n_16137)
);

AND2x2_ASAP7_75t_L g16138 ( 
.A(n_15181),
.B(n_11404),
.Y(n_16138)
);

NAND2xp5_ASAP7_75t_L g16139 ( 
.A(n_15641),
.B(n_10655),
.Y(n_16139)
);

AOI22xp33_ASAP7_75t_L g16140 ( 
.A1(n_15845),
.A2(n_10791),
.B1(n_10513),
.B2(n_10718),
.Y(n_16140)
);

NAND2xp5_ASAP7_75t_L g16141 ( 
.A(n_15663),
.B(n_10655),
.Y(n_16141)
);

AND2x2_ASAP7_75t_L g16142 ( 
.A(n_15479),
.B(n_11404),
.Y(n_16142)
);

NAND4xp25_ASAP7_75t_L g16143 ( 
.A(n_15050),
.B(n_10063),
.C(n_9351),
.D(n_9448),
.Y(n_16143)
);

NAND2xp5_ASAP7_75t_SL g16144 ( 
.A(n_15647),
.B(n_10753),
.Y(n_16144)
);

NAND2xp5_ASAP7_75t_L g16145 ( 
.A(n_15668),
.B(n_10655),
.Y(n_16145)
);

OAI21xp5_ASAP7_75t_SL g16146 ( 
.A1(n_15267),
.A2(n_11028),
.B(n_10972),
.Y(n_16146)
);

AOI22xp5_ASAP7_75t_L g16147 ( 
.A1(n_15633),
.A2(n_11520),
.B1(n_10159),
.B2(n_10137),
.Y(n_16147)
);

AND2x2_ASAP7_75t_L g16148 ( 
.A(n_15691),
.B(n_11458),
.Y(n_16148)
);

NAND2xp5_ASAP7_75t_L g16149 ( 
.A(n_15134),
.B(n_10737),
.Y(n_16149)
);

AND2x2_ASAP7_75t_L g16150 ( 
.A(n_15584),
.B(n_11458),
.Y(n_16150)
);

OAI221xp5_ASAP7_75t_SL g16151 ( 
.A1(n_15640),
.A2(n_9397),
.B1(n_10307),
.B2(n_10335),
.C(n_10304),
.Y(n_16151)
);

AND2x2_ASAP7_75t_L g16152 ( 
.A(n_15194),
.B(n_11458),
.Y(n_16152)
);

NAND2xp5_ASAP7_75t_L g16153 ( 
.A(n_15142),
.B(n_10737),
.Y(n_16153)
);

NAND2xp5_ASAP7_75t_L g16154 ( 
.A(n_15142),
.B(n_10737),
.Y(n_16154)
);

NAND4xp25_ASAP7_75t_L g16155 ( 
.A(n_15661),
.B(n_9448),
.C(n_9697),
.D(n_9531),
.Y(n_16155)
);

AOI21xp5_ASAP7_75t_L g16156 ( 
.A1(n_15230),
.A2(n_14751),
.B(n_14829),
.Y(n_16156)
);

AND2x2_ASAP7_75t_L g16157 ( 
.A(n_15383),
.B(n_10997),
.Y(n_16157)
);

NAND2xp5_ASAP7_75t_L g16158 ( 
.A(n_15114),
.B(n_10792),
.Y(n_16158)
);

OAI22x1_ASAP7_75t_L g16159 ( 
.A1(n_15269),
.A2(n_9563),
.B1(n_9848),
.B2(n_9675),
.Y(n_16159)
);

NAND2xp5_ASAP7_75t_L g16160 ( 
.A(n_15118),
.B(n_10792),
.Y(n_16160)
);

AND2x2_ASAP7_75t_L g16161 ( 
.A(n_15054),
.B(n_10997),
.Y(n_16161)
);

AND2x2_ASAP7_75t_L g16162 ( 
.A(n_15054),
.B(n_11018),
.Y(n_16162)
);

AND2x2_ASAP7_75t_L g16163 ( 
.A(n_15152),
.B(n_11018),
.Y(n_16163)
);

AND2x2_ASAP7_75t_L g16164 ( 
.A(n_15161),
.B(n_11020),
.Y(n_16164)
);

NOR3xp33_ASAP7_75t_L g16165 ( 
.A(n_15496),
.B(n_10381),
.C(n_10314),
.Y(n_16165)
);

OA21x2_ASAP7_75t_L g16166 ( 
.A1(n_15662),
.A2(n_10880),
.B(n_10860),
.Y(n_16166)
);

OAI22xp5_ASAP7_75t_L g16167 ( 
.A1(n_15205),
.A2(n_9941),
.B1(n_9967),
.B2(n_9954),
.Y(n_16167)
);

AND2x2_ASAP7_75t_L g16168 ( 
.A(n_15162),
.B(n_11020),
.Y(n_16168)
);

NAND2xp5_ASAP7_75t_L g16169 ( 
.A(n_15015),
.B(n_10792),
.Y(n_16169)
);

NAND2xp5_ASAP7_75t_L g16170 ( 
.A(n_15019),
.B(n_10904),
.Y(n_16170)
);

OA211x2_ASAP7_75t_L g16171 ( 
.A1(n_15326),
.A2(n_9335),
.B(n_9249),
.C(n_9870),
.Y(n_16171)
);

OR2x2_ASAP7_75t_L g16172 ( 
.A(n_15244),
.B(n_11025),
.Y(n_16172)
);

NAND2xp5_ASAP7_75t_L g16173 ( 
.A(n_15022),
.B(n_10904),
.Y(n_16173)
);

NAND2xp5_ASAP7_75t_L g16174 ( 
.A(n_15025),
.B(n_10904),
.Y(n_16174)
);

AND2x2_ASAP7_75t_L g16175 ( 
.A(n_15734),
.B(n_11025),
.Y(n_16175)
);

INVx2_ASAP7_75t_L g16176 ( 
.A(n_15202),
.Y(n_16176)
);

AND2x2_ASAP7_75t_L g16177 ( 
.A(n_15121),
.B(n_11027),
.Y(n_16177)
);

NOR2xp33_ASAP7_75t_SL g16178 ( 
.A(n_15202),
.B(n_11606),
.Y(n_16178)
);

NAND2xp33_ASAP7_75t_SL g16179 ( 
.A(n_15391),
.B(n_10753),
.Y(n_16179)
);

OAI221xp5_ASAP7_75t_L g16180 ( 
.A1(n_15340),
.A2(n_11183),
.B1(n_11227),
.B2(n_11028),
.C(n_10972),
.Y(n_16180)
);

OA21x2_ASAP7_75t_L g16181 ( 
.A1(n_15662),
.A2(n_10889),
.B(n_10880),
.Y(n_16181)
);

NAND2xp5_ASAP7_75t_L g16182 ( 
.A(n_15034),
.B(n_10926),
.Y(n_16182)
);

OAI21xp33_ASAP7_75t_SL g16183 ( 
.A1(n_15040),
.A2(n_14909),
.B(n_14932),
.Y(n_16183)
);

NAND2xp5_ASAP7_75t_L g16184 ( 
.A(n_15038),
.B(n_10926),
.Y(n_16184)
);

OAI21xp5_ASAP7_75t_SL g16185 ( 
.A1(n_15746),
.A2(n_11028),
.B(n_10972),
.Y(n_16185)
);

NAND3xp33_ASAP7_75t_L g16186 ( 
.A(n_15844),
.B(n_10791),
.C(n_13417),
.Y(n_16186)
);

OAI21xp5_ASAP7_75t_SL g16187 ( 
.A1(n_15445),
.A2(n_11227),
.B(n_11183),
.Y(n_16187)
);

NAND2xp5_ASAP7_75t_L g16188 ( 
.A(n_15163),
.B(n_10926),
.Y(n_16188)
);

NAND2xp5_ASAP7_75t_SL g16189 ( 
.A(n_15469),
.B(n_10753),
.Y(n_16189)
);

OAI21xp5_ASAP7_75t_L g16190 ( 
.A1(n_15106),
.A2(n_10781),
.B(n_13990),
.Y(n_16190)
);

OAI221xp5_ASAP7_75t_SL g16191 ( 
.A1(n_15387),
.A2(n_10348),
.B1(n_10444),
.B2(n_10335),
.C(n_10304),
.Y(n_16191)
);

AND2x2_ASAP7_75t_L g16192 ( 
.A(n_15084),
.B(n_11027),
.Y(n_16192)
);

NAND2xp5_ASAP7_75t_L g16193 ( 
.A(n_15180),
.B(n_10928),
.Y(n_16193)
);

NAND2xp5_ASAP7_75t_SL g16194 ( 
.A(n_15469),
.B(n_15557),
.Y(n_16194)
);

AND2x2_ASAP7_75t_L g16195 ( 
.A(n_15442),
.B(n_11032),
.Y(n_16195)
);

NAND2xp5_ASAP7_75t_SL g16196 ( 
.A(n_15557),
.B(n_10753),
.Y(n_16196)
);

NAND2xp5_ASAP7_75t_L g16197 ( 
.A(n_15184),
.B(n_10928),
.Y(n_16197)
);

OAI22xp5_ASAP7_75t_L g16198 ( 
.A1(n_15047),
.A2(n_9941),
.B1(n_9967),
.B2(n_9954),
.Y(n_16198)
);

AND2x2_ASAP7_75t_L g16199 ( 
.A(n_15444),
.B(n_11032),
.Y(n_16199)
);

NAND3xp33_ASAP7_75t_L g16200 ( 
.A(n_15507),
.B(n_15474),
.C(n_15450),
.Y(n_16200)
);

AND2x2_ASAP7_75t_L g16201 ( 
.A(n_15455),
.B(n_11035),
.Y(n_16201)
);

NAND2xp5_ASAP7_75t_L g16202 ( 
.A(n_15199),
.B(n_10928),
.Y(n_16202)
);

AND2x2_ASAP7_75t_L g16203 ( 
.A(n_15460),
.B(n_11035),
.Y(n_16203)
);

INVx2_ASAP7_75t_L g16204 ( 
.A(n_15202),
.Y(n_16204)
);

NAND3xp33_ASAP7_75t_L g16205 ( 
.A(n_15274),
.B(n_10791),
.C(n_10718),
.Y(n_16205)
);

NAND3xp33_ASAP7_75t_L g16206 ( 
.A(n_15693),
.B(n_10791),
.C(n_10718),
.Y(n_16206)
);

AOI22xp33_ASAP7_75t_L g16207 ( 
.A1(n_15488),
.A2(n_10513),
.B1(n_10718),
.B2(n_10709),
.Y(n_16207)
);

NAND2xp5_ASAP7_75t_L g16208 ( 
.A(n_15164),
.B(n_10929),
.Y(n_16208)
);

NAND2xp5_ASAP7_75t_L g16209 ( 
.A(n_15167),
.B(n_10929),
.Y(n_16209)
);

OAI221xp5_ASAP7_75t_SL g16210 ( 
.A1(n_15541),
.A2(n_10444),
.B1(n_10570),
.B2(n_10348),
.C(n_10335),
.Y(n_16210)
);

OAI21xp5_ASAP7_75t_L g16211 ( 
.A1(n_15027),
.A2(n_13944),
.B(n_13875),
.Y(n_16211)
);

NAND2xp5_ASAP7_75t_L g16212 ( 
.A(n_15226),
.B(n_15132),
.Y(n_16212)
);

AND2x2_ASAP7_75t_L g16213 ( 
.A(n_15462),
.B(n_11036),
.Y(n_16213)
);

AOI22xp33_ASAP7_75t_L g16214 ( 
.A1(n_15490),
.A2(n_10513),
.B1(n_10718),
.B2(n_10709),
.Y(n_16214)
);

NAND2xp5_ASAP7_75t_SL g16215 ( 
.A(n_15579),
.B(n_10753),
.Y(n_16215)
);

NAND2xp5_ASAP7_75t_L g16216 ( 
.A(n_15249),
.B(n_15256),
.Y(n_16216)
);

NAND2xp5_ASAP7_75t_L g16217 ( 
.A(n_15259),
.B(n_10929),
.Y(n_16217)
);

NAND3xp33_ASAP7_75t_L g16218 ( 
.A(n_15726),
.B(n_10740),
.C(n_10709),
.Y(n_16218)
);

AOI22xp5_ASAP7_75t_L g16219 ( 
.A1(n_15859),
.A2(n_10159),
.B1(n_10137),
.B2(n_9775),
.Y(n_16219)
);

NAND2xp5_ASAP7_75t_L g16220 ( 
.A(n_15260),
.B(n_11021),
.Y(n_16220)
);

NAND4xp25_ASAP7_75t_L g16221 ( 
.A(n_15677),
.B(n_9448),
.C(n_9697),
.D(n_9573),
.Y(n_16221)
);

NAND3xp33_ASAP7_75t_L g16222 ( 
.A(n_15814),
.B(n_10740),
.C(n_10709),
.Y(n_16222)
);

NAND3xp33_ASAP7_75t_L g16223 ( 
.A(n_15712),
.B(n_10740),
.C(n_10709),
.Y(n_16223)
);

OAI221xp5_ASAP7_75t_SL g16224 ( 
.A1(n_15699),
.A2(n_10570),
.B1(n_10572),
.B2(n_10444),
.C(n_10348),
.Y(n_16224)
);

OAI22xp5_ASAP7_75t_L g16225 ( 
.A1(n_15542),
.A2(n_9954),
.B1(n_10024),
.B2(n_9967),
.Y(n_16225)
);

AOI22xp33_ASAP7_75t_L g16226 ( 
.A1(n_15521),
.A2(n_10513),
.B1(n_10740),
.B2(n_10709),
.Y(n_16226)
);

NAND2xp5_ASAP7_75t_L g16227 ( 
.A(n_15175),
.B(n_11021),
.Y(n_16227)
);

AND2x2_ASAP7_75t_L g16228 ( 
.A(n_15797),
.B(n_11036),
.Y(n_16228)
);

NAND2xp5_ASAP7_75t_L g16229 ( 
.A(n_15493),
.B(n_11021),
.Y(n_16229)
);

AND2x2_ASAP7_75t_L g16230 ( 
.A(n_15266),
.B(n_11050),
.Y(n_16230)
);

AND2x2_ASAP7_75t_L g16231 ( 
.A(n_15288),
.B(n_11050),
.Y(n_16231)
);

NAND3xp33_ASAP7_75t_L g16232 ( 
.A(n_15671),
.B(n_10740),
.C(n_13875),
.Y(n_16232)
);

OAI221xp5_ASAP7_75t_SL g16233 ( 
.A1(n_15281),
.A2(n_10593),
.B1(n_10758),
.B2(n_10572),
.C(n_10570),
.Y(n_16233)
);

AND2x2_ASAP7_75t_L g16234 ( 
.A(n_15333),
.B(n_11061),
.Y(n_16234)
);

NAND2xp5_ASAP7_75t_L g16235 ( 
.A(n_15558),
.B(n_11070),
.Y(n_16235)
);

AOI22xp33_ASAP7_75t_SL g16236 ( 
.A1(n_15215),
.A2(n_9967),
.B1(n_10024),
.B2(n_9954),
.Y(n_16236)
);

NAND2xp5_ASAP7_75t_L g16237 ( 
.A(n_15559),
.B(n_11070),
.Y(n_16237)
);

INVx2_ASAP7_75t_L g16238 ( 
.A(n_15227),
.Y(n_16238)
);

NAND3xp33_ASAP7_75t_L g16239 ( 
.A(n_15011),
.B(n_15026),
.C(n_15020),
.Y(n_16239)
);

NAND2xp5_ASAP7_75t_L g16240 ( 
.A(n_15270),
.B(n_11070),
.Y(n_16240)
);

NAND2xp5_ASAP7_75t_SL g16241 ( 
.A(n_15579),
.B(n_10821),
.Y(n_16241)
);

AOI22xp33_ASAP7_75t_L g16242 ( 
.A1(n_15722),
.A2(n_10513),
.B1(n_10740),
.B2(n_10906),
.Y(n_16242)
);

AND2x2_ASAP7_75t_L g16243 ( 
.A(n_15412),
.B(n_11061),
.Y(n_16243)
);

NAND2xp5_ASAP7_75t_L g16244 ( 
.A(n_15270),
.B(n_15598),
.Y(n_16244)
);

NAND2xp5_ASAP7_75t_L g16245 ( 
.A(n_15250),
.B(n_11064),
.Y(n_16245)
);

AND2x2_ASAP7_75t_L g16246 ( 
.A(n_15160),
.B(n_11064),
.Y(n_16246)
);

AND2x2_ASAP7_75t_L g16247 ( 
.A(n_15494),
.B(n_11068),
.Y(n_16247)
);

INVx2_ASAP7_75t_L g16248 ( 
.A(n_15046),
.Y(n_16248)
);

NAND2xp5_ASAP7_75t_SL g16249 ( 
.A(n_15344),
.B(n_10821),
.Y(n_16249)
);

AND2x2_ASAP7_75t_L g16250 ( 
.A(n_15508),
.B(n_11068),
.Y(n_16250)
);

NAND3xp33_ASAP7_75t_L g16251 ( 
.A(n_15207),
.B(n_13944),
.C(n_12077),
.Y(n_16251)
);

AND2x2_ASAP7_75t_L g16252 ( 
.A(n_15371),
.B(n_15373),
.Y(n_16252)
);

NAND2xp5_ASAP7_75t_L g16253 ( 
.A(n_15200),
.B(n_11078),
.Y(n_16253)
);

OAI221xp5_ASAP7_75t_SL g16254 ( 
.A1(n_15866),
.A2(n_10758),
.B1(n_10814),
.B2(n_10593),
.C(n_10572),
.Y(n_16254)
);

NAND3xp33_ASAP7_75t_L g16255 ( 
.A(n_15209),
.B(n_15223),
.C(n_15196),
.Y(n_16255)
);

NAND2xp5_ASAP7_75t_SL g16256 ( 
.A(n_15344),
.B(n_10821),
.Y(n_16256)
);

NAND3xp33_ASAP7_75t_L g16257 ( 
.A(n_15739),
.B(n_12077),
.C(n_11606),
.Y(n_16257)
);

AOI22xp33_ASAP7_75t_L g16258 ( 
.A1(n_15745),
.A2(n_10942),
.B1(n_10906),
.B2(n_9965),
.Y(n_16258)
);

NAND3xp33_ASAP7_75t_L g16259 ( 
.A(n_15603),
.B(n_12077),
.C(n_11606),
.Y(n_16259)
);

NAND2xp5_ASAP7_75t_L g16260 ( 
.A(n_15216),
.B(n_11078),
.Y(n_16260)
);

NAND2xp5_ASAP7_75t_L g16261 ( 
.A(n_15098),
.B(n_11086),
.Y(n_16261)
);

AOI211xp5_ASAP7_75t_L g16262 ( 
.A1(n_15645),
.A2(n_10834),
.B(n_11002),
.C(n_10821),
.Y(n_16262)
);

NAND2xp5_ASAP7_75t_L g16263 ( 
.A(n_15137),
.B(n_15159),
.Y(n_16263)
);

NAND2xp5_ASAP7_75t_SL g16264 ( 
.A(n_15658),
.B(n_10821),
.Y(n_16264)
);

NAND2xp5_ASAP7_75t_L g16265 ( 
.A(n_15241),
.B(n_11086),
.Y(n_16265)
);

OAI221xp5_ASAP7_75t_L g16266 ( 
.A1(n_15532),
.A2(n_11242),
.B1(n_11287),
.B2(n_11227),
.C(n_11183),
.Y(n_16266)
);

NAND3xp33_ASAP7_75t_L g16267 ( 
.A(n_15651),
.B(n_11606),
.C(n_10497),
.Y(n_16267)
);

NAND2xp5_ASAP7_75t_L g16268 ( 
.A(n_15243),
.B(n_11096),
.Y(n_16268)
);

NAND2xp5_ASAP7_75t_L g16269 ( 
.A(n_15673),
.B(n_11096),
.Y(n_16269)
);

NAND3xp33_ASAP7_75t_L g16270 ( 
.A(n_15659),
.B(n_11606),
.C(n_10497),
.Y(n_16270)
);

NAND2xp5_ASAP7_75t_L g16271 ( 
.A(n_15674),
.B(n_11098),
.Y(n_16271)
);

NAND2xp5_ASAP7_75t_L g16272 ( 
.A(n_15675),
.B(n_11098),
.Y(n_16272)
);

NAND3xp33_ASAP7_75t_L g16273 ( 
.A(n_15562),
.B(n_10497),
.C(n_11822),
.Y(n_16273)
);

AND2x2_ASAP7_75t_L g16274 ( 
.A(n_15376),
.B(n_11103),
.Y(n_16274)
);

NAND2xp5_ASAP7_75t_SL g16275 ( 
.A(n_15658),
.B(n_10821),
.Y(n_16275)
);

OAI22xp33_ASAP7_75t_L g16276 ( 
.A1(n_15831),
.A2(n_10024),
.B1(n_10033),
.B2(n_9967),
.Y(n_16276)
);

NAND2xp5_ASAP7_75t_L g16277 ( 
.A(n_15648),
.B(n_11103),
.Y(n_16277)
);

NAND2xp5_ASAP7_75t_L g16278 ( 
.A(n_15650),
.B(n_11104),
.Y(n_16278)
);

NAND2xp5_ASAP7_75t_L g16279 ( 
.A(n_15665),
.B(n_11104),
.Y(n_16279)
);

NAND2xp5_ASAP7_75t_L g16280 ( 
.A(n_15669),
.B(n_11106),
.Y(n_16280)
);

AND2x2_ASAP7_75t_L g16281 ( 
.A(n_15380),
.B(n_11106),
.Y(n_16281)
);

NAND3xp33_ASAP7_75t_L g16282 ( 
.A(n_15562),
.B(n_10497),
.C(n_11822),
.Y(n_16282)
);

AND2x2_ASAP7_75t_L g16283 ( 
.A(n_15385),
.B(n_11109),
.Y(n_16283)
);

AND2x2_ASAP7_75t_L g16284 ( 
.A(n_15339),
.B(n_11109),
.Y(n_16284)
);

AOI22xp33_ASAP7_75t_L g16285 ( 
.A1(n_15343),
.A2(n_15611),
.B1(n_15676),
.B2(n_15670),
.Y(n_16285)
);

OAI22xp5_ASAP7_75t_L g16286 ( 
.A1(n_15072),
.A2(n_9967),
.B1(n_10033),
.B2(n_10024),
.Y(n_16286)
);

AOI221xp5_ASAP7_75t_L g16287 ( 
.A1(n_15451),
.A2(n_14998),
.B1(n_10033),
.B2(n_10024),
.C(n_9967),
.Y(n_16287)
);

AND2x2_ASAP7_75t_L g16288 ( 
.A(n_15237),
.B(n_11110),
.Y(n_16288)
);

NAND3xp33_ASAP7_75t_L g16289 ( 
.A(n_15794),
.B(n_10497),
.C(n_11822),
.Y(n_16289)
);

NAND2xp5_ASAP7_75t_L g16290 ( 
.A(n_15253),
.B(n_11110),
.Y(n_16290)
);

AND2x2_ASAP7_75t_L g16291 ( 
.A(n_15238),
.B(n_11111),
.Y(n_16291)
);

NAND4xp25_ASAP7_75t_L g16292 ( 
.A(n_15035),
.B(n_9561),
.C(n_9582),
.D(n_9573),
.Y(n_16292)
);

AND2x2_ASAP7_75t_L g16293 ( 
.A(n_15240),
.B(n_11111),
.Y(n_16293)
);

NAND2xp5_ASAP7_75t_L g16294 ( 
.A(n_15271),
.B(n_11117),
.Y(n_16294)
);

NAND2xp5_ASAP7_75t_L g16295 ( 
.A(n_15282),
.B(n_11117),
.Y(n_16295)
);

NAND3xp33_ASAP7_75t_L g16296 ( 
.A(n_15834),
.B(n_10497),
.C(n_13445),
.Y(n_16296)
);

NAND3xp33_ASAP7_75t_L g16297 ( 
.A(n_15666),
.B(n_13468),
.C(n_10865),
.Y(n_16297)
);

NOR2xp33_ASAP7_75t_L g16298 ( 
.A(n_15431),
.B(n_10135),
.Y(n_16298)
);

AND2x2_ASAP7_75t_L g16299 ( 
.A(n_15245),
.B(n_11132),
.Y(n_16299)
);

NAND2xp5_ASAP7_75t_L g16300 ( 
.A(n_15285),
.B(n_11132),
.Y(n_16300)
);

NAND2xp5_ASAP7_75t_L g16301 ( 
.A(n_15293),
.B(n_11142),
.Y(n_16301)
);

AOI22xp33_ASAP7_75t_SL g16302 ( 
.A1(n_15310),
.A2(n_10024),
.B1(n_10033),
.B2(n_9967),
.Y(n_16302)
);

AOI221xp5_ASAP7_75t_L g16303 ( 
.A1(n_15520),
.A2(n_10033),
.B1(n_10024),
.B2(n_9967),
.C(n_10821),
.Y(n_16303)
);

NAND2xp5_ASAP7_75t_L g16304 ( 
.A(n_15296),
.B(n_11142),
.Y(n_16304)
);

AOI22xp33_ASAP7_75t_SL g16305 ( 
.A1(n_15390),
.A2(n_10024),
.B1(n_10033),
.B2(n_9967),
.Y(n_16305)
);

NAND2xp5_ASAP7_75t_L g16306 ( 
.A(n_15303),
.B(n_9364),
.Y(n_16306)
);

INVx2_ASAP7_75t_L g16307 ( 
.A(n_15046),
.Y(n_16307)
);

NAND3xp33_ASAP7_75t_L g16308 ( 
.A(n_15511),
.B(n_13468),
.C(n_10865),
.Y(n_16308)
);

NAND2xp5_ASAP7_75t_L g16309 ( 
.A(n_15308),
.B(n_15311),
.Y(n_16309)
);

NAND2xp5_ASAP7_75t_SL g16310 ( 
.A(n_15681),
.B(n_10834),
.Y(n_16310)
);

NAND2xp5_ASAP7_75t_L g16311 ( 
.A(n_15104),
.B(n_9364),
.Y(n_16311)
);

NAND2xp5_ASAP7_75t_L g16312 ( 
.A(n_15361),
.B(n_9364),
.Y(n_16312)
);

NOR2xp33_ASAP7_75t_L g16313 ( 
.A(n_15433),
.B(n_9019),
.Y(n_16313)
);

NAND2xp5_ASAP7_75t_L g16314 ( 
.A(n_15435),
.B(n_9364),
.Y(n_16314)
);

OAI22xp5_ASAP7_75t_L g16315 ( 
.A1(n_15471),
.A2(n_9967),
.B1(n_10033),
.B2(n_10024),
.Y(n_16315)
);

AND2x2_ASAP7_75t_L g16316 ( 
.A(n_15625),
.B(n_14565),
.Y(n_16316)
);

NAND2xp5_ASAP7_75t_L g16317 ( 
.A(n_15272),
.B(n_9364),
.Y(n_16317)
);

NAND2xp5_ASAP7_75t_L g16318 ( 
.A(n_15236),
.B(n_9376),
.Y(n_16318)
);

OAI221xp5_ASAP7_75t_SL g16319 ( 
.A1(n_15534),
.A2(n_10814),
.B1(n_10858),
.B2(n_10758),
.C(n_10593),
.Y(n_16319)
);

AND2x2_ASAP7_75t_L g16320 ( 
.A(n_15632),
.B(n_14565),
.Y(n_16320)
);

NAND3xp33_ASAP7_75t_L g16321 ( 
.A(n_15225),
.B(n_10865),
.C(n_10857),
.Y(n_16321)
);

NAND2xp5_ASAP7_75t_L g16322 ( 
.A(n_15225),
.B(n_9376),
.Y(n_16322)
);

AND2x2_ASAP7_75t_L g16323 ( 
.A(n_15799),
.B(n_11470),
.Y(n_16323)
);

INVx1_ASAP7_75t_L g16324 ( 
.A(n_15309),
.Y(n_16324)
);

AND2x2_ASAP7_75t_L g16325 ( 
.A(n_15545),
.B(n_11470),
.Y(n_16325)
);

NAND2xp5_ASAP7_75t_L g16326 ( 
.A(n_15289),
.B(n_9376),
.Y(n_16326)
);

NAND2xp5_ASAP7_75t_L g16327 ( 
.A(n_15289),
.B(n_9376),
.Y(n_16327)
);

AND2x2_ASAP7_75t_L g16328 ( 
.A(n_15547),
.B(n_11470),
.Y(n_16328)
);

OAI221xp5_ASAP7_75t_L g16329 ( 
.A1(n_15535),
.A2(n_11183),
.B1(n_11287),
.B2(n_11242),
.C(n_11227),
.Y(n_16329)
);

AND2x2_ASAP7_75t_L g16330 ( 
.A(n_15555),
.B(n_11489),
.Y(n_16330)
);

NAND2xp5_ASAP7_75t_SL g16331 ( 
.A(n_15681),
.B(n_10834),
.Y(n_16331)
);

NAND2xp5_ASAP7_75t_L g16332 ( 
.A(n_15298),
.B(n_9376),
.Y(n_16332)
);

NAND2xp5_ASAP7_75t_L g16333 ( 
.A(n_15298),
.B(n_9320),
.Y(n_16333)
);

OAI221xp5_ASAP7_75t_L g16334 ( 
.A1(n_15629),
.A2(n_11312),
.B1(n_11327),
.B2(n_11287),
.C(n_11242),
.Y(n_16334)
);

NAND3xp33_ASAP7_75t_L g16335 ( 
.A(n_15828),
.B(n_10865),
.C(n_10857),
.Y(n_16335)
);

OAI22xp5_ASAP7_75t_L g16336 ( 
.A1(n_15471),
.A2(n_9967),
.B1(n_10033),
.B2(n_10024),
.Y(n_16336)
);

OAI221xp5_ASAP7_75t_SL g16337 ( 
.A1(n_15837),
.A2(n_10858),
.B1(n_10814),
.B2(n_9117),
.C(n_11340),
.Y(n_16337)
);

AOI221xp5_ASAP7_75t_L g16338 ( 
.A1(n_15787),
.A2(n_10033),
.B1(n_10024),
.B2(n_9967),
.C(n_10834),
.Y(n_16338)
);

NAND3xp33_ASAP7_75t_L g16339 ( 
.A(n_15841),
.B(n_10865),
.C(n_10857),
.Y(n_16339)
);

OAI21xp5_ASAP7_75t_SL g16340 ( 
.A1(n_15741),
.A2(n_11287),
.B(n_11242),
.Y(n_16340)
);

OAI22xp5_ASAP7_75t_L g16341 ( 
.A1(n_15634),
.A2(n_10024),
.B1(n_10033),
.B2(n_9117),
.Y(n_16341)
);

OAI221xp5_ASAP7_75t_L g16342 ( 
.A1(n_15400),
.A2(n_11352),
.B1(n_11361),
.B2(n_11327),
.C(n_11312),
.Y(n_16342)
);

NAND2xp5_ASAP7_75t_L g16343 ( 
.A(n_15325),
.B(n_9320),
.Y(n_16343)
);

AND2x2_ASAP7_75t_L g16344 ( 
.A(n_15561),
.B(n_11489),
.Y(n_16344)
);

OAI221xp5_ASAP7_75t_L g16345 ( 
.A1(n_15721),
.A2(n_11352),
.B1(n_11361),
.B2(n_11327),
.C(n_11312),
.Y(n_16345)
);

NAND3xp33_ASAP7_75t_L g16346 ( 
.A(n_15263),
.B(n_10865),
.C(n_10857),
.Y(n_16346)
);

NAND2xp5_ASAP7_75t_L g16347 ( 
.A(n_15325),
.B(n_9320),
.Y(n_16347)
);

NAND3xp33_ASAP7_75t_L g16348 ( 
.A(n_15049),
.B(n_10857),
.C(n_11927),
.Y(n_16348)
);

AND2x2_ASAP7_75t_L g16349 ( 
.A(n_15575),
.B(n_11489),
.Y(n_16349)
);

NAND2xp5_ASAP7_75t_L g16350 ( 
.A(n_15331),
.B(n_9320),
.Y(n_16350)
);

NAND2xp5_ASAP7_75t_L g16351 ( 
.A(n_15331),
.B(n_9320),
.Y(n_16351)
);

NOR2x1_ASAP7_75t_SL g16352 ( 
.A(n_15228),
.B(n_10834),
.Y(n_16352)
);

AND2x2_ASAP7_75t_SL g16353 ( 
.A(n_15173),
.B(n_9792),
.Y(n_16353)
);

NAND2xp5_ASAP7_75t_SL g16354 ( 
.A(n_15694),
.B(n_10834),
.Y(n_16354)
);

NAND2xp5_ASAP7_75t_L g16355 ( 
.A(n_15769),
.B(n_11461),
.Y(n_16355)
);

NAND2xp5_ASAP7_75t_L g16356 ( 
.A(n_15176),
.B(n_11461),
.Y(n_16356)
);

NAND2xp5_ASAP7_75t_L g16357 ( 
.A(n_15318),
.B(n_15393),
.Y(n_16357)
);

NAND2xp5_ASAP7_75t_L g16358 ( 
.A(n_15403),
.B(n_11461),
.Y(n_16358)
);

OAI22xp33_ASAP7_75t_SL g16359 ( 
.A1(n_15642),
.A2(n_11327),
.B1(n_11352),
.B2(n_11312),
.Y(n_16359)
);

NAND2xp5_ASAP7_75t_L g16360 ( 
.A(n_15422),
.B(n_9209),
.Y(n_16360)
);

OAI221xp5_ASAP7_75t_L g16361 ( 
.A1(n_15470),
.A2(n_11362),
.B1(n_11575),
.B2(n_11361),
.C(n_11352),
.Y(n_16361)
);

OAI22xp5_ASAP7_75t_L g16362 ( 
.A1(n_15744),
.A2(n_10024),
.B1(n_10033),
.B2(n_9117),
.Y(n_16362)
);

AOI22xp33_ASAP7_75t_L g16363 ( 
.A1(n_15678),
.A2(n_10942),
.B1(n_10906),
.B2(n_9965),
.Y(n_16363)
);

NAND2xp5_ASAP7_75t_L g16364 ( 
.A(n_15305),
.B(n_9209),
.Y(n_16364)
);

NAND3xp33_ASAP7_75t_L g16365 ( 
.A(n_15049),
.B(n_10857),
.C(n_11927),
.Y(n_16365)
);

AND2x2_ASAP7_75t_L g16366 ( 
.A(n_15576),
.B(n_11490),
.Y(n_16366)
);

NAND2xp5_ASAP7_75t_L g16367 ( 
.A(n_15307),
.B(n_9209),
.Y(n_16367)
);

AND2x2_ASAP7_75t_L g16368 ( 
.A(n_15577),
.B(n_15582),
.Y(n_16368)
);

NAND3xp33_ASAP7_75t_L g16369 ( 
.A(n_15056),
.B(n_11948),
.C(n_11927),
.Y(n_16369)
);

NAND2xp5_ASAP7_75t_L g16370 ( 
.A(n_15314),
.B(n_9209),
.Y(n_16370)
);

AND2x2_ASAP7_75t_L g16371 ( 
.A(n_15312),
.B(n_11490),
.Y(n_16371)
);

NAND2xp5_ASAP7_75t_L g16372 ( 
.A(n_15315),
.B(n_9209),
.Y(n_16372)
);

HB1xp67_ASAP7_75t_L g16373 ( 
.A(n_15056),
.Y(n_16373)
);

NAND2xp5_ASAP7_75t_L g16374 ( 
.A(n_15426),
.B(n_9224),
.Y(n_16374)
);

NAND2xp5_ASAP7_75t_SL g16375 ( 
.A(n_15694),
.B(n_10834),
.Y(n_16375)
);

NAND2xp5_ASAP7_75t_L g16376 ( 
.A(n_15362),
.B(n_9224),
.Y(n_16376)
);

NAND2xp5_ASAP7_75t_L g16377 ( 
.A(n_15295),
.B(n_9224),
.Y(n_16377)
);

NAND2xp5_ASAP7_75t_L g16378 ( 
.A(n_15713),
.B(n_9224),
.Y(n_16378)
);

NAND2xp5_ASAP7_75t_L g16379 ( 
.A(n_15714),
.B(n_9224),
.Y(n_16379)
);

NAND2xp5_ASAP7_75t_L g16380 ( 
.A(n_15277),
.B(n_15292),
.Y(n_16380)
);

NAND2xp5_ASAP7_75t_L g16381 ( 
.A(n_15723),
.B(n_9264),
.Y(n_16381)
);

AOI211xp5_ASAP7_75t_L g16382 ( 
.A1(n_15760),
.A2(n_11002),
.B(n_11224),
.C(n_10834),
.Y(n_16382)
);

INVx1_ASAP7_75t_L g16383 ( 
.A(n_15320),
.Y(n_16383)
);

OA21x2_ASAP7_75t_L g16384 ( 
.A1(n_15320),
.A2(n_10895),
.B(n_10889),
.Y(n_16384)
);

OAI21xp5_ASAP7_75t_L g16385 ( 
.A1(n_15323),
.A2(n_10873),
.B(n_10872),
.Y(n_16385)
);

OAI21xp33_ASAP7_75t_L g16386 ( 
.A1(n_15478),
.A2(n_9573),
.B(n_9561),
.Y(n_16386)
);

OAI22xp5_ASAP7_75t_L g16387 ( 
.A1(n_15744),
.A2(n_10033),
.B1(n_9117),
.B2(n_10036),
.Y(n_16387)
);

AND2x2_ASAP7_75t_L g16388 ( 
.A(n_15360),
.B(n_11490),
.Y(n_16388)
);

NAND3xp33_ASAP7_75t_L g16389 ( 
.A(n_15221),
.B(n_11948),
.C(n_10569),
.Y(n_16389)
);

NAND2xp5_ASAP7_75t_L g16390 ( 
.A(n_15737),
.B(n_9264),
.Y(n_16390)
);

NAND2xp5_ASAP7_75t_L g16391 ( 
.A(n_15757),
.B(n_9264),
.Y(n_16391)
);

OR2x2_ASAP7_75t_L g16392 ( 
.A(n_15290),
.B(n_11452),
.Y(n_16392)
);

AND2x2_ASAP7_75t_L g16393 ( 
.A(n_15370),
.B(n_10642),
.Y(n_16393)
);

NAND2xp5_ASAP7_75t_L g16394 ( 
.A(n_15759),
.B(n_9264),
.Y(n_16394)
);

OAI221xp5_ASAP7_75t_L g16395 ( 
.A1(n_15485),
.A2(n_11575),
.B1(n_11610),
.B2(n_11362),
.C(n_11361),
.Y(n_16395)
);

AND2x2_ASAP7_75t_L g16396 ( 
.A(n_15394),
.B(n_10642),
.Y(n_16396)
);

NAND3xp33_ASAP7_75t_L g16397 ( 
.A(n_15221),
.B(n_11948),
.C(n_10569),
.Y(n_16397)
);

NAND2xp5_ASAP7_75t_L g16398 ( 
.A(n_15328),
.B(n_9264),
.Y(n_16398)
);

AND2x2_ASAP7_75t_L g16399 ( 
.A(n_15407),
.B(n_10642),
.Y(n_16399)
);

AOI221xp5_ASAP7_75t_L g16400 ( 
.A1(n_15825),
.A2(n_10033),
.B1(n_11224),
.B2(n_11276),
.C(n_11002),
.Y(n_16400)
);

NAND2xp5_ASAP7_75t_L g16401 ( 
.A(n_15336),
.B(n_9343),
.Y(n_16401)
);

NAND2xp5_ASAP7_75t_L g16402 ( 
.A(n_15337),
.B(n_15446),
.Y(n_16402)
);

AND2x2_ASAP7_75t_L g16403 ( 
.A(n_15409),
.B(n_15410),
.Y(n_16403)
);

NOR3xp33_ASAP7_75t_L g16404 ( 
.A(n_15097),
.B(n_10314),
.C(n_10591),
.Y(n_16404)
);

OA211x2_ASAP7_75t_L g16405 ( 
.A1(n_15621),
.A2(n_9335),
.B(n_9249),
.C(n_9870),
.Y(n_16405)
);

NAND3xp33_ASAP7_75t_L g16406 ( 
.A(n_15827),
.B(n_15624),
.C(n_15074),
.Y(n_16406)
);

AND2x2_ASAP7_75t_L g16407 ( 
.A(n_15428),
.B(n_15719),
.Y(n_16407)
);

AND2x2_ASAP7_75t_L g16408 ( 
.A(n_15452),
.B(n_9343),
.Y(n_16408)
);

AOI221xp5_ASAP7_75t_L g16409 ( 
.A1(n_15421),
.A2(n_11002),
.B1(n_11469),
.B2(n_11276),
.C(n_11224),
.Y(n_16409)
);

OA21x2_ASAP7_75t_L g16410 ( 
.A1(n_15341),
.A2(n_10903),
.B(n_10895),
.Y(n_16410)
);

NAND3xp33_ASAP7_75t_L g16411 ( 
.A(n_15070),
.B(n_10569),
.C(n_9741),
.Y(n_16411)
);

OA21x2_ASAP7_75t_L g16412 ( 
.A1(n_15341),
.A2(n_10905),
.B(n_10903),
.Y(n_16412)
);

NAND2xp5_ASAP7_75t_L g16413 ( 
.A(n_15350),
.B(n_9343),
.Y(n_16413)
);

NAND3xp33_ASAP7_75t_L g16414 ( 
.A(n_15076),
.B(n_15081),
.C(n_15077),
.Y(n_16414)
);

AOI221xp5_ASAP7_75t_L g16415 ( 
.A1(n_15086),
.A2(n_11002),
.B1(n_11469),
.B2(n_11276),
.C(n_11224),
.Y(n_16415)
);

NAND2xp5_ASAP7_75t_L g16416 ( 
.A(n_15351),
.B(n_9343),
.Y(n_16416)
);

AND2x2_ASAP7_75t_SL g16417 ( 
.A(n_15425),
.B(n_9792),
.Y(n_16417)
);

AOI22xp33_ASAP7_75t_SL g16418 ( 
.A1(n_15716),
.A2(n_10159),
.B1(n_10137),
.B2(n_10048),
.Y(n_16418)
);

AND2x2_ASAP7_75t_L g16419 ( 
.A(n_15552),
.B(n_15556),
.Y(n_16419)
);

AND2x2_ASAP7_75t_L g16420 ( 
.A(n_15570),
.B(n_9343),
.Y(n_16420)
);

NAND2xp5_ASAP7_75t_L g16421 ( 
.A(n_15356),
.B(n_9112),
.Y(n_16421)
);

NAND3xp33_ASAP7_75t_L g16422 ( 
.A(n_15090),
.B(n_10569),
.C(n_9741),
.Y(n_16422)
);

AOI221xp5_ASAP7_75t_L g16423 ( 
.A1(n_15100),
.A2(n_11002),
.B1(n_11469),
.B2(n_11276),
.C(n_11224),
.Y(n_16423)
);

OA211x2_ASAP7_75t_L g16424 ( 
.A1(n_15094),
.A2(n_9335),
.B(n_9249),
.C(n_9870),
.Y(n_16424)
);

OAI21xp5_ASAP7_75t_L g16425 ( 
.A1(n_15710),
.A2(n_15573),
.B(n_15818),
.Y(n_16425)
);

NAND2xp5_ASAP7_75t_SL g16426 ( 
.A(n_15516),
.B(n_11002),
.Y(n_16426)
);

NAND3xp33_ASAP7_75t_L g16427 ( 
.A(n_15103),
.B(n_10569),
.C(n_9741),
.Y(n_16427)
);

AND2x2_ASAP7_75t_L g16428 ( 
.A(n_15605),
.B(n_10083),
.Y(n_16428)
);

OAI21xp5_ASAP7_75t_L g16429 ( 
.A1(n_15553),
.A2(n_10761),
.B(n_10767),
.Y(n_16429)
);

AND2x2_ASAP7_75t_L g16430 ( 
.A(n_15613),
.B(n_10083),
.Y(n_16430)
);

OAI21xp5_ASAP7_75t_SL g16431 ( 
.A1(n_15751),
.A2(n_15440),
.B(n_15438),
.Y(n_16431)
);

NAND3xp33_ASAP7_75t_L g16432 ( 
.A(n_15119),
.B(n_10569),
.C(n_9741),
.Y(n_16432)
);

NOR3xp33_ASAP7_75t_SL g16433 ( 
.A(n_15107),
.B(n_8737),
.C(n_9502),
.Y(n_16433)
);

NAND2xp33_ASAP7_75t_L g16434 ( 
.A(n_15146),
.B(n_11002),
.Y(n_16434)
);

AND2x2_ASAP7_75t_L g16435 ( 
.A(n_15620),
.B(n_15685),
.Y(n_16435)
);

NAND2xp5_ASAP7_75t_L g16436 ( 
.A(n_15441),
.B(n_9112),
.Y(n_16436)
);

AND2x2_ASAP7_75t_L g16437 ( 
.A(n_15700),
.B(n_10083),
.Y(n_16437)
);

OAI21xp33_ASAP7_75t_L g16438 ( 
.A1(n_15609),
.A2(n_9573),
.B(n_9561),
.Y(n_16438)
);

OAI221xp5_ASAP7_75t_SL g16439 ( 
.A1(n_15829),
.A2(n_15427),
.B1(n_15692),
.B2(n_15275),
.C(n_15009),
.Y(n_16439)
);

AND2x2_ASAP7_75t_L g16440 ( 
.A(n_15707),
.B(n_10083),
.Y(n_16440)
);

OAI22xp5_ASAP7_75t_L g16441 ( 
.A1(n_15016),
.A2(n_9117),
.B1(n_10048),
.B2(n_10036),
.Y(n_16441)
);

AND2x2_ASAP7_75t_L g16442 ( 
.A(n_15708),
.B(n_15711),
.Y(n_16442)
);

AND2x2_ASAP7_75t_L g16443 ( 
.A(n_15715),
.B(n_10083),
.Y(n_16443)
);

OAI221xp5_ASAP7_75t_SL g16444 ( 
.A1(n_15427),
.A2(n_10858),
.B1(n_11380),
.B2(n_11340),
.C(n_11408),
.Y(n_16444)
);

NAND2xp5_ASAP7_75t_L g16445 ( 
.A(n_15550),
.B(n_9112),
.Y(n_16445)
);

NAND2xp5_ASAP7_75t_L g16446 ( 
.A(n_15255),
.B(n_9112),
.Y(n_16446)
);

AND2x2_ASAP7_75t_L g16447 ( 
.A(n_15638),
.B(n_10187),
.Y(n_16447)
);

NAND2xp5_ASAP7_75t_L g16448 ( 
.A(n_15347),
.B(n_9112),
.Y(n_16448)
);

AND2x2_ASAP7_75t_L g16449 ( 
.A(n_15724),
.B(n_15727),
.Y(n_16449)
);

OAI221xp5_ASAP7_75t_SL g16450 ( 
.A1(n_15316),
.A2(n_11380),
.B1(n_11544),
.B2(n_11408),
.C(n_11578),
.Y(n_16450)
);

AND2x2_ASAP7_75t_L g16451 ( 
.A(n_15735),
.B(n_10187),
.Y(n_16451)
);

NAND2xp5_ASAP7_75t_L g16452 ( 
.A(n_15749),
.B(n_9121),
.Y(n_16452)
);

INVx1_ASAP7_75t_L g16453 ( 
.A(n_15353),
.Y(n_16453)
);

OAI21xp5_ASAP7_75t_SL g16454 ( 
.A1(n_15349),
.A2(n_11575),
.B(n_11362),
.Y(n_16454)
);

AOI221xp5_ASAP7_75t_L g16455 ( 
.A1(n_15126),
.A2(n_11224),
.B1(n_11478),
.B2(n_11469),
.C(n_11276),
.Y(n_16455)
);

AND2x2_ASAP7_75t_L g16456 ( 
.A(n_15750),
.B(n_10187),
.Y(n_16456)
);

AND2x2_ASAP7_75t_L g16457 ( 
.A(n_15754),
.B(n_10187),
.Y(n_16457)
);

AND2x2_ASAP7_75t_L g16458 ( 
.A(n_15765),
.B(n_10187),
.Y(n_16458)
);

OAI22xp5_ASAP7_75t_L g16459 ( 
.A1(n_15024),
.A2(n_10048),
.B1(n_10110),
.B2(n_10036),
.Y(n_16459)
);

OAI22xp5_ASAP7_75t_L g16460 ( 
.A1(n_15456),
.A2(n_10048),
.B1(n_10110),
.B2(n_10036),
.Y(n_16460)
);

NAND2xp5_ASAP7_75t_L g16461 ( 
.A(n_15768),
.B(n_9121),
.Y(n_16461)
);

AND2x2_ASAP7_75t_L g16462 ( 
.A(n_15772),
.B(n_9019),
.Y(n_16462)
);

NAND2xp5_ASAP7_75t_L g16463 ( 
.A(n_15788),
.B(n_9121),
.Y(n_16463)
);

NAND3xp33_ASAP7_75t_L g16464 ( 
.A(n_15127),
.B(n_9741),
.C(n_9723),
.Y(n_16464)
);

AND2x2_ASAP7_75t_L g16465 ( 
.A(n_15803),
.B(n_9019),
.Y(n_16465)
);

NAND2xp5_ASAP7_75t_L g16466 ( 
.A(n_15809),
.B(n_9121),
.Y(n_16466)
);

AND2x2_ASAP7_75t_L g16467 ( 
.A(n_15815),
.B(n_9019),
.Y(n_16467)
);

AND2x2_ASAP7_75t_L g16468 ( 
.A(n_15822),
.B(n_9019),
.Y(n_16468)
);

NAND3xp33_ASAP7_75t_L g16469 ( 
.A(n_15133),
.B(n_9741),
.C(n_9723),
.Y(n_16469)
);

AND2x2_ASAP7_75t_L g16470 ( 
.A(n_15720),
.B(n_9019),
.Y(n_16470)
);

INVx1_ASAP7_75t_L g16471 ( 
.A(n_15353),
.Y(n_16471)
);

OAI21xp5_ASAP7_75t_L g16472 ( 
.A1(n_15538),
.A2(n_10761),
.B(n_10767),
.Y(n_16472)
);

AND2x2_ASAP7_75t_L g16473 ( 
.A(n_15533),
.B(n_15563),
.Y(n_16473)
);

NAND2xp5_ASAP7_75t_L g16474 ( 
.A(n_15136),
.B(n_9121),
.Y(n_16474)
);

OAI221xp5_ASAP7_75t_L g16475 ( 
.A1(n_15622),
.A2(n_11362),
.B1(n_11616),
.B2(n_11610),
.C(n_11575),
.Y(n_16475)
);

NAND3xp33_ASAP7_75t_L g16476 ( 
.A(n_15139),
.B(n_9741),
.C(n_9723),
.Y(n_16476)
);

OAI221xp5_ASAP7_75t_L g16477 ( 
.A1(n_15672),
.A2(n_11616),
.B1(n_11610),
.B2(n_11469),
.C(n_11478),
.Y(n_16477)
);

OAI21xp33_ASAP7_75t_SL g16478 ( 
.A1(n_15539),
.A2(n_12905),
.B(n_11614),
.Y(n_16478)
);

AND2x2_ASAP7_75t_L g16479 ( 
.A(n_15748),
.B(n_9019),
.Y(n_16479)
);

AND2x2_ASAP7_75t_L g16480 ( 
.A(n_15449),
.B(n_9019),
.Y(n_16480)
);

AND2x2_ASAP7_75t_L g16481 ( 
.A(n_15461),
.B(n_15467),
.Y(n_16481)
);

AND2x2_ASAP7_75t_L g16482 ( 
.A(n_15510),
.B(n_9040),
.Y(n_16482)
);

AND2x2_ASAP7_75t_L g16483 ( 
.A(n_15568),
.B(n_9040),
.Y(n_16483)
);

AND2x2_ASAP7_75t_L g16484 ( 
.A(n_15736),
.B(n_9040),
.Y(n_16484)
);

NAND2xp5_ASAP7_75t_L g16485 ( 
.A(n_15145),
.B(n_9126),
.Y(n_16485)
);

NAND2xp5_ASAP7_75t_L g16486 ( 
.A(n_15149),
.B(n_9126),
.Y(n_16486)
);

NAND2xp5_ASAP7_75t_L g16487 ( 
.A(n_15154),
.B(n_9126),
.Y(n_16487)
);

AOI22xp5_ASAP7_75t_L g16488 ( 
.A1(n_15476),
.A2(n_15770),
.B1(n_15524),
.B2(n_15702),
.Y(n_16488)
);

NAND2xp33_ASAP7_75t_SL g16489 ( 
.A(n_15229),
.B(n_11224),
.Y(n_16489)
);

NAND2xp5_ASAP7_75t_L g16490 ( 
.A(n_15166),
.B(n_9126),
.Y(n_16490)
);

NAND3xp33_ASAP7_75t_L g16491 ( 
.A(n_15178),
.B(n_9741),
.C(n_9723),
.Y(n_16491)
);

AOI22xp5_ASAP7_75t_L g16492 ( 
.A1(n_15476),
.A2(n_10159),
.B1(n_10137),
.B2(n_9775),
.Y(n_16492)
);

OAI21xp33_ASAP7_75t_L g16493 ( 
.A1(n_15262),
.A2(n_9573),
.B(n_9561),
.Y(n_16493)
);

AND2x2_ASAP7_75t_L g16494 ( 
.A(n_15690),
.B(n_9040),
.Y(n_16494)
);

AND2x2_ASAP7_75t_L g16495 ( 
.A(n_15169),
.B(n_9040),
.Y(n_16495)
);

NAND2xp5_ASAP7_75t_L g16496 ( 
.A(n_15186),
.B(n_9126),
.Y(n_16496)
);

AOI22xp33_ASAP7_75t_L g16497 ( 
.A1(n_15777),
.A2(n_10942),
.B1(n_10906),
.B2(n_9965),
.Y(n_16497)
);

NAND2xp5_ASAP7_75t_L g16498 ( 
.A(n_15192),
.B(n_9153),
.Y(n_16498)
);

NAND2xp5_ASAP7_75t_SL g16499 ( 
.A(n_15516),
.B(n_11224),
.Y(n_16499)
);

NAND4xp25_ASAP7_75t_L g16500 ( 
.A(n_15763),
.B(n_9561),
.C(n_9582),
.D(n_9573),
.Y(n_16500)
);

NOR2xp67_ASAP7_75t_L g16501 ( 
.A(n_15386),
.B(n_15174),
.Y(n_16501)
);

NAND2xp5_ASAP7_75t_L g16502 ( 
.A(n_15201),
.B(n_9153),
.Y(n_16502)
);

AND2x2_ASAP7_75t_L g16503 ( 
.A(n_15789),
.B(n_9040),
.Y(n_16503)
);

AND2x2_ASAP7_75t_L g16504 ( 
.A(n_15664),
.B(n_9040),
.Y(n_16504)
);

AND2x2_ASAP7_75t_L g16505 ( 
.A(n_15664),
.B(n_9040),
.Y(n_16505)
);

NAND2xp5_ASAP7_75t_L g16506 ( 
.A(n_15203),
.B(n_9153),
.Y(n_16506)
);

OAI221xp5_ASAP7_75t_SL g16507 ( 
.A1(n_15322),
.A2(n_11380),
.B1(n_11544),
.B2(n_11408),
.C(n_11578),
.Y(n_16507)
);

AOI22xp33_ASAP7_75t_L g16508 ( 
.A1(n_15847),
.A2(n_10942),
.B1(n_10906),
.B2(n_9965),
.Y(n_16508)
);

AOI21xp5_ASAP7_75t_L g16509 ( 
.A1(n_15548),
.A2(n_14829),
.B(n_14828),
.Y(n_16509)
);

NAND2xp5_ASAP7_75t_L g16510 ( 
.A(n_15208),
.B(n_9153),
.Y(n_16510)
);

NAND3xp33_ASAP7_75t_L g16511 ( 
.A(n_15211),
.B(n_9741),
.C(n_9723),
.Y(n_16511)
);

OAI221xp5_ASAP7_75t_L g16512 ( 
.A1(n_15278),
.A2(n_15424),
.B1(n_15195),
.B2(n_15368),
.C(n_15355),
.Y(n_16512)
);

AND2x2_ASAP7_75t_L g16513 ( 
.A(n_15756),
.B(n_9054),
.Y(n_16513)
);

NAND2xp5_ASAP7_75t_L g16514 ( 
.A(n_15217),
.B(n_9153),
.Y(n_16514)
);

OAI22xp5_ASAP7_75t_L g16515 ( 
.A1(n_15080),
.A2(n_10048),
.B1(n_10110),
.B2(n_10036),
.Y(n_16515)
);

NAND2xp5_ASAP7_75t_L g16516 ( 
.A(n_15234),
.B(n_9163),
.Y(n_16516)
);

NOR3xp33_ASAP7_75t_L g16517 ( 
.A(n_15108),
.B(n_10591),
.C(n_10023),
.Y(n_16517)
);

AND2x2_ASAP7_75t_L g16518 ( 
.A(n_15758),
.B(n_9054),
.Y(n_16518)
);

NAND2xp5_ASAP7_75t_L g16519 ( 
.A(n_15242),
.B(n_9163),
.Y(n_16519)
);

OAI21xp33_ASAP7_75t_L g16520 ( 
.A1(n_15832),
.A2(n_9582),
.B(n_9561),
.Y(n_16520)
);

AOI21xp5_ASAP7_75t_SL g16521 ( 
.A1(n_15566),
.A2(n_14828),
.B(n_14784),
.Y(n_16521)
);

NOR2xp33_ASAP7_75t_L g16522 ( 
.A(n_15419),
.B(n_9054),
.Y(n_16522)
);

NAND2xp5_ASAP7_75t_L g16523 ( 
.A(n_15248),
.B(n_9163),
.Y(n_16523)
);

NAND2xp33_ASAP7_75t_SL g16524 ( 
.A(n_15747),
.B(n_11276),
.Y(n_16524)
);

AND2x2_ASAP7_75t_L g16525 ( 
.A(n_15551),
.B(n_9054),
.Y(n_16525)
);

NAND2xp5_ASAP7_75t_L g16526 ( 
.A(n_15183),
.B(n_9163),
.Y(n_16526)
);

NAND2xp5_ASAP7_75t_L g16527 ( 
.A(n_15187),
.B(n_9163),
.Y(n_16527)
);

OAI221xp5_ASAP7_75t_SL g16528 ( 
.A1(n_15587),
.A2(n_11544),
.B1(n_11614),
.B2(n_11578),
.C(n_9294),
.Y(n_16528)
);

NAND2xp5_ASAP7_75t_L g16529 ( 
.A(n_15191),
.B(n_9164),
.Y(n_16529)
);

AND2x2_ASAP7_75t_L g16530 ( 
.A(n_15747),
.B(n_9054),
.Y(n_16530)
);

OR2x2_ASAP7_75t_L g16531 ( 
.A(n_15128),
.B(n_11452),
.Y(n_16531)
);

NAND2xp5_ASAP7_75t_L g16532 ( 
.A(n_15232),
.B(n_9164),
.Y(n_16532)
);

NOR3xp33_ASAP7_75t_L g16533 ( 
.A(n_15235),
.B(n_10591),
.C(n_10023),
.Y(n_16533)
);

NAND4xp25_ASAP7_75t_L g16534 ( 
.A(n_15513),
.B(n_9582),
.C(n_8935),
.D(n_9918),
.Y(n_16534)
);

NAND2xp5_ASAP7_75t_L g16535 ( 
.A(n_15135),
.B(n_9164),
.Y(n_16535)
);

OA211x2_ASAP7_75t_L g16536 ( 
.A1(n_15143),
.A2(n_9092),
.B(n_9174),
.C(n_8762),
.Y(n_16536)
);

OAI21xp5_ASAP7_75t_L g16537 ( 
.A1(n_15549),
.A2(n_10761),
.B(n_10767),
.Y(n_16537)
);

AND2x2_ASAP7_75t_L g16538 ( 
.A(n_15566),
.B(n_9054),
.Y(n_16538)
);

NAND3xp33_ASAP7_75t_L g16539 ( 
.A(n_15144),
.B(n_9723),
.C(n_10616),
.Y(n_16539)
);

NAND2xp5_ASAP7_75t_L g16540 ( 
.A(n_15147),
.B(n_9164),
.Y(n_16540)
);

NAND2xp5_ASAP7_75t_SL g16541 ( 
.A(n_15623),
.B(n_11276),
.Y(n_16541)
);

NAND2xp5_ASAP7_75t_L g16542 ( 
.A(n_15157),
.B(n_9164),
.Y(n_16542)
);

AND2x2_ASAP7_75t_L g16543 ( 
.A(n_15623),
.B(n_15766),
.Y(n_16543)
);

AND2x2_ASAP7_75t_L g16544 ( 
.A(n_15702),
.B(n_9054),
.Y(n_16544)
);

NAND3xp33_ASAP7_75t_L g16545 ( 
.A(n_15530),
.B(n_9723),
.C(n_10616),
.Y(n_16545)
);

NAND2xp5_ASAP7_75t_L g16546 ( 
.A(n_15112),
.B(n_11082),
.Y(n_16546)
);

AND2x2_ASAP7_75t_L g16547 ( 
.A(n_15525),
.B(n_9054),
.Y(n_16547)
);

NAND3xp33_ASAP7_75t_L g16548 ( 
.A(n_15276),
.B(n_9723),
.C(n_10616),
.Y(n_16548)
);

HB1xp67_ASAP7_75t_L g16549 ( 
.A(n_15375),
.Y(n_16549)
);

INVx1_ASAP7_75t_L g16550 ( 
.A(n_15258),
.Y(n_16550)
);

AOI22xp5_ASAP7_75t_L g16551 ( 
.A1(n_15764),
.A2(n_10159),
.B1(n_10137),
.B2(n_9775),
.Y(n_16551)
);

AOI22xp5_ASAP7_75t_L g16552 ( 
.A1(n_15764),
.A2(n_10159),
.B1(n_10137),
.B2(n_9775),
.Y(n_16552)
);

NOR3xp33_ASAP7_75t_L g16553 ( 
.A(n_15280),
.B(n_10023),
.C(n_9993),
.Y(n_16553)
);

NAND2xp5_ASAP7_75t_L g16554 ( 
.A(n_15286),
.B(n_11082),
.Y(n_16554)
);

AND2x2_ASAP7_75t_L g16555 ( 
.A(n_15732),
.B(n_9072),
.Y(n_16555)
);

AND2x2_ASAP7_75t_L g16556 ( 
.A(n_15740),
.B(n_9072),
.Y(n_16556)
);

NAND3xp33_ASAP7_75t_L g16557 ( 
.A(n_15291),
.B(n_9723),
.C(n_10616),
.Y(n_16557)
);

NAND3xp33_ASAP7_75t_L g16558 ( 
.A(n_15294),
.B(n_10616),
.C(n_11985),
.Y(n_16558)
);

NAND2xp5_ASAP7_75t_L g16559 ( 
.A(n_15299),
.B(n_11082),
.Y(n_16559)
);

NAND2xp5_ASAP7_75t_L g16560 ( 
.A(n_15317),
.B(n_11082),
.Y(n_16560)
);

NAND2xp5_ASAP7_75t_L g16561 ( 
.A(n_15321),
.B(n_11082),
.Y(n_16561)
);

NAND2xp5_ASAP7_75t_L g16562 ( 
.A(n_15327),
.B(n_11082),
.Y(n_16562)
);

NAND2xp5_ASAP7_75t_L g16563 ( 
.A(n_15329),
.B(n_11082),
.Y(n_16563)
);

NAND2xp5_ASAP7_75t_L g16564 ( 
.A(n_15330),
.B(n_11082),
.Y(n_16564)
);

NAND2xp5_ASAP7_75t_L g16565 ( 
.A(n_15332),
.B(n_15335),
.Y(n_16565)
);

OAI21xp33_ASAP7_75t_L g16566 ( 
.A1(n_15087),
.A2(n_9582),
.B(n_11610),
.Y(n_16566)
);

AND2x2_ASAP7_75t_L g16567 ( 
.A(n_15743),
.B(n_9072),
.Y(n_16567)
);

AOI21xp5_ASAP7_75t_L g16568 ( 
.A1(n_15833),
.A2(n_12015),
.B(n_11985),
.Y(n_16568)
);

NOR3xp33_ASAP7_75t_L g16569 ( 
.A(n_15342),
.B(n_10023),
.C(n_9993),
.Y(n_16569)
);

AND2x2_ASAP7_75t_L g16570 ( 
.A(n_15448),
.B(n_9072),
.Y(n_16570)
);

OAI221xp5_ASAP7_75t_SL g16571 ( 
.A1(n_15589),
.A2(n_11614),
.B1(n_9294),
.B2(n_9329),
.C(n_9108),
.Y(n_16571)
);

AND2x2_ASAP7_75t_L g16572 ( 
.A(n_15755),
.B(n_15762),
.Y(n_16572)
);

OA21x2_ASAP7_75t_L g16573 ( 
.A1(n_15683),
.A2(n_10913),
.B(n_10905),
.Y(n_16573)
);

INVxp67_ASAP7_75t_L g16574 ( 
.A(n_15141),
.Y(n_16574)
);

NAND3xp33_ASAP7_75t_L g16575 ( 
.A(n_15345),
.B(n_10616),
.C(n_11985),
.Y(n_16575)
);

NAND2xp5_ASAP7_75t_SL g16576 ( 
.A(n_15843),
.B(n_11276),
.Y(n_16576)
);

NAND2xp5_ASAP7_75t_L g16577 ( 
.A(n_15348),
.B(n_11085),
.Y(n_16577)
);

OAI21xp5_ASAP7_75t_SL g16578 ( 
.A1(n_15843),
.A2(n_11616),
.B(n_10038),
.Y(n_16578)
);

NAND2xp5_ASAP7_75t_SL g16579 ( 
.A(n_15729),
.B(n_11469),
.Y(n_16579)
);

NAND2xp5_ASAP7_75t_L g16580 ( 
.A(n_15357),
.B(n_11085),
.Y(n_16580)
);

NAND2xp5_ASAP7_75t_L g16581 ( 
.A(n_15367),
.B(n_11085),
.Y(n_16581)
);

NAND3xp33_ASAP7_75t_L g16582 ( 
.A(n_15397),
.B(n_12015),
.C(n_10807),
.Y(n_16582)
);

AND2x2_ASAP7_75t_L g16583 ( 
.A(n_15755),
.B(n_9072),
.Y(n_16583)
);

AOI221xp5_ASAP7_75t_L g16584 ( 
.A1(n_15405),
.A2(n_11478),
.B1(n_11469),
.B2(n_10942),
.C(n_10110),
.Y(n_16584)
);

AND2x2_ASAP7_75t_L g16585 ( 
.A(n_15762),
.B(n_9072),
.Y(n_16585)
);

NAND2xp5_ASAP7_75t_L g16586 ( 
.A(n_15406),
.B(n_11085),
.Y(n_16586)
);

NAND2xp5_ASAP7_75t_L g16587 ( 
.A(n_15408),
.B(n_11085),
.Y(n_16587)
);

NOR2xp33_ASAP7_75t_L g16588 ( 
.A(n_15399),
.B(n_9072),
.Y(n_16588)
);

AOI221xp5_ASAP7_75t_SL g16589 ( 
.A1(n_15824),
.A2(n_11478),
.B1(n_11469),
.B2(n_10110),
.C(n_10181),
.Y(n_16589)
);

NAND3xp33_ASAP7_75t_L g16590 ( 
.A(n_15411),
.B(n_12015),
.C(n_10807),
.Y(n_16590)
);

NAND2xp5_ASAP7_75t_L g16591 ( 
.A(n_15415),
.B(n_11085),
.Y(n_16591)
);

OAI21xp33_ASAP7_75t_L g16592 ( 
.A1(n_15601),
.A2(n_9582),
.B(n_11616),
.Y(n_16592)
);

NAND2xp5_ASAP7_75t_SL g16593 ( 
.A(n_15729),
.B(n_11478),
.Y(n_16593)
);

AND2x2_ASAP7_75t_L g16594 ( 
.A(n_15773),
.B(n_9072),
.Y(n_16594)
);

NAND2xp5_ASAP7_75t_L g16595 ( 
.A(n_15420),
.B(n_11085),
.Y(n_16595)
);

AND2x2_ASAP7_75t_L g16596 ( 
.A(n_15773),
.B(n_9102),
.Y(n_16596)
);

NAND2xp5_ASAP7_75t_L g16597 ( 
.A(n_15423),
.B(n_11085),
.Y(n_16597)
);

NAND2xp5_ASAP7_75t_L g16598 ( 
.A(n_15434),
.B(n_9046),
.Y(n_16598)
);

NAND2xp5_ASAP7_75t_L g16599 ( 
.A(n_15436),
.B(n_15447),
.Y(n_16599)
);

AND2x2_ASAP7_75t_L g16600 ( 
.A(n_15792),
.B(n_9102),
.Y(n_16600)
);

OA21x2_ASAP7_75t_L g16601 ( 
.A1(n_15684),
.A2(n_15703),
.B(n_15688),
.Y(n_16601)
);

NAND3xp33_ASAP7_75t_L g16602 ( 
.A(n_15453),
.B(n_10807),
.C(n_10805),
.Y(n_16602)
);

NAND3xp33_ASAP7_75t_L g16603 ( 
.A(n_15459),
.B(n_10807),
.C(n_10805),
.Y(n_16603)
);

AND2x2_ASAP7_75t_L g16604 ( 
.A(n_15792),
.B(n_9102),
.Y(n_16604)
);

NAND2xp5_ASAP7_75t_L g16605 ( 
.A(n_15465),
.B(n_9046),
.Y(n_16605)
);

NAND3xp33_ASAP7_75t_L g16606 ( 
.A(n_15482),
.B(n_10807),
.C(n_10805),
.Y(n_16606)
);

NAND4xp25_ASAP7_75t_L g16607 ( 
.A(n_15491),
.B(n_8935),
.C(n_9946),
.D(n_9918),
.Y(n_16607)
);

NAND4xp25_ASAP7_75t_L g16608 ( 
.A(n_15492),
.B(n_9918),
.C(n_9982),
.D(n_9946),
.Y(n_16608)
);

NAND3xp33_ASAP7_75t_L g16609 ( 
.A(n_15504),
.B(n_10807),
.C(n_10805),
.Y(n_16609)
);

NAND3xp33_ASAP7_75t_L g16610 ( 
.A(n_15505),
.B(n_10813),
.C(n_10805),
.Y(n_16610)
);

NAND2xp5_ASAP7_75t_L g16611 ( 
.A(n_15165),
.B(n_9046),
.Y(n_16611)
);

NAND3xp33_ASAP7_75t_L g16612 ( 
.A(n_15212),
.B(n_10813),
.C(n_10805),
.Y(n_16612)
);

AND2x2_ASAP7_75t_L g16613 ( 
.A(n_15495),
.B(n_15503),
.Y(n_16613)
);

AND2x2_ASAP7_75t_L g16614 ( 
.A(n_15628),
.B(n_9102),
.Y(n_16614)
);

NAND3xp33_ASAP7_75t_L g16615 ( 
.A(n_15377),
.B(n_10813),
.C(n_11478),
.Y(n_16615)
);

OAI21xp5_ASAP7_75t_L g16616 ( 
.A1(n_15680),
.A2(n_10774),
.B(n_10771),
.Y(n_16616)
);

AND2x2_ASAP7_75t_SL g16617 ( 
.A(n_15544),
.B(n_9792),
.Y(n_16617)
);

NAND2xp5_ASAP7_75t_L g16618 ( 
.A(n_15381),
.B(n_9046),
.Y(n_16618)
);

NAND2xp5_ASAP7_75t_L g16619 ( 
.A(n_15384),
.B(n_15388),
.Y(n_16619)
);

INVxp67_ASAP7_75t_SL g16620 ( 
.A(n_16125),
.Y(n_16620)
);

AND2x2_ASAP7_75t_L g16621 ( 
.A(n_15993),
.B(n_15631),
.Y(n_16621)
);

NAND2xp5_ASAP7_75t_L g16622 ( 
.A(n_16248),
.B(n_15389),
.Y(n_16622)
);

AND2x2_ASAP7_75t_L g16623 ( 
.A(n_15999),
.B(n_15636),
.Y(n_16623)
);

INVx2_ASAP7_75t_L g16624 ( 
.A(n_15998),
.Y(n_16624)
);

INVx1_ASAP7_75t_L g16625 ( 
.A(n_16007),
.Y(n_16625)
);

HB1xp67_ASAP7_75t_L g16626 ( 
.A(n_16034),
.Y(n_16626)
);

INVx1_ASAP7_75t_L g16627 ( 
.A(n_16373),
.Y(n_16627)
);

INVxp67_ASAP7_75t_L g16628 ( 
.A(n_15880),
.Y(n_16628)
);

AND2x2_ASAP7_75t_L g16629 ( 
.A(n_15927),
.B(n_15643),
.Y(n_16629)
);

NAND2xp5_ASAP7_75t_L g16630 ( 
.A(n_16307),
.B(n_15392),
.Y(n_16630)
);

NAND3xp33_ASAP7_75t_L g16631 ( 
.A(n_15881),
.B(n_15287),
.C(n_15284),
.Y(n_16631)
);

AND2x2_ASAP7_75t_L g16632 ( 
.A(n_15937),
.B(n_15656),
.Y(n_16632)
);

AND2x2_ASAP7_75t_L g16633 ( 
.A(n_16045),
.B(n_15660),
.Y(n_16633)
);

INVx1_ASAP7_75t_L g16634 ( 
.A(n_16076),
.Y(n_16634)
);

NAND2xp5_ASAP7_75t_L g16635 ( 
.A(n_15888),
.B(n_15554),
.Y(n_16635)
);

INVxp67_ASAP7_75t_L g16636 ( 
.A(n_15994),
.Y(n_16636)
);

INVx2_ASAP7_75t_L g16637 ( 
.A(n_16065),
.Y(n_16637)
);

AND2x2_ASAP7_75t_L g16638 ( 
.A(n_16066),
.B(n_15667),
.Y(n_16638)
);

AND2x2_ASAP7_75t_L g16639 ( 
.A(n_15895),
.B(n_15593),
.Y(n_16639)
);

AND2x2_ASAP7_75t_L g16640 ( 
.A(n_16419),
.B(n_16543),
.Y(n_16640)
);

NAND2xp5_ASAP7_75t_L g16641 ( 
.A(n_16095),
.B(n_15528),
.Y(n_16641)
);

AND2x2_ASAP7_75t_L g16642 ( 
.A(n_16043),
.B(n_15599),
.Y(n_16642)
);

AND2x4_ASAP7_75t_L g16643 ( 
.A(n_16238),
.B(n_15652),
.Y(n_16643)
);

NAND2xp5_ASAP7_75t_L g16644 ( 
.A(n_15926),
.B(n_15761),
.Y(n_16644)
);

AND2x2_ASAP7_75t_L g16645 ( 
.A(n_15894),
.B(n_15608),
.Y(n_16645)
);

NAND2xp5_ASAP7_75t_L g16646 ( 
.A(n_15957),
.B(n_15849),
.Y(n_16646)
);

NAND2xp5_ASAP7_75t_L g16647 ( 
.A(n_15946),
.B(n_16006),
.Y(n_16647)
);

OR2x2_ASAP7_75t_L g16648 ( 
.A(n_15896),
.B(n_15464),
.Y(n_16648)
);

HB1xp67_ASAP7_75t_L g16649 ( 
.A(n_16034),
.Y(n_16649)
);

INVxp67_ASAP7_75t_L g16650 ( 
.A(n_16178),
.Y(n_16650)
);

AND2x4_ASAP7_75t_SL g16651 ( 
.A(n_16572),
.B(n_15517),
.Y(n_16651)
);

AND2x4_ASAP7_75t_L g16652 ( 
.A(n_16252),
.B(n_16003),
.Y(n_16652)
);

NAND2xp5_ASAP7_75t_L g16653 ( 
.A(n_16026),
.B(n_15853),
.Y(n_16653)
);

INVx1_ASAP7_75t_L g16654 ( 
.A(n_16324),
.Y(n_16654)
);

NAND2xp5_ASAP7_75t_L g16655 ( 
.A(n_15969),
.B(n_15854),
.Y(n_16655)
);

AND2x4_ASAP7_75t_SL g16656 ( 
.A(n_16473),
.B(n_16488),
.Y(n_16656)
);

INVx2_ASAP7_75t_L g16657 ( 
.A(n_16065),
.Y(n_16657)
);

INVx1_ASAP7_75t_L g16658 ( 
.A(n_16383),
.Y(n_16658)
);

INVx2_ASAP7_75t_L g16659 ( 
.A(n_16082),
.Y(n_16659)
);

BUFx2_ASAP7_75t_L g16660 ( 
.A(n_16082),
.Y(n_16660)
);

OR2x2_ASAP7_75t_L g16661 ( 
.A(n_15979),
.B(n_15109),
.Y(n_16661)
);

INVx1_ASAP7_75t_L g16662 ( 
.A(n_16453),
.Y(n_16662)
);

OR2x2_ASAP7_75t_L g16663 ( 
.A(n_16009),
.B(n_15793),
.Y(n_16663)
);

INVx3_ASAP7_75t_L g16664 ( 
.A(n_16115),
.Y(n_16664)
);

NAND2xp5_ASAP7_75t_L g16665 ( 
.A(n_15970),
.B(n_15855),
.Y(n_16665)
);

INVx1_ASAP7_75t_L g16666 ( 
.A(n_16471),
.Y(n_16666)
);

INVx1_ASAP7_75t_L g16667 ( 
.A(n_16549),
.Y(n_16667)
);

AND2x2_ASAP7_75t_L g16668 ( 
.A(n_16481),
.B(n_15610),
.Y(n_16668)
);

INVx1_ASAP7_75t_L g16669 ( 
.A(n_16601),
.Y(n_16669)
);

HB1xp67_ASAP7_75t_L g16670 ( 
.A(n_16027),
.Y(n_16670)
);

INVx2_ASAP7_75t_L g16671 ( 
.A(n_15951),
.Y(n_16671)
);

AND2x4_ASAP7_75t_L g16672 ( 
.A(n_16407),
.B(n_15454),
.Y(n_16672)
);

NAND2xp5_ASAP7_75t_L g16673 ( 
.A(n_15891),
.B(n_15967),
.Y(n_16673)
);

AND2x2_ASAP7_75t_L g16674 ( 
.A(n_16077),
.B(n_15590),
.Y(n_16674)
);

AND2x2_ASAP7_75t_L g16675 ( 
.A(n_15884),
.B(n_15591),
.Y(n_16675)
);

AND2x2_ASAP7_75t_L g16676 ( 
.A(n_15882),
.B(n_15509),
.Y(n_16676)
);

AND2x2_ASAP7_75t_L g16677 ( 
.A(n_15885),
.B(n_15512),
.Y(n_16677)
);

INVx2_ASAP7_75t_SL g16678 ( 
.A(n_16117),
.Y(n_16678)
);

NAND2xp5_ASAP7_75t_L g16679 ( 
.A(n_16010),
.B(n_15864),
.Y(n_16679)
);

OR2x2_ASAP7_75t_L g16680 ( 
.A(n_16263),
.B(n_15398),
.Y(n_16680)
);

AND2x2_ASAP7_75t_L g16681 ( 
.A(n_15906),
.B(n_15515),
.Y(n_16681)
);

INVx2_ASAP7_75t_L g16682 ( 
.A(n_16352),
.Y(n_16682)
);

NOR2x1_ASAP7_75t_L g16683 ( 
.A(n_16014),
.B(n_15725),
.Y(n_16683)
);

HB1xp67_ASAP7_75t_L g16684 ( 
.A(n_16027),
.Y(n_16684)
);

AND2x4_ASAP7_75t_L g16685 ( 
.A(n_15945),
.B(n_15300),
.Y(n_16685)
);

INVx1_ASAP7_75t_L g16686 ( 
.A(n_16601),
.Y(n_16686)
);

INVx1_ASAP7_75t_L g16687 ( 
.A(n_16550),
.Y(n_16687)
);

AND2x4_ASAP7_75t_L g16688 ( 
.A(n_16024),
.B(n_15334),
.Y(n_16688)
);

INVx1_ASAP7_75t_L g16689 ( 
.A(n_16216),
.Y(n_16689)
);

OR2x2_ASAP7_75t_L g16690 ( 
.A(n_15960),
.B(n_15398),
.Y(n_16690)
);

HB1xp67_ASAP7_75t_L g16691 ( 
.A(n_16105),
.Y(n_16691)
);

INVx1_ASAP7_75t_L g16692 ( 
.A(n_15952),
.Y(n_16692)
);

INVx2_ASAP7_75t_L g16693 ( 
.A(n_16176),
.Y(n_16693)
);

INVx1_ASAP7_75t_L g16694 ( 
.A(n_15909),
.Y(n_16694)
);

INVx1_ASAP7_75t_L g16695 ( 
.A(n_15936),
.Y(n_16695)
);

INVx1_ASAP7_75t_L g16696 ( 
.A(n_16050),
.Y(n_16696)
);

INVx1_ASAP7_75t_L g16697 ( 
.A(n_15916),
.Y(n_16697)
);

INVx2_ASAP7_75t_L g16698 ( 
.A(n_16204),
.Y(n_16698)
);

INVx2_ASAP7_75t_L g16699 ( 
.A(n_16051),
.Y(n_16699)
);

HB1xp67_ASAP7_75t_L g16700 ( 
.A(n_16501),
.Y(n_16700)
);

INVx2_ASAP7_75t_L g16701 ( 
.A(n_16062),
.Y(n_16701)
);

INVx1_ASAP7_75t_L g16702 ( 
.A(n_16255),
.Y(n_16702)
);

AND2x2_ASAP7_75t_L g16703 ( 
.A(n_15925),
.B(n_15919),
.Y(n_16703)
);

HB1xp67_ASAP7_75t_L g16704 ( 
.A(n_15972),
.Y(n_16704)
);

INVx2_ASAP7_75t_L g16705 ( 
.A(n_15987),
.Y(n_16705)
);

AND2x2_ASAP7_75t_L g16706 ( 
.A(n_15908),
.B(n_15457),
.Y(n_16706)
);

AND2x2_ASAP7_75t_L g16707 ( 
.A(n_16033),
.B(n_15767),
.Y(n_16707)
);

INVx2_ASAP7_75t_L g16708 ( 
.A(n_16068),
.Y(n_16708)
);

HB1xp67_ASAP7_75t_L g16709 ( 
.A(n_15988),
.Y(n_16709)
);

HB1xp67_ASAP7_75t_L g16710 ( 
.A(n_15978),
.Y(n_16710)
);

INVx2_ASAP7_75t_L g16711 ( 
.A(n_16119),
.Y(n_16711)
);

NAND2xp5_ASAP7_75t_L g16712 ( 
.A(n_15948),
.B(n_15867),
.Y(n_16712)
);

AND2x2_ASAP7_75t_L g16713 ( 
.A(n_16403),
.B(n_15771),
.Y(n_16713)
);

AND2x4_ASAP7_75t_L g16714 ( 
.A(n_16239),
.B(n_15526),
.Y(n_16714)
);

HB1xp67_ASAP7_75t_L g16715 ( 
.A(n_15981),
.Y(n_16715)
);

AND2x2_ASAP7_75t_L g16716 ( 
.A(n_16368),
.B(n_15779),
.Y(n_16716)
);

INVx1_ASAP7_75t_L g16717 ( 
.A(n_16355),
.Y(n_16717)
);

INVx1_ASAP7_75t_L g16718 ( 
.A(n_16020),
.Y(n_16718)
);

AND2x4_ASAP7_75t_L g16719 ( 
.A(n_16194),
.B(n_15527),
.Y(n_16719)
);

AND2x2_ASAP7_75t_L g16720 ( 
.A(n_16135),
.B(n_15782),
.Y(n_16720)
);

INVx1_ASAP7_75t_L g16721 ( 
.A(n_16025),
.Y(n_16721)
);

NAND2xp5_ASAP7_75t_L g16722 ( 
.A(n_16096),
.B(n_15817),
.Y(n_16722)
);

AND2x2_ASAP7_75t_L g16723 ( 
.A(n_16138),
.B(n_15783),
.Y(n_16723)
);

HB1xp67_ASAP7_75t_L g16724 ( 
.A(n_16316),
.Y(n_16724)
);

INVx2_ASAP7_75t_L g16725 ( 
.A(n_15989),
.Y(n_16725)
);

NAND2xp5_ASAP7_75t_SL g16726 ( 
.A(n_15887),
.B(n_15838),
.Y(n_16726)
);

INVx2_ASAP7_75t_L g16727 ( 
.A(n_16133),
.Y(n_16727)
);

AND2x2_ASAP7_75t_L g16728 ( 
.A(n_15900),
.B(n_15785),
.Y(n_16728)
);

INVx1_ASAP7_75t_L g16729 ( 
.A(n_15986),
.Y(n_16729)
);

NAND2xp5_ASAP7_75t_L g16730 ( 
.A(n_15874),
.B(n_15717),
.Y(n_16730)
);

HB1xp67_ASAP7_75t_L g16731 ( 
.A(n_16320),
.Y(n_16731)
);

AND2x2_ASAP7_75t_L g16732 ( 
.A(n_16435),
.B(n_15796),
.Y(n_16732)
);

INVx2_ASAP7_75t_L g16733 ( 
.A(n_16142),
.Y(n_16733)
);

INVx2_ASAP7_75t_SL g16734 ( 
.A(n_15931),
.Y(n_16734)
);

INVx1_ASAP7_75t_L g16735 ( 
.A(n_15990),
.Y(n_16735)
);

AND2x2_ASAP7_75t_L g16736 ( 
.A(n_16442),
.B(n_16613),
.Y(n_16736)
);

AND2x4_ASAP7_75t_L g16737 ( 
.A(n_16449),
.B(n_15801),
.Y(n_16737)
);

HB1xp67_ASAP7_75t_L g16738 ( 
.A(n_16212),
.Y(n_16738)
);

AND2x2_ASAP7_75t_L g16739 ( 
.A(n_15968),
.B(n_15802),
.Y(n_16739)
);

OR2x2_ASAP7_75t_L g16740 ( 
.A(n_15872),
.B(n_15468),
.Y(n_16740)
);

OR2x2_ASAP7_75t_L g16741 ( 
.A(n_15963),
.B(n_15498),
.Y(n_16741)
);

INVx1_ASAP7_75t_L g16742 ( 
.A(n_16031),
.Y(n_16742)
);

AND2x2_ASAP7_75t_L g16743 ( 
.A(n_15898),
.B(n_15812),
.Y(n_16743)
);

NAND2xp5_ASAP7_75t_L g16744 ( 
.A(n_15878),
.B(n_15718),
.Y(n_16744)
);

AND2x2_ASAP7_75t_L g16745 ( 
.A(n_15869),
.B(n_15813),
.Y(n_16745)
);

OR2x2_ASAP7_75t_L g16746 ( 
.A(n_15964),
.B(n_15499),
.Y(n_16746)
);

INVx2_ASAP7_75t_SL g16747 ( 
.A(n_16074),
.Y(n_16747)
);

INVx1_ASAP7_75t_L g16748 ( 
.A(n_15949),
.Y(n_16748)
);

AND2x2_ASAP7_75t_L g16749 ( 
.A(n_16102),
.B(n_16114),
.Y(n_16749)
);

INVx1_ASAP7_75t_L g16750 ( 
.A(n_15976),
.Y(n_16750)
);

NAND2xp5_ASAP7_75t_L g16751 ( 
.A(n_15879),
.B(n_15804),
.Y(n_16751)
);

INVx1_ASAP7_75t_L g16752 ( 
.A(n_16100),
.Y(n_16752)
);

INVx2_ASAP7_75t_SL g16753 ( 
.A(n_16011),
.Y(n_16753)
);

AND2x2_ASAP7_75t_L g16754 ( 
.A(n_16037),
.B(n_15821),
.Y(n_16754)
);

AND2x2_ASAP7_75t_L g16755 ( 
.A(n_16285),
.B(n_15823),
.Y(n_16755)
);

AND2x2_ASAP7_75t_L g16756 ( 
.A(n_16079),
.B(n_15578),
.Y(n_16756)
);

INVx1_ASAP7_75t_L g16757 ( 
.A(n_16169),
.Y(n_16757)
);

NAND2xp5_ASAP7_75t_L g16758 ( 
.A(n_15928),
.B(n_15805),
.Y(n_16758)
);

AND2x2_ASAP7_75t_L g16759 ( 
.A(n_16040),
.B(n_15581),
.Y(n_16759)
);

NAND2xp5_ASAP7_75t_SL g16760 ( 
.A(n_15876),
.B(n_15838),
.Y(n_16760)
);

INVx2_ASAP7_75t_SL g16761 ( 
.A(n_16417),
.Y(n_16761)
);

OR2x2_ASAP7_75t_L g16762 ( 
.A(n_16380),
.B(n_15501),
.Y(n_16762)
);

AND2x2_ASAP7_75t_L g16763 ( 
.A(n_16121),
.B(n_15585),
.Y(n_16763)
);

NAND4xp25_ASAP7_75t_L g16764 ( 
.A(n_15870),
.B(n_15774),
.C(n_15781),
.D(n_15776),
.Y(n_16764)
);

AND2x2_ASAP7_75t_L g16765 ( 
.A(n_16036),
.B(n_15679),
.Y(n_16765)
);

INVx1_ASAP7_75t_L g16766 ( 
.A(n_16170),
.Y(n_16766)
);

AND2x2_ASAP7_75t_L g16767 ( 
.A(n_15877),
.B(n_15695),
.Y(n_16767)
);

HB1xp67_ASAP7_75t_L g16768 ( 
.A(n_16123),
.Y(n_16768)
);

INVx1_ASAP7_75t_L g16769 ( 
.A(n_16173),
.Y(n_16769)
);

AND2x2_ASAP7_75t_L g16770 ( 
.A(n_15901),
.B(n_15698),
.Y(n_16770)
);

AND2x2_ASAP7_75t_L g16771 ( 
.A(n_16136),
.B(n_15705),
.Y(n_16771)
);

AND2x2_ASAP7_75t_L g16772 ( 
.A(n_15920),
.B(n_15807),
.Y(n_16772)
);

INVx1_ASAP7_75t_L g16773 ( 
.A(n_16174),
.Y(n_16773)
);

INVx1_ASAP7_75t_L g16774 ( 
.A(n_16182),
.Y(n_16774)
);

NOR2xp33_ASAP7_75t_L g16775 ( 
.A(n_16103),
.B(n_15522),
.Y(n_16775)
);

INVx1_ASAP7_75t_L g16776 ( 
.A(n_16184),
.Y(n_16776)
);

NAND2xp5_ASAP7_75t_SL g16777 ( 
.A(n_16124),
.B(n_15830),
.Y(n_16777)
);

INVx1_ASAP7_75t_L g16778 ( 
.A(n_16414),
.Y(n_16778)
);

NAND2xp5_ASAP7_75t_SL g16779 ( 
.A(n_16107),
.B(n_15851),
.Y(n_16779)
);

AND2x2_ASAP7_75t_L g16780 ( 
.A(n_15902),
.B(n_15811),
.Y(n_16780)
);

HB1xp67_ASAP7_75t_L g16781 ( 
.A(n_15959),
.Y(n_16781)
);

INVx1_ASAP7_75t_L g16782 ( 
.A(n_16217),
.Y(n_16782)
);

AND2x2_ASAP7_75t_L g16783 ( 
.A(n_16112),
.B(n_15784),
.Y(n_16783)
);

NOR2xp33_ASAP7_75t_L g16784 ( 
.A(n_16512),
.B(n_15523),
.Y(n_16784)
);

AND2x2_ASAP7_75t_L g16785 ( 
.A(n_16152),
.B(n_15798),
.Y(n_16785)
);

NAND2xp5_ASAP7_75t_L g16786 ( 
.A(n_16057),
.B(n_15800),
.Y(n_16786)
);

AND2x2_ASAP7_75t_L g16787 ( 
.A(n_16126),
.B(n_15334),
.Y(n_16787)
);

OR2x2_ASAP7_75t_L g16788 ( 
.A(n_16244),
.B(n_15506),
.Y(n_16788)
);

AND2x2_ASAP7_75t_L g16789 ( 
.A(n_16128),
.B(n_15858),
.Y(n_16789)
);

INVx1_ASAP7_75t_L g16790 ( 
.A(n_16220),
.Y(n_16790)
);

NOR2xp33_ASAP7_75t_L g16791 ( 
.A(n_16402),
.B(n_15689),
.Y(n_16791)
);

AND2x2_ASAP7_75t_L g16792 ( 
.A(n_16132),
.B(n_15861),
.Y(n_16792)
);

AOI22xp33_ASAP7_75t_L g16793 ( 
.A1(n_15932),
.A2(n_15778),
.B1(n_15704),
.B2(n_15731),
.Y(n_16793)
);

INVxp67_ASAP7_75t_SL g16794 ( 
.A(n_16016),
.Y(n_16794)
);

INVx1_ASAP7_75t_L g16795 ( 
.A(n_16309),
.Y(n_16795)
);

OR2x2_ASAP7_75t_L g16796 ( 
.A(n_16356),
.B(n_15733),
.Y(n_16796)
);

HB1xp67_ASAP7_75t_L g16797 ( 
.A(n_16574),
.Y(n_16797)
);

AND2x2_ASAP7_75t_L g16798 ( 
.A(n_16150),
.B(n_15569),
.Y(n_16798)
);

NAND2x1_ASAP7_75t_SL g16799 ( 
.A(n_15953),
.B(n_15571),
.Y(n_16799)
);

INVx1_ASAP7_75t_L g16800 ( 
.A(n_15973),
.Y(n_16800)
);

INVx2_ASAP7_75t_L g16801 ( 
.A(n_16148),
.Y(n_16801)
);

INVx1_ASAP7_75t_L g16802 ( 
.A(n_16000),
.Y(n_16802)
);

OR2x2_ASAP7_75t_L g16803 ( 
.A(n_15899),
.B(n_15775),
.Y(n_16803)
);

INVx2_ASAP7_75t_L g16804 ( 
.A(n_16384),
.Y(n_16804)
);

INVx1_ASAP7_75t_L g16805 ( 
.A(n_16229),
.Y(n_16805)
);

INVx3_ASAP7_75t_L g16806 ( 
.A(n_16538),
.Y(n_16806)
);

INVx1_ASAP7_75t_SL g16807 ( 
.A(n_15923),
.Y(n_16807)
);

NOR2xp67_ASAP7_75t_L g16808 ( 
.A(n_16039),
.B(n_15574),
.Y(n_16808)
);

NAND2xp5_ASAP7_75t_L g16809 ( 
.A(n_15903),
.B(n_16357),
.Y(n_16809)
);

AND2x2_ASAP7_75t_L g16810 ( 
.A(n_16163),
.B(n_15580),
.Y(n_16810)
);

AND2x2_ASAP7_75t_L g16811 ( 
.A(n_16164),
.B(n_15586),
.Y(n_16811)
);

INVx1_ASAP7_75t_L g16812 ( 
.A(n_15950),
.Y(n_16812)
);

INVxp67_ASAP7_75t_SL g16813 ( 
.A(n_15942),
.Y(n_16813)
);

AND2x2_ASAP7_75t_L g16814 ( 
.A(n_16168),
.B(n_15597),
.Y(n_16814)
);

INVx1_ASAP7_75t_L g16815 ( 
.A(n_16015),
.Y(n_16815)
);

NAND2x1p5_ASAP7_75t_L g16816 ( 
.A(n_16032),
.B(n_8191),
.Y(n_16816)
);

INVx4_ASAP7_75t_L g16817 ( 
.A(n_16353),
.Y(n_16817)
);

AND2x2_ASAP7_75t_L g16818 ( 
.A(n_16425),
.B(n_15604),
.Y(n_16818)
);

AND2x2_ASAP7_75t_L g16819 ( 
.A(n_16298),
.B(n_15614),
.Y(n_16819)
);

HB1xp67_ASAP7_75t_L g16820 ( 
.A(n_16022),
.Y(n_16820)
);

AND2x4_ASAP7_75t_L g16821 ( 
.A(n_15995),
.B(n_15696),
.Y(n_16821)
);

INVx2_ASAP7_75t_L g16822 ( 
.A(n_16384),
.Y(n_16822)
);

AND2x4_ASAP7_75t_L g16823 ( 
.A(n_15971),
.B(n_15933),
.Y(n_16823)
);

OR2x2_ASAP7_75t_L g16824 ( 
.A(n_15965),
.B(n_15696),
.Y(n_16824)
);

AND2x2_ASAP7_75t_L g16825 ( 
.A(n_16246),
.B(n_15616),
.Y(n_16825)
);

INVx2_ASAP7_75t_SL g16826 ( 
.A(n_16617),
.Y(n_16826)
);

OAI22xp5_ASAP7_75t_L g16827 ( 
.A1(n_15873),
.A2(n_15883),
.B1(n_15871),
.B2(n_15929),
.Y(n_16827)
);

AND2x2_ASAP7_75t_L g16828 ( 
.A(n_16091),
.B(n_15618),
.Y(n_16828)
);

INVx1_ASAP7_75t_L g16829 ( 
.A(n_16410),
.Y(n_16829)
);

INVx2_ASAP7_75t_L g16830 ( 
.A(n_16410),
.Y(n_16830)
);

AND2x2_ASAP7_75t_L g16831 ( 
.A(n_16247),
.B(n_16323),
.Y(n_16831)
);

INVx1_ASAP7_75t_L g16832 ( 
.A(n_16412),
.Y(n_16832)
);

INVx1_ASAP7_75t_L g16833 ( 
.A(n_16412),
.Y(n_16833)
);

NOR2x1p5_ASAP7_75t_L g16834 ( 
.A(n_15922),
.B(n_15910),
.Y(n_16834)
);

INVx4_ASAP7_75t_L g16835 ( 
.A(n_16504),
.Y(n_16835)
);

INVx1_ASAP7_75t_L g16836 ( 
.A(n_16565),
.Y(n_16836)
);

NAND2xp5_ASAP7_75t_L g16837 ( 
.A(n_15930),
.B(n_15626),
.Y(n_16837)
);

INVx2_ASAP7_75t_SL g16838 ( 
.A(n_16161),
.Y(n_16838)
);

INVxp67_ASAP7_75t_L g16839 ( 
.A(n_15958),
.Y(n_16839)
);

INVx2_ASAP7_75t_L g16840 ( 
.A(n_16420),
.Y(n_16840)
);

INVx4_ASAP7_75t_L g16841 ( 
.A(n_16505),
.Y(n_16841)
);

AND2x2_ASAP7_75t_L g16842 ( 
.A(n_16393),
.B(n_15627),
.Y(n_16842)
);

INVx1_ASAP7_75t_L g16843 ( 
.A(n_16599),
.Y(n_16843)
);

INVx1_ASAP7_75t_L g16844 ( 
.A(n_16619),
.Y(n_16844)
);

AND2x2_ASAP7_75t_L g16845 ( 
.A(n_16396),
.B(n_15630),
.Y(n_16845)
);

AND2x2_ASAP7_75t_L g16846 ( 
.A(n_16399),
.B(n_15635),
.Y(n_16846)
);

INVx1_ASAP7_75t_L g16847 ( 
.A(n_16153),
.Y(n_16847)
);

AND2x2_ASAP7_75t_L g16848 ( 
.A(n_16371),
.B(n_15780),
.Y(n_16848)
);

INVx1_ASAP7_75t_L g16849 ( 
.A(n_16154),
.Y(n_16849)
);

AND2x2_ASAP7_75t_L g16850 ( 
.A(n_16388),
.B(n_15820),
.Y(n_16850)
);

INVx2_ASAP7_75t_L g16851 ( 
.A(n_16162),
.Y(n_16851)
);

BUFx3_ASAP7_75t_L g16852 ( 
.A(n_15974),
.Y(n_16852)
);

AND2x4_ASAP7_75t_L g16853 ( 
.A(n_15975),
.B(n_10539),
.Y(n_16853)
);

OR2x2_ASAP7_75t_L g16854 ( 
.A(n_15966),
.B(n_16111),
.Y(n_16854)
);

INVx2_ASAP7_75t_L g16855 ( 
.A(n_16408),
.Y(n_16855)
);

AND2x2_ASAP7_75t_L g16856 ( 
.A(n_16325),
.B(n_16328),
.Y(n_16856)
);

INVxp67_ASAP7_75t_SL g16857 ( 
.A(n_16048),
.Y(n_16857)
);

INVx2_ASAP7_75t_L g16858 ( 
.A(n_16594),
.Y(n_16858)
);

AND2x2_ASAP7_75t_L g16859 ( 
.A(n_16330),
.B(n_15860),
.Y(n_16859)
);

AND2x2_ASAP7_75t_L g16860 ( 
.A(n_16344),
.B(n_9102),
.Y(n_16860)
);

INVx1_ASAP7_75t_L g16861 ( 
.A(n_15983),
.Y(n_16861)
);

INVx2_ASAP7_75t_L g16862 ( 
.A(n_16596),
.Y(n_16862)
);

AND2x2_ASAP7_75t_L g16863 ( 
.A(n_16349),
.B(n_9102),
.Y(n_16863)
);

INVxp67_ASAP7_75t_SL g16864 ( 
.A(n_16005),
.Y(n_16864)
);

AND2x2_ASAP7_75t_L g16865 ( 
.A(n_16366),
.B(n_9102),
.Y(n_16865)
);

INVx2_ASAP7_75t_L g16866 ( 
.A(n_16600),
.Y(n_16866)
);

HB1xp67_ASAP7_75t_L g16867 ( 
.A(n_16023),
.Y(n_16867)
);

HB1xp67_ASAP7_75t_L g16868 ( 
.A(n_16070),
.Y(n_16868)
);

INVx2_ASAP7_75t_L g16869 ( 
.A(n_16604),
.Y(n_16869)
);

INVx1_ASAP7_75t_L g16870 ( 
.A(n_15985),
.Y(n_16870)
);

INVx1_ASAP7_75t_L g16871 ( 
.A(n_16240),
.Y(n_16871)
);

AND2x4_ASAP7_75t_L g16872 ( 
.A(n_16406),
.B(n_10539),
.Y(n_16872)
);

NAND2xp5_ASAP7_75t_L g16873 ( 
.A(n_16054),
.B(n_9046),
.Y(n_16873)
);

OR2x2_ASAP7_75t_L g16874 ( 
.A(n_15954),
.B(n_11452),
.Y(n_16874)
);

NAND2xp5_ASAP7_75t_L g16875 ( 
.A(n_15938),
.B(n_9171),
.Y(n_16875)
);

INVx1_ASAP7_75t_L g16876 ( 
.A(n_16235),
.Y(n_16876)
);

NAND2xp5_ASAP7_75t_L g16877 ( 
.A(n_15939),
.B(n_9171),
.Y(n_16877)
);

OAI22xp5_ASAP7_75t_L g16878 ( 
.A1(n_15914),
.A2(n_10048),
.B1(n_10110),
.B2(n_10036),
.Y(n_16878)
);

BUFx2_ASAP7_75t_L g16879 ( 
.A(n_16179),
.Y(n_16879)
);

INVx1_ASAP7_75t_L g16880 ( 
.A(n_16237),
.Y(n_16880)
);

INVx1_ASAP7_75t_L g16881 ( 
.A(n_16573),
.Y(n_16881)
);

INVx3_ASAP7_75t_L g16882 ( 
.A(n_16175),
.Y(n_16882)
);

INVx4_ASAP7_75t_L g16883 ( 
.A(n_16530),
.Y(n_16883)
);

BUFx2_ASAP7_75t_L g16884 ( 
.A(n_16166),
.Y(n_16884)
);

NOR2x1_ASAP7_75t_L g16885 ( 
.A(n_16200),
.B(n_13206),
.Y(n_16885)
);

BUFx2_ASAP7_75t_L g16886 ( 
.A(n_16166),
.Y(n_16886)
);

INVx2_ASAP7_75t_L g16887 ( 
.A(n_16583),
.Y(n_16887)
);

INVx1_ASAP7_75t_L g16888 ( 
.A(n_16573),
.Y(n_16888)
);

INVx1_ASAP7_75t_L g16889 ( 
.A(n_16109),
.Y(n_16889)
);

INVx1_ASAP7_75t_L g16890 ( 
.A(n_16181),
.Y(n_16890)
);

AND2x4_ASAP7_75t_L g16891 ( 
.A(n_16008),
.B(n_10539),
.Y(n_16891)
);

INVx1_ASAP7_75t_L g16892 ( 
.A(n_16181),
.Y(n_16892)
);

INVx3_ASAP7_75t_L g16893 ( 
.A(n_16228),
.Y(n_16893)
);

INVx2_ASAP7_75t_L g16894 ( 
.A(n_16585),
.Y(n_16894)
);

AND2x2_ASAP7_75t_L g16895 ( 
.A(n_16157),
.B(n_16284),
.Y(n_16895)
);

AND2x2_ASAP7_75t_L g16896 ( 
.A(n_15935),
.B(n_16274),
.Y(n_16896)
);

INVx2_ASAP7_75t_L g16897 ( 
.A(n_16544),
.Y(n_16897)
);

AND2x2_ASAP7_75t_L g16898 ( 
.A(n_16281),
.B(n_9102),
.Y(n_16898)
);

AND2x2_ASAP7_75t_L g16899 ( 
.A(n_16283),
.B(n_9172),
.Y(n_16899)
);

OR2x2_ASAP7_75t_L g16900 ( 
.A(n_15956),
.B(n_11452),
.Y(n_16900)
);

AND2x4_ASAP7_75t_L g16901 ( 
.A(n_16071),
.B(n_10539),
.Y(n_16901)
);

AND2x2_ASAP7_75t_L g16902 ( 
.A(n_16017),
.B(n_16021),
.Y(n_16902)
);

AND2x2_ASAP7_75t_L g16903 ( 
.A(n_16495),
.B(n_9172),
.Y(n_16903)
);

NAND2x1p5_ASAP7_75t_L g16904 ( 
.A(n_16075),
.B(n_8191),
.Y(n_16904)
);

INVx1_ASAP7_75t_L g16905 ( 
.A(n_16127),
.Y(n_16905)
);

AND2x2_ASAP7_75t_L g16906 ( 
.A(n_16192),
.B(n_9172),
.Y(n_16906)
);

AND2x2_ASAP7_75t_L g16907 ( 
.A(n_16195),
.B(n_9172),
.Y(n_16907)
);

AND2x2_ASAP7_75t_L g16908 ( 
.A(n_16199),
.B(n_9172),
.Y(n_16908)
);

NAND2xp5_ASAP7_75t_L g16909 ( 
.A(n_16431),
.B(n_9171),
.Y(n_16909)
);

AND2x2_ASAP7_75t_L g16910 ( 
.A(n_16201),
.B(n_9172),
.Y(n_16910)
);

INVx2_ASAP7_75t_L g16911 ( 
.A(n_16230),
.Y(n_16911)
);

INVx1_ASAP7_75t_L g16912 ( 
.A(n_16139),
.Y(n_16912)
);

AND2x2_ASAP7_75t_L g16913 ( 
.A(n_16203),
.B(n_9172),
.Y(n_16913)
);

INVx2_ASAP7_75t_L g16914 ( 
.A(n_16231),
.Y(n_16914)
);

INVx1_ASAP7_75t_L g16915 ( 
.A(n_16141),
.Y(n_16915)
);

INVx2_ASAP7_75t_L g16916 ( 
.A(n_16234),
.Y(n_16916)
);

NAND2xp5_ASAP7_75t_L g16917 ( 
.A(n_15890),
.B(n_9171),
.Y(n_16917)
);

AND2x4_ASAP7_75t_L g16918 ( 
.A(n_16078),
.B(n_16083),
.Y(n_16918)
);

INVx2_ASAP7_75t_L g16919 ( 
.A(n_16243),
.Y(n_16919)
);

AND2x2_ASAP7_75t_L g16920 ( 
.A(n_16213),
.B(n_9172),
.Y(n_16920)
);

HB1xp67_ASAP7_75t_L g16921 ( 
.A(n_16073),
.Y(n_16921)
);

INVx1_ASAP7_75t_L g16922 ( 
.A(n_16145),
.Y(n_16922)
);

OR2x2_ASAP7_75t_L g16923 ( 
.A(n_16089),
.B(n_11452),
.Y(n_16923)
);

AND2x2_ASAP7_75t_L g16924 ( 
.A(n_15996),
.B(n_10539),
.Y(n_16924)
);

NAND2xp5_ASAP7_75t_L g16925 ( 
.A(n_16053),
.B(n_9171),
.Y(n_16925)
);

INVx2_ASAP7_75t_L g16926 ( 
.A(n_16451),
.Y(n_16926)
);

AND2x2_ASAP7_75t_L g16927 ( 
.A(n_16004),
.B(n_10539),
.Y(n_16927)
);

INVx2_ASAP7_75t_L g16928 ( 
.A(n_16456),
.Y(n_16928)
);

NAND2xp5_ASAP7_75t_L g16929 ( 
.A(n_15897),
.B(n_11478),
.Y(n_16929)
);

HB1xp67_ASAP7_75t_L g16930 ( 
.A(n_15997),
.Y(n_16930)
);

BUFx2_ASAP7_75t_L g16931 ( 
.A(n_15955),
.Y(n_16931)
);

AND2x4_ASAP7_75t_L g16932 ( 
.A(n_16249),
.B(n_10539),
.Y(n_16932)
);

INVx1_ASAP7_75t_L g16933 ( 
.A(n_16158),
.Y(n_16933)
);

INVx1_ASAP7_75t_L g16934 ( 
.A(n_16160),
.Y(n_16934)
);

INVx1_ASAP7_75t_L g16935 ( 
.A(n_16188),
.Y(n_16935)
);

INVx3_ASAP7_75t_L g16936 ( 
.A(n_16503),
.Y(n_16936)
);

AND2x2_ASAP7_75t_L g16937 ( 
.A(n_16313),
.B(n_10598),
.Y(n_16937)
);

OR2x2_ASAP7_75t_L g16938 ( 
.A(n_16193),
.B(n_11452),
.Y(n_16938)
);

INVx1_ASAP7_75t_L g16939 ( 
.A(n_16197),
.Y(n_16939)
);

HB1xp67_ASAP7_75t_L g16940 ( 
.A(n_16013),
.Y(n_16940)
);

INVx2_ASAP7_75t_L g16941 ( 
.A(n_16457),
.Y(n_16941)
);

INVx1_ASAP7_75t_SL g16942 ( 
.A(n_16524),
.Y(n_16942)
);

NAND2xp5_ASAP7_75t_L g16943 ( 
.A(n_15984),
.B(n_11478),
.Y(n_16943)
);

OR2x2_ASAP7_75t_L g16944 ( 
.A(n_16202),
.B(n_11452),
.Y(n_16944)
);

AND2x2_ASAP7_75t_L g16945 ( 
.A(n_16250),
.B(n_10598),
.Y(n_16945)
);

OR2x2_ASAP7_75t_L g16946 ( 
.A(n_16208),
.B(n_11452),
.Y(n_16946)
);

HB1xp67_ASAP7_75t_L g16947 ( 
.A(n_15915),
.Y(n_16947)
);

INVx2_ASAP7_75t_L g16948 ( 
.A(n_16458),
.Y(n_16948)
);

INVx1_ASAP7_75t_L g16949 ( 
.A(n_16209),
.Y(n_16949)
);

INVx1_ASAP7_75t_L g16950 ( 
.A(n_16227),
.Y(n_16950)
);

INVx3_ASAP7_75t_L g16951 ( 
.A(n_16470),
.Y(n_16951)
);

NAND4xp25_ASAP7_75t_L g16952 ( 
.A(n_16439),
.B(n_9946),
.C(n_9982),
.D(n_9918),
.Y(n_16952)
);

AND2x2_ASAP7_75t_L g16953 ( 
.A(n_16358),
.B(n_10598),
.Y(n_16953)
);

HB1xp67_ASAP7_75t_L g16954 ( 
.A(n_16256),
.Y(n_16954)
);

AOI22xp33_ASAP7_75t_L g16955 ( 
.A1(n_15886),
.A2(n_10897),
.B1(n_11172),
.B2(n_11169),
.Y(n_16955)
);

INVx1_ASAP7_75t_L g16956 ( 
.A(n_16269),
.Y(n_16956)
);

INVx1_ASAP7_75t_L g16957 ( 
.A(n_16271),
.Y(n_16957)
);

OR2x2_ASAP7_75t_L g16958 ( 
.A(n_15961),
.B(n_11605),
.Y(n_16958)
);

AND2x2_ASAP7_75t_L g16959 ( 
.A(n_16428),
.B(n_10598),
.Y(n_16959)
);

AND2x2_ASAP7_75t_L g16960 ( 
.A(n_16430),
.B(n_10598),
.Y(n_16960)
);

INVx2_ASAP7_75t_L g16961 ( 
.A(n_16437),
.Y(n_16961)
);

INVx1_ASAP7_75t_L g16962 ( 
.A(n_16272),
.Y(n_16962)
);

INVx1_ASAP7_75t_L g16963 ( 
.A(n_16277),
.Y(n_16963)
);

OR2x2_ASAP7_75t_L g16964 ( 
.A(n_16149),
.B(n_16278),
.Y(n_16964)
);

AND2x2_ASAP7_75t_L g16965 ( 
.A(n_16440),
.B(n_10598),
.Y(n_16965)
);

NAND2xp5_ASAP7_75t_SL g16966 ( 
.A(n_16359),
.B(n_10132),
.Y(n_16966)
);

INVx2_ASAP7_75t_L g16967 ( 
.A(n_16443),
.Y(n_16967)
);

AND2x2_ASAP7_75t_L g16968 ( 
.A(n_16447),
.B(n_10598),
.Y(n_16968)
);

NAND2xp5_ASAP7_75t_L g16969 ( 
.A(n_15941),
.B(n_11013),
.Y(n_16969)
);

AND2x2_ASAP7_75t_L g16970 ( 
.A(n_16484),
.B(n_11605),
.Y(n_16970)
);

INVx2_ASAP7_75t_L g16971 ( 
.A(n_16513),
.Y(n_16971)
);

CKINVDCx5p33_ASAP7_75t_R g16972 ( 
.A(n_16386),
.Y(n_16972)
);

AND2x2_ASAP7_75t_L g16973 ( 
.A(n_16177),
.B(n_11605),
.Y(n_16973)
);

HB1xp67_ASAP7_75t_L g16974 ( 
.A(n_16392),
.Y(n_16974)
);

INVx1_ASAP7_75t_L g16975 ( 
.A(n_16279),
.Y(n_16975)
);

BUFx2_ASAP7_75t_L g16976 ( 
.A(n_16183),
.Y(n_16976)
);

NAND2xp5_ASAP7_75t_L g16977 ( 
.A(n_16156),
.B(n_11013),
.Y(n_16977)
);

AND2x2_ASAP7_75t_L g16978 ( 
.A(n_16482),
.B(n_16029),
.Y(n_16978)
);

NAND2xp5_ASAP7_75t_L g16979 ( 
.A(n_15892),
.B(n_11013),
.Y(n_16979)
);

HB1xp67_ASAP7_75t_L g16980 ( 
.A(n_16104),
.Y(n_16980)
);

OR2x2_ASAP7_75t_L g16981 ( 
.A(n_16280),
.B(n_11605),
.Y(n_16981)
);

NOR2x1_ASAP7_75t_L g16982 ( 
.A(n_16012),
.B(n_13206),
.Y(n_16982)
);

AND2x2_ASAP7_75t_L g16983 ( 
.A(n_16046),
.B(n_11605),
.Y(n_16983)
);

OR2x2_ASAP7_75t_L g16984 ( 
.A(n_16172),
.B(n_11605),
.Y(n_16984)
);

BUFx3_ASAP7_75t_L g16985 ( 
.A(n_16052),
.Y(n_16985)
);

OR2x2_ASAP7_75t_L g16986 ( 
.A(n_16055),
.B(n_11605),
.Y(n_16986)
);

HB1xp67_ASAP7_75t_SL g16987 ( 
.A(n_16433),
.Y(n_16987)
);

INVx1_ASAP7_75t_L g16988 ( 
.A(n_16378),
.Y(n_16988)
);

INVx3_ASAP7_75t_SL g16989 ( 
.A(n_16189),
.Y(n_16989)
);

NAND2xp5_ASAP7_75t_L g16990 ( 
.A(n_15962),
.B(n_11013),
.Y(n_16990)
);

INVx1_ASAP7_75t_L g16991 ( 
.A(n_16379),
.Y(n_16991)
);

INVx2_ASAP7_75t_L g16992 ( 
.A(n_16518),
.Y(n_16992)
);

OR2x2_ASAP7_75t_L g16993 ( 
.A(n_16056),
.B(n_11605),
.Y(n_16993)
);

INVx1_ASAP7_75t_L g16994 ( 
.A(n_16381),
.Y(n_16994)
);

INVx2_ASAP7_75t_L g16995 ( 
.A(n_16547),
.Y(n_16995)
);

INVx1_ASAP7_75t_L g16996 ( 
.A(n_16390),
.Y(n_16996)
);

AND2x2_ASAP7_75t_L g16997 ( 
.A(n_16060),
.B(n_9918),
.Y(n_16997)
);

BUFx2_ASAP7_75t_L g16998 ( 
.A(n_15889),
.Y(n_16998)
);

INVxp67_ASAP7_75t_L g16999 ( 
.A(n_16434),
.Y(n_16999)
);

INVx2_ASAP7_75t_L g17000 ( 
.A(n_16479),
.Y(n_17000)
);

INVx1_ASAP7_75t_L g17001 ( 
.A(n_16391),
.Y(n_17001)
);

INVx2_ASAP7_75t_L g17002 ( 
.A(n_16531),
.Y(n_17002)
);

AND2x2_ASAP7_75t_L g17003 ( 
.A(n_16063),
.B(n_16067),
.Y(n_17003)
);

INVx1_ASAP7_75t_L g17004 ( 
.A(n_16394),
.Y(n_17004)
);

INVx1_ASAP7_75t_L g17005 ( 
.A(n_16265),
.Y(n_17005)
);

INVx2_ASAP7_75t_L g17006 ( 
.A(n_16480),
.Y(n_17006)
);

AND2x2_ASAP7_75t_L g17007 ( 
.A(n_16069),
.B(n_9918),
.Y(n_17007)
);

INVx1_ASAP7_75t_L g17008 ( 
.A(n_16268),
.Y(n_17008)
);

AND2x4_ASAP7_75t_L g17009 ( 
.A(n_16144),
.B(n_11013),
.Y(n_17009)
);

INVx1_ASAP7_75t_L g17010 ( 
.A(n_16261),
.Y(n_17010)
);

AND2x2_ASAP7_75t_L g17011 ( 
.A(n_16147),
.B(n_9946),
.Y(n_17011)
);

INVx1_ASAP7_75t_L g17012 ( 
.A(n_16260),
.Y(n_17012)
);

INVx2_ASAP7_75t_L g17013 ( 
.A(n_16462),
.Y(n_17013)
);

INVx1_ASAP7_75t_L g17014 ( 
.A(n_16374),
.Y(n_17014)
);

AND2x2_ASAP7_75t_L g17015 ( 
.A(n_16520),
.B(n_9946),
.Y(n_17015)
);

AND2x2_ASAP7_75t_L g17016 ( 
.A(n_16522),
.B(n_9946),
.Y(n_17016)
);

INVx1_ASAP7_75t_L g17017 ( 
.A(n_16253),
.Y(n_17017)
);

AND2x2_ASAP7_75t_L g17018 ( 
.A(n_16448),
.B(n_9982),
.Y(n_17018)
);

INVx1_ASAP7_75t_L g17019 ( 
.A(n_16245),
.Y(n_17019)
);

INVx1_ASAP7_75t_L g17020 ( 
.A(n_16288),
.Y(n_17020)
);

INVx2_ASAP7_75t_L g17021 ( 
.A(n_16465),
.Y(n_17021)
);

INVx1_ASAP7_75t_L g17022 ( 
.A(n_16291),
.Y(n_17022)
);

AND2x2_ASAP7_75t_L g17023 ( 
.A(n_16438),
.B(n_9982),
.Y(n_17023)
);

AND2x2_ASAP7_75t_L g17024 ( 
.A(n_16293),
.B(n_9982),
.Y(n_17024)
);

INVx4_ASAP7_75t_L g17025 ( 
.A(n_16299),
.Y(n_17025)
);

BUFx3_ASAP7_75t_L g17026 ( 
.A(n_16092),
.Y(n_17026)
);

HB1xp67_ASAP7_75t_L g17027 ( 
.A(n_16196),
.Y(n_17027)
);

OR2x2_ASAP7_75t_L g17028 ( 
.A(n_16097),
.B(n_10787),
.Y(n_17028)
);

INVx1_ASAP7_75t_L g17029 ( 
.A(n_16474),
.Y(n_17029)
);

INVx1_ASAP7_75t_L g17030 ( 
.A(n_16485),
.Y(n_17030)
);

AND2x2_ASAP7_75t_L g17031 ( 
.A(n_16467),
.B(n_9982),
.Y(n_17031)
);

INVx2_ASAP7_75t_L g17032 ( 
.A(n_16468),
.Y(n_17032)
);

AND2x2_ASAP7_75t_L g17033 ( 
.A(n_16322),
.B(n_9990),
.Y(n_17033)
);

AND2x2_ASAP7_75t_L g17034 ( 
.A(n_16493),
.B(n_9990),
.Y(n_17034)
);

OR2x2_ASAP7_75t_L g17035 ( 
.A(n_16376),
.B(n_10787),
.Y(n_17035)
);

NOR2xp33_ASAP7_75t_L g17036 ( 
.A(n_15921),
.B(n_10137),
.Y(n_17036)
);

NAND2xp5_ASAP7_75t_L g17037 ( 
.A(n_15917),
.B(n_15893),
.Y(n_17037)
);

INVx2_ASAP7_75t_L g17038 ( 
.A(n_16494),
.Y(n_17038)
);

AND2x2_ASAP7_75t_L g17039 ( 
.A(n_16398),
.B(n_9990),
.Y(n_17039)
);

HB1xp67_ASAP7_75t_L g17040 ( 
.A(n_16215),
.Y(n_17040)
);

INVx1_ASAP7_75t_L g17041 ( 
.A(n_16486),
.Y(n_17041)
);

OR2x2_ASAP7_75t_L g17042 ( 
.A(n_16526),
.B(n_10787),
.Y(n_17042)
);

INVx2_ASAP7_75t_L g17043 ( 
.A(n_16570),
.Y(n_17043)
);

AND2x2_ASAP7_75t_L g17044 ( 
.A(n_16401),
.B(n_9990),
.Y(n_17044)
);

OR2x2_ASAP7_75t_L g17045 ( 
.A(n_16527),
.B(n_10787),
.Y(n_17045)
);

INVx2_ASAP7_75t_SL g17046 ( 
.A(n_16264),
.Y(n_17046)
);

INVx2_ASAP7_75t_L g17047 ( 
.A(n_16483),
.Y(n_17047)
);

BUFx3_ASAP7_75t_L g17048 ( 
.A(n_16290),
.Y(n_17048)
);

NOR2xp33_ASAP7_75t_L g17049 ( 
.A(n_15992),
.B(n_10137),
.Y(n_17049)
);

INVx1_ASAP7_75t_L g17050 ( 
.A(n_16487),
.Y(n_17050)
);

NAND2x1_ASAP7_75t_L g17051 ( 
.A(n_16521),
.B(n_13212),
.Y(n_17051)
);

OR2x2_ASAP7_75t_L g17052 ( 
.A(n_16529),
.B(n_10787),
.Y(n_17052)
);

OR2x2_ASAP7_75t_L g17053 ( 
.A(n_16532),
.B(n_10787),
.Y(n_17053)
);

INVx2_ASAP7_75t_L g17054 ( 
.A(n_16555),
.Y(n_17054)
);

INVx1_ASAP7_75t_L g17055 ( 
.A(n_16490),
.Y(n_17055)
);

NOR2x1_ASAP7_75t_L g17056 ( 
.A(n_15905),
.B(n_13212),
.Y(n_17056)
);

INVx2_ASAP7_75t_SL g17057 ( 
.A(n_16275),
.Y(n_17057)
);

NAND2xp5_ASAP7_75t_L g17058 ( 
.A(n_16099),
.B(n_11013),
.Y(n_17058)
);

INVx1_ASAP7_75t_L g17059 ( 
.A(n_16496),
.Y(n_17059)
);

INVx1_ASAP7_75t_L g17060 ( 
.A(n_16498),
.Y(n_17060)
);

INVx1_ASAP7_75t_L g17061 ( 
.A(n_16502),
.Y(n_17061)
);

INVx2_ASAP7_75t_L g17062 ( 
.A(n_16556),
.Y(n_17062)
);

INVx1_ASAP7_75t_L g17063 ( 
.A(n_16506),
.Y(n_17063)
);

AND2x4_ASAP7_75t_L g17064 ( 
.A(n_16310),
.B(n_11013),
.Y(n_17064)
);

INVx2_ASAP7_75t_L g17065 ( 
.A(n_16567),
.Y(n_17065)
);

AND2x2_ASAP7_75t_L g17066 ( 
.A(n_16413),
.B(n_9990),
.Y(n_17066)
);

INVx1_ASAP7_75t_L g17067 ( 
.A(n_16510),
.Y(n_17067)
);

INVx2_ASAP7_75t_L g17068 ( 
.A(n_16331),
.Y(n_17068)
);

NAND2xp67_ASAP7_75t_L g17069 ( 
.A(n_16509),
.B(n_9792),
.Y(n_17069)
);

NAND2xp5_ASAP7_75t_SL g17070 ( 
.A(n_16131),
.B(n_10132),
.Y(n_17070)
);

INVx1_ASAP7_75t_L g17071 ( 
.A(n_16514),
.Y(n_17071)
);

AND2x4_ASAP7_75t_L g17072 ( 
.A(n_16354),
.B(n_11013),
.Y(n_17072)
);

INVx2_ASAP7_75t_SL g17073 ( 
.A(n_16375),
.Y(n_17073)
);

INVx1_ASAP7_75t_L g17074 ( 
.A(n_16516),
.Y(n_17074)
);

AND2x2_ASAP7_75t_L g17075 ( 
.A(n_16416),
.B(n_9990),
.Y(n_17075)
);

INVx2_ASAP7_75t_SL g17076 ( 
.A(n_16426),
.Y(n_17076)
);

HB1xp67_ASAP7_75t_L g17077 ( 
.A(n_16241),
.Y(n_17077)
);

AND2x2_ASAP7_75t_SL g17078 ( 
.A(n_16087),
.B(n_9792),
.Y(n_17078)
);

AND2x2_ASAP7_75t_L g17079 ( 
.A(n_16421),
.B(n_10004),
.Y(n_17079)
);

INVx1_ASAP7_75t_L g17080 ( 
.A(n_16519),
.Y(n_17080)
);

NAND2xp5_ASAP7_75t_L g17081 ( 
.A(n_16588),
.B(n_11022),
.Y(n_17081)
);

INVx1_ASAP7_75t_L g17082 ( 
.A(n_16523),
.Y(n_17082)
);

INVx1_ASAP7_75t_L g17083 ( 
.A(n_16598),
.Y(n_17083)
);

AND2x2_ASAP7_75t_L g17084 ( 
.A(n_16436),
.B(n_10004),
.Y(n_17084)
);

AND2x2_ASAP7_75t_L g17085 ( 
.A(n_16108),
.B(n_10004),
.Y(n_17085)
);

AND2x2_ASAP7_75t_L g17086 ( 
.A(n_16333),
.B(n_10004),
.Y(n_17086)
);

INVx1_ASAP7_75t_L g17087 ( 
.A(n_16605),
.Y(n_17087)
);

INVx1_ASAP7_75t_L g17088 ( 
.A(n_16618),
.Y(n_17088)
);

INVx2_ASAP7_75t_L g17089 ( 
.A(n_16499),
.Y(n_17089)
);

OR2x2_ASAP7_75t_L g17090 ( 
.A(n_16535),
.B(n_10787),
.Y(n_17090)
);

INVx1_ASAP7_75t_L g17091 ( 
.A(n_16294),
.Y(n_17091)
);

INVx1_ASAP7_75t_L g17092 ( 
.A(n_16295),
.Y(n_17092)
);

NOR2x1p5_ASAP7_75t_L g17093 ( 
.A(n_16500),
.B(n_9092),
.Y(n_17093)
);

INVx1_ASAP7_75t_L g17094 ( 
.A(n_16300),
.Y(n_17094)
);

INVx1_ASAP7_75t_L g17095 ( 
.A(n_16301),
.Y(n_17095)
);

NAND2xp5_ASAP7_75t_L g17096 ( 
.A(n_15912),
.B(n_11022),
.Y(n_17096)
);

HB1xp67_ASAP7_75t_L g17097 ( 
.A(n_16541),
.Y(n_17097)
);

AND2x2_ASAP7_75t_L g17098 ( 
.A(n_16343),
.B(n_10004),
.Y(n_17098)
);

INVx2_ASAP7_75t_L g17099 ( 
.A(n_16326),
.Y(n_17099)
);

AND2x2_ASAP7_75t_L g17100 ( 
.A(n_16347),
.B(n_10004),
.Y(n_17100)
);

AND2x2_ASAP7_75t_L g17101 ( 
.A(n_16350),
.B(n_10056),
.Y(n_17101)
);

HB1xp67_ASAP7_75t_L g17102 ( 
.A(n_15924),
.Y(n_17102)
);

INVx1_ASAP7_75t_L g17103 ( 
.A(n_16304),
.Y(n_17103)
);

INVx1_ASAP7_75t_L g17104 ( 
.A(n_16351),
.Y(n_17104)
);

INVx2_ASAP7_75t_L g17105 ( 
.A(n_16327),
.Y(n_17105)
);

AND2x2_ASAP7_75t_L g17106 ( 
.A(n_16311),
.B(n_10056),
.Y(n_17106)
);

INVx2_ASAP7_75t_L g17107 ( 
.A(n_16332),
.Y(n_17107)
);

AND2x2_ASAP7_75t_L g17108 ( 
.A(n_16317),
.B(n_10056),
.Y(n_17108)
);

INVx1_ASAP7_75t_L g17109 ( 
.A(n_16611),
.Y(n_17109)
);

AND2x4_ASAP7_75t_SL g17110 ( 
.A(n_16525),
.B(n_7831),
.Y(n_17110)
);

NAND2xp5_ASAP7_75t_L g17111 ( 
.A(n_16382),
.B(n_16002),
.Y(n_17111)
);

INVx1_ASAP7_75t_L g17112 ( 
.A(n_16452),
.Y(n_17112)
);

CKINVDCx20_ASAP7_75t_R g17113 ( 
.A(n_16489),
.Y(n_17113)
);

AND2x4_ASAP7_75t_L g17114 ( 
.A(n_16576),
.B(n_16579),
.Y(n_17114)
);

AND2x2_ASAP7_75t_L g17115 ( 
.A(n_16312),
.B(n_10056),
.Y(n_17115)
);

INVx1_ASAP7_75t_L g17116 ( 
.A(n_16461),
.Y(n_17116)
);

INVx1_ASAP7_75t_L g17117 ( 
.A(n_16463),
.Y(n_17117)
);

INVx1_ASAP7_75t_L g17118 ( 
.A(n_16466),
.Y(n_17118)
);

INVx2_ASAP7_75t_L g17119 ( 
.A(n_16424),
.Y(n_17119)
);

HB1xp67_ASAP7_75t_L g17120 ( 
.A(n_15934),
.Y(n_17120)
);

NOR2x1_ASAP7_75t_L g17121 ( 
.A(n_15875),
.B(n_16038),
.Y(n_17121)
);

INVx2_ASAP7_75t_L g17122 ( 
.A(n_16614),
.Y(n_17122)
);

AND2x2_ASAP7_75t_L g17123 ( 
.A(n_16314),
.B(n_16318),
.Y(n_17123)
);

AND2x4_ASAP7_75t_SL g17124 ( 
.A(n_16553),
.B(n_7831),
.Y(n_17124)
);

INVx1_ASAP7_75t_L g17125 ( 
.A(n_16306),
.Y(n_17125)
);

INVx1_ASAP7_75t_L g17126 ( 
.A(n_16445),
.Y(n_17126)
);

NAND2xp5_ASAP7_75t_L g17127 ( 
.A(n_16088),
.B(n_11022),
.Y(n_17127)
);

AND2x4_ASAP7_75t_L g17128 ( 
.A(n_16593),
.B(n_11022),
.Y(n_17128)
);

NAND2xp5_ASAP7_75t_L g17129 ( 
.A(n_16236),
.B(n_11022),
.Y(n_17129)
);

INVx1_ASAP7_75t_L g17130 ( 
.A(n_16377),
.Y(n_17130)
);

INVx1_ASAP7_75t_L g17131 ( 
.A(n_16360),
.Y(n_17131)
);

INVx1_ASAP7_75t_L g17132 ( 
.A(n_16540),
.Y(n_17132)
);

AND2x4_ASAP7_75t_L g17133 ( 
.A(n_16569),
.B(n_11022),
.Y(n_17133)
);

INVxp67_ASAP7_75t_L g17134 ( 
.A(n_15991),
.Y(n_17134)
);

HB1xp67_ASAP7_75t_L g17135 ( 
.A(n_16030),
.Y(n_17135)
);

NAND2xp5_ASAP7_75t_L g17136 ( 
.A(n_16292),
.B(n_11022),
.Y(n_17136)
);

OR2x2_ASAP7_75t_L g17137 ( 
.A(n_16542),
.B(n_10787),
.Y(n_17137)
);

AND2x2_ASAP7_75t_L g17138 ( 
.A(n_16364),
.B(n_16367),
.Y(n_17138)
);

AND2x2_ASAP7_75t_L g17139 ( 
.A(n_16370),
.B(n_10056),
.Y(n_17139)
);

AND2x2_ASAP7_75t_L g17140 ( 
.A(n_16372),
.B(n_10056),
.Y(n_17140)
);

NAND2xp5_ASAP7_75t_L g17141 ( 
.A(n_16001),
.B(n_11022),
.Y(n_17141)
);

INVx2_ASAP7_75t_SL g17142 ( 
.A(n_16554),
.Y(n_17142)
);

OR2x2_ASAP7_75t_L g17143 ( 
.A(n_16446),
.B(n_11107),
.Y(n_17143)
);

BUFx2_ASAP7_75t_SL g17144 ( 
.A(n_15918),
.Y(n_17144)
);

INVx1_ASAP7_75t_L g17145 ( 
.A(n_16559),
.Y(n_17145)
);

AND2x2_ASAP7_75t_SL g17146 ( 
.A(n_16404),
.B(n_9775),
.Y(n_17146)
);

OR2x6_ASAP7_75t_SL g17147 ( 
.A(n_16257),
.B(n_8962),
.Y(n_17147)
);

AND2x2_ASAP7_75t_L g17148 ( 
.A(n_16047),
.B(n_9974),
.Y(n_17148)
);

AND2x2_ASAP7_75t_L g17149 ( 
.A(n_16340),
.B(n_9974),
.Y(n_17149)
);

INVx2_ASAP7_75t_L g17150 ( 
.A(n_16405),
.Y(n_17150)
);

HB1xp67_ASAP7_75t_L g17151 ( 
.A(n_15947),
.Y(n_17151)
);

NAND2xp5_ASAP7_75t_L g17152 ( 
.A(n_16262),
.B(n_11026),
.Y(n_17152)
);

AND2x2_ASAP7_75t_L g17153 ( 
.A(n_16187),
.B(n_16418),
.Y(n_17153)
);

INVx1_ASAP7_75t_L g17154 ( 
.A(n_16560),
.Y(n_17154)
);

AND2x2_ASAP7_75t_L g17155 ( 
.A(n_16018),
.B(n_9974),
.Y(n_17155)
);

INVx2_ASAP7_75t_L g17156 ( 
.A(n_16090),
.Y(n_17156)
);

CKINVDCx20_ASAP7_75t_R g17157 ( 
.A(n_16546),
.Y(n_17157)
);

INVx2_ASAP7_75t_L g17158 ( 
.A(n_16090),
.Y(n_17158)
);

INVx2_ASAP7_75t_SL g17159 ( 
.A(n_16561),
.Y(n_17159)
);

INVxp67_ASAP7_75t_SL g17160 ( 
.A(n_16044),
.Y(n_17160)
);

INVx1_ASAP7_75t_L g17161 ( 
.A(n_16562),
.Y(n_17161)
);

INVx2_ASAP7_75t_L g17162 ( 
.A(n_16171),
.Y(n_17162)
);

INVx1_ASAP7_75t_L g17163 ( 
.A(n_16563),
.Y(n_17163)
);

HB1xp67_ASAP7_75t_L g17164 ( 
.A(n_15947),
.Y(n_17164)
);

AND2x2_ASAP7_75t_L g17165 ( 
.A(n_16592),
.B(n_9974),
.Y(n_17165)
);

AND2x2_ASAP7_75t_L g17166 ( 
.A(n_16028),
.B(n_9974),
.Y(n_17166)
);

AND2x2_ASAP7_75t_L g17167 ( 
.A(n_16566),
.B(n_9974),
.Y(n_17167)
);

NAND2xp5_ASAP7_75t_L g17168 ( 
.A(n_15940),
.B(n_11026),
.Y(n_17168)
);

AND2x2_ASAP7_75t_L g17169 ( 
.A(n_16454),
.B(n_9974),
.Y(n_17169)
);

AND2x2_ASAP7_75t_L g17170 ( 
.A(n_16302),
.B(n_9974),
.Y(n_17170)
);

INVxp67_ASAP7_75t_L g17171 ( 
.A(n_15977),
.Y(n_17171)
);

AND2x2_ASAP7_75t_L g17172 ( 
.A(n_16305),
.B(n_16578),
.Y(n_17172)
);

OR2x2_ASAP7_75t_L g17173 ( 
.A(n_15911),
.B(n_11107),
.Y(n_17173)
);

INVx1_ASAP7_75t_L g17174 ( 
.A(n_16564),
.Y(n_17174)
);

AND2x2_ASAP7_75t_L g17175 ( 
.A(n_16185),
.B(n_9974),
.Y(n_17175)
);

BUFx3_ASAP7_75t_L g17176 ( 
.A(n_16266),
.Y(n_17176)
);

AND2x4_ASAP7_75t_L g17177 ( 
.A(n_16259),
.B(n_11026),
.Y(n_17177)
);

AND2x2_ASAP7_75t_L g17178 ( 
.A(n_16146),
.B(n_10034),
.Y(n_17178)
);

INVx2_ASAP7_75t_SL g17179 ( 
.A(n_16577),
.Y(n_17179)
);

AND2x2_ASAP7_75t_L g17180 ( 
.A(n_16315),
.B(n_10034),
.Y(n_17180)
);

INVx3_ASAP7_75t_L g17181 ( 
.A(n_16580),
.Y(n_17181)
);

INVx1_ASAP7_75t_L g17182 ( 
.A(n_16581),
.Y(n_17182)
);

AND2x2_ASAP7_75t_L g17183 ( 
.A(n_16336),
.B(n_16198),
.Y(n_17183)
);

NAND2xp5_ASAP7_75t_L g17184 ( 
.A(n_16586),
.B(n_11026),
.Y(n_17184)
);

INVx1_ASAP7_75t_L g17185 ( 
.A(n_16587),
.Y(n_17185)
);

AND2x4_ASAP7_75t_L g17186 ( 
.A(n_16267),
.B(n_11026),
.Y(n_17186)
);

AND2x2_ASAP7_75t_L g17187 ( 
.A(n_16113),
.B(n_16341),
.Y(n_17187)
);

INVx1_ASAP7_75t_L g17188 ( 
.A(n_16591),
.Y(n_17188)
);

INVxp67_ASAP7_75t_SL g17189 ( 
.A(n_16042),
.Y(n_17189)
);

AND2x2_ASAP7_75t_L g17190 ( 
.A(n_16219),
.B(n_10034),
.Y(n_17190)
);

AND2x4_ASAP7_75t_SL g17191 ( 
.A(n_16533),
.B(n_7831),
.Y(n_17191)
);

INVx2_ASAP7_75t_L g17192 ( 
.A(n_16536),
.Y(n_17192)
);

AND2x2_ASAP7_75t_L g17193 ( 
.A(n_16595),
.B(n_10034),
.Y(n_17193)
);

INVx2_ASAP7_75t_L g17194 ( 
.A(n_15913),
.Y(n_17194)
);

NAND2xp5_ASAP7_75t_L g17195 ( 
.A(n_16597),
.B(n_11026),
.Y(n_17195)
);

NOR2xp33_ASAP7_75t_L g17196 ( 
.A(n_15907),
.B(n_10137),
.Y(n_17196)
);

AND2x2_ASAP7_75t_L g17197 ( 
.A(n_16362),
.B(n_10034),
.Y(n_17197)
);

HB1xp67_ASAP7_75t_L g17198 ( 
.A(n_15913),
.Y(n_17198)
);

INVx1_ASAP7_75t_L g17199 ( 
.A(n_16286),
.Y(n_17199)
);

NAND2xp5_ASAP7_75t_L g17200 ( 
.A(n_16190),
.B(n_11026),
.Y(n_17200)
);

INVx2_ASAP7_75t_L g17201 ( 
.A(n_16180),
.Y(n_17201)
);

AND2x4_ASAP7_75t_L g17202 ( 
.A(n_16270),
.B(n_11026),
.Y(n_17202)
);

INVx1_ASAP7_75t_L g17203 ( 
.A(n_16276),
.Y(n_17203)
);

INVx1_ASAP7_75t_L g17204 ( 
.A(n_16134),
.Y(n_17204)
);

BUFx2_ASAP7_75t_L g17205 ( 
.A(n_16369),
.Y(n_17205)
);

OR2x2_ASAP7_75t_L g17206 ( 
.A(n_16151),
.B(n_11107),
.Y(n_17206)
);

AND2x2_ASAP7_75t_L g17207 ( 
.A(n_16387),
.B(n_16338),
.Y(n_17207)
);

INVx1_ASAP7_75t_L g17208 ( 
.A(n_15943),
.Y(n_17208)
);

INVx2_ASAP7_75t_L g17209 ( 
.A(n_16329),
.Y(n_17209)
);

NAND2xp5_ASAP7_75t_L g17210 ( 
.A(n_16400),
.B(n_10754),
.Y(n_17210)
);

OR2x2_ASAP7_75t_L g17211 ( 
.A(n_16607),
.B(n_11107),
.Y(n_17211)
);

AND2x2_ASAP7_75t_L g17212 ( 
.A(n_16061),
.B(n_10034),
.Y(n_17212)
);

AND2x2_ASAP7_75t_L g17213 ( 
.A(n_16064),
.B(n_10034),
.Y(n_17213)
);

AND2x2_ASAP7_75t_L g17214 ( 
.A(n_16517),
.B(n_10034),
.Y(n_17214)
);

AND2x2_ASAP7_75t_L g17215 ( 
.A(n_16080),
.B(n_10034),
.Y(n_17215)
);

INVx1_ASAP7_75t_L g17216 ( 
.A(n_16459),
.Y(n_17216)
);

HB1xp67_ASAP7_75t_L g17217 ( 
.A(n_16608),
.Y(n_17217)
);

HB1xp67_ASAP7_75t_L g17218 ( 
.A(n_16251),
.Y(n_17218)
);

INVx3_ASAP7_75t_L g17219 ( 
.A(n_16084),
.Y(n_17219)
);

NAND2xp5_ASAP7_75t_L g17220 ( 
.A(n_16019),
.B(n_10754),
.Y(n_17220)
);

OR2x2_ASAP7_75t_L g17221 ( 
.A(n_16534),
.B(n_11107),
.Y(n_17221)
);

AND2x2_ASAP7_75t_L g17222 ( 
.A(n_16551),
.B(n_10059),
.Y(n_17222)
);

AND2x2_ASAP7_75t_L g17223 ( 
.A(n_16552),
.B(n_10059),
.Y(n_17223)
);

OR2x2_ASAP7_75t_L g17224 ( 
.A(n_16254),
.B(n_11107),
.Y(n_17224)
);

BUFx3_ASAP7_75t_L g17225 ( 
.A(n_16334),
.Y(n_17225)
);

AND2x2_ASAP7_75t_L g17226 ( 
.A(n_16492),
.B(n_10059),
.Y(n_17226)
);

AND2x2_ASAP7_75t_L g17227 ( 
.A(n_16086),
.B(n_10059),
.Y(n_17227)
);

AND2x2_ASAP7_75t_L g17228 ( 
.A(n_16303),
.B(n_10059),
.Y(n_17228)
);

AND2x2_ASAP7_75t_L g17229 ( 
.A(n_16409),
.B(n_10059),
.Y(n_17229)
);

INVx1_ASAP7_75t_L g17230 ( 
.A(n_16460),
.Y(n_17230)
);

OR2x2_ASAP7_75t_L g17231 ( 
.A(n_15980),
.B(n_11107),
.Y(n_17231)
);

OR2x2_ASAP7_75t_L g17232 ( 
.A(n_16444),
.B(n_11107),
.Y(n_17232)
);

HB1xp67_ASAP7_75t_L g17233 ( 
.A(n_16389),
.Y(n_17233)
);

INVx2_ASAP7_75t_L g17234 ( 
.A(n_16477),
.Y(n_17234)
);

NOR2xp33_ASAP7_75t_L g17235 ( 
.A(n_15944),
.B(n_10137),
.Y(n_17235)
);

INVx1_ASAP7_75t_L g17236 ( 
.A(n_16335),
.Y(n_17236)
);

OR2x2_ASAP7_75t_L g17237 ( 
.A(n_16167),
.B(n_16155),
.Y(n_17237)
);

INVx1_ASAP7_75t_L g17238 ( 
.A(n_16339),
.Y(n_17238)
);

NAND2xp5_ASAP7_75t_SL g17239 ( 
.A(n_16287),
.B(n_10154),
.Y(n_17239)
);

INVx4_ASAP7_75t_L g17240 ( 
.A(n_16415),
.Y(n_17240)
);

OR2x2_ASAP7_75t_L g17241 ( 
.A(n_16210),
.B(n_11202),
.Y(n_17241)
);

INVx1_ASAP7_75t_L g17242 ( 
.A(n_16515),
.Y(n_17242)
);

AND2x2_ASAP7_75t_L g17243 ( 
.A(n_16225),
.B(n_10059),
.Y(n_17243)
);

NAND2x1_ASAP7_75t_SL g17244 ( 
.A(n_16589),
.B(n_10154),
.Y(n_17244)
);

HB1xp67_ASAP7_75t_L g17245 ( 
.A(n_16397),
.Y(n_17245)
);

INVxp67_ASAP7_75t_L g17246 ( 
.A(n_15904),
.Y(n_17246)
);

AND2x2_ASAP7_75t_L g17247 ( 
.A(n_16423),
.B(n_10059),
.Y(n_17247)
);

NAND2xp5_ASAP7_75t_L g17248 ( 
.A(n_16455),
.B(n_10754),
.Y(n_17248)
);

INVx2_ASAP7_75t_SL g17249 ( 
.A(n_16159),
.Y(n_17249)
);

AND2x4_ASAP7_75t_SL g17250 ( 
.A(n_16165),
.B(n_8124),
.Y(n_17250)
);

INVx1_ASAP7_75t_L g17251 ( 
.A(n_16308),
.Y(n_17251)
);

INVx1_ASAP7_75t_SL g17252 ( 
.A(n_16297),
.Y(n_17252)
);

INVx2_ASAP7_75t_L g17253 ( 
.A(n_16361),
.Y(n_17253)
);

INVx2_ASAP7_75t_L g17254 ( 
.A(n_16395),
.Y(n_17254)
);

INVx1_ASAP7_75t_L g17255 ( 
.A(n_16478),
.Y(n_17255)
);

AND2x2_ASAP7_75t_L g17256 ( 
.A(n_16211),
.B(n_10059),
.Y(n_17256)
);

CKINVDCx20_ASAP7_75t_R g17257 ( 
.A(n_16072),
.Y(n_17257)
);

INVx2_ASAP7_75t_L g17258 ( 
.A(n_16342),
.Y(n_17258)
);

INVx1_ASAP7_75t_L g17259 ( 
.A(n_16464),
.Y(n_17259)
);

INVx1_ASAP7_75t_L g17260 ( 
.A(n_16469),
.Y(n_17260)
);

AND2x2_ASAP7_75t_L g17261 ( 
.A(n_16441),
.B(n_10632),
.Y(n_17261)
);

INVx2_ASAP7_75t_SL g17262 ( 
.A(n_16321),
.Y(n_17262)
);

AND2x2_ASAP7_75t_L g17263 ( 
.A(n_16508),
.B(n_10632),
.Y(n_17263)
);

HB1xp67_ASAP7_75t_L g17264 ( 
.A(n_16273),
.Y(n_17264)
);

INVx1_ASAP7_75t_L g17265 ( 
.A(n_16476),
.Y(n_17265)
);

INVxp67_ASAP7_75t_L g17266 ( 
.A(n_15982),
.Y(n_17266)
);

NAND4xp25_ASAP7_75t_L g17267 ( 
.A(n_16221),
.B(n_9472),
.C(n_9526),
.D(n_9461),
.Y(n_17267)
);

HB1xp67_ASAP7_75t_L g17268 ( 
.A(n_16282),
.Y(n_17268)
);

AND2x2_ASAP7_75t_SL g17269 ( 
.A(n_16106),
.B(n_16049),
.Y(n_17269)
);

INVx1_ASAP7_75t_L g17270 ( 
.A(n_16491),
.Y(n_17270)
);

INVxp67_ASAP7_75t_L g17271 ( 
.A(n_16289),
.Y(n_17271)
);

INVx1_ASAP7_75t_L g17272 ( 
.A(n_16511),
.Y(n_17272)
);

AND2x2_ASAP7_75t_L g17273 ( 
.A(n_16137),
.B(n_10632),
.Y(n_17273)
);

NAND2xp5_ASAP7_75t_L g17274 ( 
.A(n_16035),
.B(n_10754),
.Y(n_17274)
);

AND2x2_ASAP7_75t_L g17275 ( 
.A(n_16385),
.B(n_10632),
.Y(n_17275)
);

OR2x2_ASAP7_75t_L g17276 ( 
.A(n_16233),
.B(n_11202),
.Y(n_17276)
);

INVx2_ASAP7_75t_L g17277 ( 
.A(n_16345),
.Y(n_17277)
);

INVx2_ASAP7_75t_L g17278 ( 
.A(n_16475),
.Y(n_17278)
);

AND2x2_ASAP7_75t_L g17279 ( 
.A(n_16130),
.B(n_10632),
.Y(n_17279)
);

AND2x2_ASAP7_75t_L g17280 ( 
.A(n_16497),
.B(n_10632),
.Y(n_17280)
);

INVx1_ASAP7_75t_L g17281 ( 
.A(n_16296),
.Y(n_17281)
);

INVx2_ASAP7_75t_L g17282 ( 
.A(n_16120),
.Y(n_17282)
);

AND2x2_ASAP7_75t_L g17283 ( 
.A(n_16429),
.B(n_10632),
.Y(n_17283)
);

AND2x2_ASAP7_75t_L g17284 ( 
.A(n_16584),
.B(n_16258),
.Y(n_17284)
);

INVx4_ASAP7_75t_L g17285 ( 
.A(n_16093),
.Y(n_17285)
);

HB1xp67_ASAP7_75t_L g17286 ( 
.A(n_16348),
.Y(n_17286)
);

OR2x2_ASAP7_75t_L g17287 ( 
.A(n_16337),
.B(n_11202),
.Y(n_17287)
);

INVx1_ASAP7_75t_SL g17288 ( 
.A(n_16346),
.Y(n_17288)
);

AND2x4_ASAP7_75t_L g17289 ( 
.A(n_16186),
.B(n_10669),
.Y(n_17289)
);

INVx1_ASAP7_75t_L g17290 ( 
.A(n_16365),
.Y(n_17290)
);

INVx1_ASAP7_75t_L g17291 ( 
.A(n_16411),
.Y(n_17291)
);

NOR2x1p5_ASAP7_75t_L g17292 ( 
.A(n_16857),
.B(n_16101),
.Y(n_17292)
);

AND2x2_ASAP7_75t_L g17293 ( 
.A(n_16640),
.B(n_16621),
.Y(n_17293)
);

INVx1_ASAP7_75t_L g17294 ( 
.A(n_16660),
.Y(n_17294)
);

INVx1_ASAP7_75t_L g17295 ( 
.A(n_16660),
.Y(n_17295)
);

INVx1_ASAP7_75t_L g17296 ( 
.A(n_16670),
.Y(n_17296)
);

AND2x2_ASAP7_75t_L g17297 ( 
.A(n_16632),
.B(n_16363),
.Y(n_17297)
);

INVx3_ASAP7_75t_L g17298 ( 
.A(n_16652),
.Y(n_17298)
);

OAI21x1_ASAP7_75t_L g17299 ( 
.A1(n_17051),
.A2(n_16568),
.B(n_16140),
.Y(n_17299)
);

BUFx2_ASAP7_75t_L g17300 ( 
.A(n_16700),
.Y(n_17300)
);

OR2x2_ASAP7_75t_L g17301 ( 
.A(n_16704),
.B(n_16715),
.Y(n_17301)
);

INVx1_ASAP7_75t_L g17302 ( 
.A(n_16684),
.Y(n_17302)
);

INVx1_ASAP7_75t_L g17303 ( 
.A(n_16626),
.Y(n_17303)
);

OAI21x1_ASAP7_75t_L g17304 ( 
.A1(n_16885),
.A2(n_16232),
.B(n_16110),
.Y(n_17304)
);

INVx1_ASAP7_75t_L g17305 ( 
.A(n_16649),
.Y(n_17305)
);

INVx1_ASAP7_75t_L g17306 ( 
.A(n_16669),
.Y(n_17306)
);

INVx1_ASAP7_75t_L g17307 ( 
.A(n_16686),
.Y(n_17307)
);

OR2x6_ASAP7_75t_L g17308 ( 
.A(n_16734),
.B(n_9756),
.Y(n_17308)
);

INVx2_ASAP7_75t_L g17309 ( 
.A(n_16879),
.Y(n_17309)
);

INVx2_ASAP7_75t_L g17310 ( 
.A(n_16879),
.Y(n_17310)
);

AND2x4_ASAP7_75t_L g17311 ( 
.A(n_16736),
.B(n_10669),
.Y(n_17311)
);

OR2x6_ASAP7_75t_L g17312 ( 
.A(n_16624),
.B(n_9756),
.Y(n_17312)
);

AND2x2_ASAP7_75t_L g17313 ( 
.A(n_16703),
.B(n_16616),
.Y(n_17313)
);

OR2x6_ASAP7_75t_L g17314 ( 
.A(n_16636),
.B(n_9756),
.Y(n_17314)
);

NAND2xp5_ASAP7_75t_L g17315 ( 
.A(n_16714),
.B(n_16206),
.Y(n_17315)
);

OA21x2_ASAP7_75t_L g17316 ( 
.A1(n_16637),
.A2(n_16129),
.B(n_16558),
.Y(n_17316)
);

OAI21xp5_ASAP7_75t_L g17317 ( 
.A1(n_16827),
.A2(n_16098),
.B(n_16118),
.Y(n_17317)
);

INVx1_ASAP7_75t_L g17318 ( 
.A(n_16657),
.Y(n_17318)
);

INVx2_ASAP7_75t_L g17319 ( 
.A(n_16688),
.Y(n_17319)
);

INVx1_ASAP7_75t_L g17320 ( 
.A(n_16659),
.Y(n_17320)
);

BUFx2_ASAP7_75t_L g17321 ( 
.A(n_16709),
.Y(n_17321)
);

BUFx3_ASAP7_75t_L g17322 ( 
.A(n_16674),
.Y(n_17322)
);

INVx1_ASAP7_75t_L g17323 ( 
.A(n_16688),
.Y(n_17323)
);

OAI21xp5_ASAP7_75t_SL g17324 ( 
.A1(n_16998),
.A2(n_16122),
.B(n_16143),
.Y(n_17324)
);

OR2x6_ASAP7_75t_L g17325 ( 
.A(n_16797),
.B(n_9756),
.Y(n_17325)
);

NAND2xp5_ASAP7_75t_SL g17326 ( 
.A(n_16998),
.B(n_16615),
.Y(n_17326)
);

AND2x6_ASAP7_75t_SL g17327 ( 
.A(n_16749),
.B(n_9333),
.Y(n_17327)
);

AND2x2_ASAP7_75t_L g17328 ( 
.A(n_16645),
.B(n_16207),
.Y(n_17328)
);

INVx1_ASAP7_75t_L g17329 ( 
.A(n_16691),
.Y(n_17329)
);

OR2x2_ASAP7_75t_L g17330 ( 
.A(n_16710),
.B(n_16319),
.Y(n_17330)
);

HB1xp67_ASAP7_75t_L g17331 ( 
.A(n_16620),
.Y(n_17331)
);

INVx1_ASAP7_75t_L g17332 ( 
.A(n_16825),
.Y(n_17332)
);

HB1xp67_ASAP7_75t_L g17333 ( 
.A(n_16682),
.Y(n_17333)
);

NOR2x1_ASAP7_75t_SL g17334 ( 
.A(n_16761),
.B(n_16826),
.Y(n_17334)
);

NAND3xp33_ASAP7_75t_L g17335 ( 
.A(n_17102),
.B(n_16041),
.C(n_16058),
.Y(n_17335)
);

INVx1_ASAP7_75t_L g17336 ( 
.A(n_16685),
.Y(n_17336)
);

INVx1_ASAP7_75t_L g17337 ( 
.A(n_16685),
.Y(n_17337)
);

BUFx3_ASAP7_75t_L g17338 ( 
.A(n_16656),
.Y(n_17338)
);

OA21x2_ASAP7_75t_L g17339 ( 
.A1(n_16884),
.A2(n_16575),
.B(n_16085),
.Y(n_17339)
);

NAND2xp5_ASAP7_75t_SL g17340 ( 
.A(n_16976),
.B(n_16545),
.Y(n_17340)
);

OAI21x1_ASAP7_75t_L g17341 ( 
.A1(n_17056),
.A2(n_16982),
.B(n_16683),
.Y(n_17341)
);

INVx1_ASAP7_75t_L g17342 ( 
.A(n_16810),
.Y(n_17342)
);

NAND2xp5_ASAP7_75t_L g17343 ( 
.A(n_16628),
.B(n_16214),
.Y(n_17343)
);

NAND3xp33_ASAP7_75t_SL g17344 ( 
.A(n_16976),
.B(n_16931),
.C(n_17037),
.Y(n_17344)
);

NOR3xp33_ASAP7_75t_SL g17345 ( 
.A(n_16779),
.B(n_16224),
.C(n_16116),
.Y(n_17345)
);

INVx2_ASAP7_75t_L g17346 ( 
.A(n_16629),
.Y(n_17346)
);

NAND2xp5_ASAP7_75t_L g17347 ( 
.A(n_16633),
.B(n_16226),
.Y(n_17347)
);

INVx1_ASAP7_75t_L g17348 ( 
.A(n_16811),
.Y(n_17348)
);

AOI21x1_ASAP7_75t_L g17349 ( 
.A1(n_16884),
.A2(n_16059),
.B(n_16582),
.Y(n_17349)
);

INVx1_ASAP7_75t_L g17350 ( 
.A(n_16814),
.Y(n_17350)
);

HB1xp67_ASAP7_75t_L g17351 ( 
.A(n_16787),
.Y(n_17351)
);

HB1xp67_ASAP7_75t_L g17352 ( 
.A(n_16886),
.Y(n_17352)
);

OA21x2_ASAP7_75t_L g17353 ( 
.A1(n_16886),
.A2(n_16590),
.B(n_16427),
.Y(n_17353)
);

INVx1_ASAP7_75t_L g17354 ( 
.A(n_16881),
.Y(n_17354)
);

INVx1_ASAP7_75t_L g17355 ( 
.A(n_16888),
.Y(n_17355)
);

OA21x2_ASAP7_75t_L g17356 ( 
.A1(n_16777),
.A2(n_16832),
.B(n_16829),
.Y(n_17356)
);

INVx2_ASAP7_75t_L g17357 ( 
.A(n_16623),
.Y(n_17357)
);

BUFx3_ASAP7_75t_L g17358 ( 
.A(n_16643),
.Y(n_17358)
);

OA21x2_ASAP7_75t_L g17359 ( 
.A1(n_16833),
.A2(n_16631),
.B(n_16931),
.Y(n_17359)
);

NAND2xp5_ASAP7_75t_SL g17360 ( 
.A(n_17194),
.B(n_16719),
.Y(n_17360)
);

NAND3xp33_ASAP7_75t_L g17361 ( 
.A(n_17120),
.B(n_16094),
.C(n_16539),
.Y(n_17361)
);

INVx2_ASAP7_75t_L g17362 ( 
.A(n_16639),
.Y(n_17362)
);

OA21x2_ASAP7_75t_L g17363 ( 
.A1(n_16804),
.A2(n_16830),
.B(n_16822),
.Y(n_17363)
);

HB1xp67_ASAP7_75t_L g17364 ( 
.A(n_16625),
.Y(n_17364)
);

INVx1_ASAP7_75t_L g17365 ( 
.A(n_16798),
.Y(n_17365)
);

INVx2_ASAP7_75t_L g17366 ( 
.A(n_16651),
.Y(n_17366)
);

INVxp67_ASAP7_75t_L g17367 ( 
.A(n_16987),
.Y(n_17367)
);

INVx4_ASAP7_75t_L g17368 ( 
.A(n_16693),
.Y(n_17368)
);

INVx1_ASAP7_75t_L g17369 ( 
.A(n_16842),
.Y(n_17369)
);

INVx1_ASAP7_75t_L g17370 ( 
.A(n_16845),
.Y(n_17370)
);

INVxp67_ASAP7_75t_SL g17371 ( 
.A(n_16799),
.Y(n_17371)
);

INVx1_ASAP7_75t_L g17372 ( 
.A(n_16846),
.Y(n_17372)
);

OA21x2_ASAP7_75t_L g17373 ( 
.A1(n_16794),
.A2(n_16432),
.B(n_16422),
.Y(n_17373)
);

OA21x2_ASAP7_75t_L g17374 ( 
.A1(n_17205),
.A2(n_16557),
.B(n_16548),
.Y(n_17374)
);

INVx1_ASAP7_75t_L g17375 ( 
.A(n_16667),
.Y(n_17375)
);

INVx1_ASAP7_75t_L g17376 ( 
.A(n_16789),
.Y(n_17376)
);

INVx1_ASAP7_75t_L g17377 ( 
.A(n_16792),
.Y(n_17377)
);

OR2x2_ASAP7_75t_L g17378 ( 
.A(n_16647),
.B(n_16191),
.Y(n_17378)
);

INVx2_ASAP7_75t_L g17379 ( 
.A(n_16668),
.Y(n_17379)
);

BUFx3_ASAP7_75t_L g17380 ( 
.A(n_16747),
.Y(n_17380)
);

INVx2_ASAP7_75t_L g17381 ( 
.A(n_16642),
.Y(n_17381)
);

INVx2_ASAP7_75t_L g17382 ( 
.A(n_16638),
.Y(n_17382)
);

INVx2_ASAP7_75t_L g17383 ( 
.A(n_16672),
.Y(n_17383)
);

AND2x2_ASAP7_75t_L g17384 ( 
.A(n_16676),
.B(n_16537),
.Y(n_17384)
);

BUFx2_ASAP7_75t_L g17385 ( 
.A(n_17113),
.Y(n_17385)
);

INVx2_ASAP7_75t_L g17386 ( 
.A(n_16743),
.Y(n_17386)
);

NAND3xp33_ASAP7_75t_L g17387 ( 
.A(n_16947),
.B(n_16205),
.C(n_16602),
.Y(n_17387)
);

OA21x2_ASAP7_75t_L g17388 ( 
.A1(n_17205),
.A2(n_16222),
.B(n_16218),
.Y(n_17388)
);

OA21x2_ASAP7_75t_L g17389 ( 
.A1(n_16890),
.A2(n_16223),
.B(n_16603),
.Y(n_17389)
);

INVx3_ASAP7_75t_L g17390 ( 
.A(n_17025),
.Y(n_17390)
);

AOI21xp5_ASAP7_75t_L g17391 ( 
.A1(n_16864),
.A2(n_16977),
.B(n_17121),
.Y(n_17391)
);

INVx1_ASAP7_75t_L g17392 ( 
.A(n_16783),
.Y(n_17392)
);

BUFx3_ASAP7_75t_L g17393 ( 
.A(n_16664),
.Y(n_17393)
);

OR2x2_ASAP7_75t_L g17394 ( 
.A(n_16646),
.B(n_16450),
.Y(n_17394)
);

BUFx2_ASAP7_75t_L g17395 ( 
.A(n_16737),
.Y(n_17395)
);

BUFx2_ASAP7_75t_L g17396 ( 
.A(n_16677),
.Y(n_17396)
);

OA21x2_ASAP7_75t_L g17397 ( 
.A1(n_16892),
.A2(n_16609),
.B(n_16606),
.Y(n_17397)
);

INVx2_ASAP7_75t_L g17398 ( 
.A(n_16713),
.Y(n_17398)
);

INVx1_ASAP7_75t_SL g17399 ( 
.A(n_16896),
.Y(n_17399)
);

NAND2xp5_ASAP7_75t_SL g17400 ( 
.A(n_17198),
.B(n_16612),
.Y(n_17400)
);

OA21x2_ASAP7_75t_L g17401 ( 
.A1(n_16813),
.A2(n_16610),
.B(n_16081),
.Y(n_17401)
);

INVx1_ASAP7_75t_L g17402 ( 
.A(n_16641),
.Y(n_17402)
);

OR2x6_ASAP7_75t_L g17403 ( 
.A(n_16702),
.B(n_10027),
.Y(n_17403)
);

BUFx2_ASAP7_75t_L g17404 ( 
.A(n_16728),
.Y(n_17404)
);

INVx2_ASAP7_75t_L g17405 ( 
.A(n_16716),
.Y(n_17405)
);

INVx4_ASAP7_75t_SL g17406 ( 
.A(n_16634),
.Y(n_17406)
);

OR2x6_ASAP7_75t_L g17407 ( 
.A(n_16698),
.B(n_16753),
.Y(n_17407)
);

INVx2_ASAP7_75t_L g17408 ( 
.A(n_16732),
.Y(n_17408)
);

HB1xp67_ASAP7_75t_L g17409 ( 
.A(n_16627),
.Y(n_17409)
);

OR2x2_ASAP7_75t_L g17410 ( 
.A(n_16724),
.B(n_16507),
.Y(n_17410)
);

INVx1_ASAP7_75t_L g17411 ( 
.A(n_16785),
.Y(n_17411)
);

OR2x2_ASAP7_75t_L g17412 ( 
.A(n_16731),
.B(n_16528),
.Y(n_17412)
);

NAND2xp5_ASAP7_75t_L g17413 ( 
.A(n_16745),
.B(n_16242),
.Y(n_17413)
);

INVx1_ASAP7_75t_L g17414 ( 
.A(n_16654),
.Y(n_17414)
);

OAI21x1_ASAP7_75t_L g17415 ( 
.A1(n_16673),
.A2(n_16472),
.B(n_11677),
.Y(n_17415)
);

NAND2xp5_ASAP7_75t_L g17416 ( 
.A(n_16768),
.B(n_10985),
.Y(n_17416)
);

INVx1_ASAP7_75t_L g17417 ( 
.A(n_16658),
.Y(n_17417)
);

INVx2_ASAP7_75t_L g17418 ( 
.A(n_16739),
.Y(n_17418)
);

INVx1_ASAP7_75t_L g17419 ( 
.A(n_16662),
.Y(n_17419)
);

INVx1_ASAP7_75t_L g17420 ( 
.A(n_16666),
.Y(n_17420)
);

INVx3_ASAP7_75t_L g17421 ( 
.A(n_16893),
.Y(n_17421)
);

INVx1_ASAP7_75t_L g17422 ( 
.A(n_16648),
.Y(n_17422)
);

AND2x2_ASAP7_75t_L g17423 ( 
.A(n_16681),
.B(n_10669),
.Y(n_17423)
);

INVx4_ASAP7_75t_SL g17424 ( 
.A(n_16692),
.Y(n_17424)
);

AND2x2_ASAP7_75t_L g17425 ( 
.A(n_16706),
.B(n_10669),
.Y(n_17425)
);

INVx2_ASAP7_75t_L g17426 ( 
.A(n_16675),
.Y(n_17426)
);

INVx1_ASAP7_75t_L g17427 ( 
.A(n_16705),
.Y(n_17427)
);

BUFx2_ASAP7_75t_L g17428 ( 
.A(n_16980),
.Y(n_17428)
);

HB1xp67_ASAP7_75t_L g17429 ( 
.A(n_16807),
.Y(n_17429)
);

BUFx2_ASAP7_75t_L g17430 ( 
.A(n_17097),
.Y(n_17430)
);

BUFx6f_ASAP7_75t_L g17431 ( 
.A(n_16687),
.Y(n_17431)
);

INVx2_ASAP7_75t_SL g17432 ( 
.A(n_16895),
.Y(n_17432)
);

AND2x2_ASAP7_75t_L g17433 ( 
.A(n_16755),
.B(n_10669),
.Y(n_17433)
);

INVx4_ASAP7_75t_SL g17434 ( 
.A(n_16989),
.Y(n_17434)
);

INVx1_ASAP7_75t_L g17435 ( 
.A(n_16725),
.Y(n_17435)
);

INVx1_ASAP7_75t_SL g17436 ( 
.A(n_16767),
.Y(n_17436)
);

INVx1_ASAP7_75t_L g17437 ( 
.A(n_16974),
.Y(n_17437)
);

INVx2_ASAP7_75t_L g17438 ( 
.A(n_16754),
.Y(n_17438)
);

INVx2_ASAP7_75t_L g17439 ( 
.A(n_16707),
.Y(n_17439)
);

AND2x2_ASAP7_75t_L g17440 ( 
.A(n_16831),
.B(n_10669),
.Y(n_17440)
);

OR2x2_ASAP7_75t_L g17441 ( 
.A(n_16712),
.B(n_16571),
.Y(n_17441)
);

INVx1_ASAP7_75t_L g17442 ( 
.A(n_16788),
.Y(n_17442)
);

INVx1_ASAP7_75t_L g17443 ( 
.A(n_16733),
.Y(n_17443)
);

BUFx2_ASAP7_75t_L g17444 ( 
.A(n_16817),
.Y(n_17444)
);

AOI21xp5_ASAP7_75t_L g17445 ( 
.A1(n_16781),
.A2(n_13640),
.B(n_13594),
.Y(n_17445)
);

INVx1_ASAP7_75t_L g17446 ( 
.A(n_16711),
.Y(n_17446)
);

INVx1_ASAP7_75t_SL g17447 ( 
.A(n_16803),
.Y(n_17447)
);

OR2x2_ASAP7_75t_L g17448 ( 
.A(n_16635),
.B(n_11202),
.Y(n_17448)
);

INVx1_ASAP7_75t_L g17449 ( 
.A(n_16622),
.Y(n_17449)
);

BUFx8_ASAP7_75t_L g17450 ( 
.A(n_16671),
.Y(n_17450)
);

INVx1_ASAP7_75t_L g17451 ( 
.A(n_16630),
.Y(n_17451)
);

INVx2_ASAP7_75t_L g17452 ( 
.A(n_16720),
.Y(n_17452)
);

INVx1_ASAP7_75t_L g17453 ( 
.A(n_16738),
.Y(n_17453)
);

INVx4_ASAP7_75t_SL g17454 ( 
.A(n_16694),
.Y(n_17454)
);

HB1xp67_ASAP7_75t_L g17455 ( 
.A(n_16808),
.Y(n_17455)
);

INVx2_ASAP7_75t_L g17456 ( 
.A(n_16882),
.Y(n_17456)
);

OA21x2_ASAP7_75t_L g17457 ( 
.A1(n_17290),
.A2(n_10930),
.B(n_10913),
.Y(n_17457)
);

INVx1_ASAP7_75t_SL g17458 ( 
.A(n_16663),
.Y(n_17458)
);

INVx2_ASAP7_75t_L g17459 ( 
.A(n_16723),
.Y(n_17459)
);

INVx2_ASAP7_75t_L g17460 ( 
.A(n_16678),
.Y(n_17460)
);

NAND3xp33_ASAP7_75t_SL g17461 ( 
.A(n_17257),
.B(n_10038),
.C(n_10011),
.Y(n_17461)
);

OA21x2_ASAP7_75t_L g17462 ( 
.A1(n_17189),
.A2(n_17251),
.B(n_17238),
.Y(n_17462)
);

INVx1_ASAP7_75t_L g17463 ( 
.A(n_16746),
.Y(n_17463)
);

INVx4_ASAP7_75t_SL g17464 ( 
.A(n_16695),
.Y(n_17464)
);

NAND2xp5_ASAP7_75t_L g17465 ( 
.A(n_16839),
.B(n_10985),
.Y(n_17465)
);

INVx2_ASAP7_75t_L g17466 ( 
.A(n_16771),
.Y(n_17466)
);

OA21x2_ASAP7_75t_L g17467 ( 
.A1(n_17236),
.A2(n_10932),
.B(n_10930),
.Y(n_17467)
);

AND2x2_ASAP7_75t_L g17468 ( 
.A(n_16759),
.B(n_10669),
.Y(n_17468)
);

BUFx2_ASAP7_75t_L g17469 ( 
.A(n_16954),
.Y(n_17469)
);

INVx1_ASAP7_75t_L g17470 ( 
.A(n_16708),
.Y(n_17470)
);

INVx1_ASAP7_75t_L g17471 ( 
.A(n_16741),
.Y(n_17471)
);

INVx1_ASAP7_75t_L g17472 ( 
.A(n_16679),
.Y(n_17472)
);

INVxp67_ASAP7_75t_SL g17473 ( 
.A(n_17151),
.Y(n_17473)
);

BUFx2_ASAP7_75t_L g17474 ( 
.A(n_16930),
.Y(n_17474)
);

INVx4_ASAP7_75t_SL g17475 ( 
.A(n_16752),
.Y(n_17475)
);

INVx4_ASAP7_75t_SL g17476 ( 
.A(n_16852),
.Y(n_17476)
);

INVx1_ASAP7_75t_L g17477 ( 
.A(n_16911),
.Y(n_17477)
);

INVx1_ASAP7_75t_L g17478 ( 
.A(n_16914),
.Y(n_17478)
);

INVx2_ASAP7_75t_L g17479 ( 
.A(n_17114),
.Y(n_17479)
);

INVxp67_ASAP7_75t_L g17480 ( 
.A(n_17164),
.Y(n_17480)
);

INVx1_ASAP7_75t_L g17481 ( 
.A(n_16916),
.Y(n_17481)
);

AOI21xp5_ASAP7_75t_L g17482 ( 
.A1(n_16760),
.A2(n_13640),
.B(n_13594),
.Y(n_17482)
);

INVx4_ASAP7_75t_SL g17483 ( 
.A(n_16802),
.Y(n_17483)
);

INVx2_ASAP7_75t_L g17484 ( 
.A(n_17114),
.Y(n_17484)
);

AND2x4_ASAP7_75t_L g17485 ( 
.A(n_16727),
.B(n_10898),
.Y(n_17485)
);

INVx1_ASAP7_75t_L g17486 ( 
.A(n_16919),
.Y(n_17486)
);

INVx3_ASAP7_75t_L g17487 ( 
.A(n_16901),
.Y(n_17487)
);

INVx2_ASAP7_75t_L g17488 ( 
.A(n_16763),
.Y(n_17488)
);

HB1xp67_ASAP7_75t_L g17489 ( 
.A(n_17069),
.Y(n_17489)
);

OAI21x1_ASAP7_75t_L g17490 ( 
.A1(n_16690),
.A2(n_12238),
.B(n_12657),
.Y(n_17490)
);

INVx1_ASAP7_75t_SL g17491 ( 
.A(n_16740),
.Y(n_17491)
);

INVx1_ASAP7_75t_SL g17492 ( 
.A(n_16942),
.Y(n_17492)
);

INVx2_ASAP7_75t_L g17493 ( 
.A(n_16801),
.Y(n_17493)
);

INVx1_ASAP7_75t_L g17494 ( 
.A(n_16848),
.Y(n_17494)
);

INVx1_ASAP7_75t_L g17495 ( 
.A(n_16859),
.Y(n_17495)
);

INVx2_ASAP7_75t_L g17496 ( 
.A(n_16838),
.Y(n_17496)
);

HB1xp67_ASAP7_75t_L g17497 ( 
.A(n_17027),
.Y(n_17497)
);

INVx2_ASAP7_75t_L g17498 ( 
.A(n_16816),
.Y(n_17498)
);

INVx1_ASAP7_75t_L g17499 ( 
.A(n_16820),
.Y(n_17499)
);

INVxp67_ASAP7_75t_SL g17500 ( 
.A(n_17255),
.Y(n_17500)
);

INVx2_ASAP7_75t_L g17501 ( 
.A(n_16904),
.Y(n_17501)
);

BUFx3_ASAP7_75t_L g17502 ( 
.A(n_16699),
.Y(n_17502)
);

INVx1_ASAP7_75t_L g17503 ( 
.A(n_16867),
.Y(n_17503)
);

HB1xp67_ASAP7_75t_L g17504 ( 
.A(n_17040),
.Y(n_17504)
);

HB1xp67_ASAP7_75t_L g17505 ( 
.A(n_17077),
.Y(n_17505)
);

HB1xp67_ASAP7_75t_L g17506 ( 
.A(n_16821),
.Y(n_17506)
);

NAND2xp5_ASAP7_75t_SL g17507 ( 
.A(n_17289),
.B(n_10154),
.Y(n_17507)
);

OA21x2_ASAP7_75t_L g17508 ( 
.A1(n_17160),
.A2(n_10935),
.B(n_10932),
.Y(n_17508)
);

INVx1_ASAP7_75t_L g17509 ( 
.A(n_16796),
.Y(n_17509)
);

INVxp67_ASAP7_75t_L g17510 ( 
.A(n_16775),
.Y(n_17510)
);

INVx1_ASAP7_75t_L g17511 ( 
.A(n_16851),
.Y(n_17511)
);

AND2x2_ASAP7_75t_L g17512 ( 
.A(n_16856),
.B(n_10898),
.Y(n_17512)
);

INVx1_ASAP7_75t_L g17513 ( 
.A(n_16655),
.Y(n_17513)
);

INVx1_ASAP7_75t_L g17514 ( 
.A(n_16665),
.Y(n_17514)
);

INVx1_ASAP7_75t_L g17515 ( 
.A(n_16840),
.Y(n_17515)
);

INVx3_ASAP7_75t_L g17516 ( 
.A(n_16901),
.Y(n_17516)
);

INVx2_ASAP7_75t_L g17517 ( 
.A(n_16756),
.Y(n_17517)
);

AO21x1_ASAP7_75t_L g17518 ( 
.A1(n_16718),
.A2(n_11162),
.B(n_11158),
.Y(n_17518)
);

OAI21x1_ASAP7_75t_L g17519 ( 
.A1(n_16726),
.A2(n_12679),
.B(n_12662),
.Y(n_17519)
);

AOI21xp5_ASAP7_75t_L g17520 ( 
.A1(n_16979),
.A2(n_13653),
.B(n_11837),
.Y(n_17520)
);

INVx2_ASAP7_75t_L g17521 ( 
.A(n_16701),
.Y(n_17521)
);

INVx1_ASAP7_75t_L g17522 ( 
.A(n_16868),
.Y(n_17522)
);

INVx2_ASAP7_75t_L g17523 ( 
.A(n_16806),
.Y(n_17523)
);

OAI21x1_ASAP7_75t_L g17524 ( 
.A1(n_16644),
.A2(n_16680),
.B(n_16653),
.Y(n_17524)
);

INVx1_ASAP7_75t_L g17525 ( 
.A(n_16921),
.Y(n_17525)
);

AND2x2_ASAP7_75t_L g17526 ( 
.A(n_16770),
.B(n_10898),
.Y(n_17526)
);

INVx3_ASAP7_75t_L g17527 ( 
.A(n_16932),
.Y(n_17527)
);

OAI21x1_ASAP7_75t_L g17528 ( 
.A1(n_16786),
.A2(n_12687),
.B(n_12126),
.Y(n_17528)
);

INVx2_ASAP7_75t_L g17529 ( 
.A(n_16936),
.Y(n_17529)
);

INVx2_ASAP7_75t_L g17530 ( 
.A(n_16951),
.Y(n_17530)
);

INVx2_ASAP7_75t_L g17531 ( 
.A(n_16855),
.Y(n_17531)
);

INVx1_ASAP7_75t_L g17532 ( 
.A(n_17020),
.Y(n_17532)
);

INVx4_ASAP7_75t_SL g17533 ( 
.A(n_16815),
.Y(n_17533)
);

HB1xp67_ASAP7_75t_L g17534 ( 
.A(n_17286),
.Y(n_17534)
);

HB1xp67_ASAP7_75t_L g17535 ( 
.A(n_17046),
.Y(n_17535)
);

INVx1_ASAP7_75t_L g17536 ( 
.A(n_17022),
.Y(n_17536)
);

INVx1_ASAP7_75t_L g17537 ( 
.A(n_16926),
.Y(n_17537)
);

INVx5_ASAP7_75t_L g17538 ( 
.A(n_16835),
.Y(n_17538)
);

INVx1_ASAP7_75t_L g17539 ( 
.A(n_16928),
.Y(n_17539)
);

AOI21xp5_ASAP7_75t_L g17540 ( 
.A1(n_16969),
.A2(n_13653),
.B(n_11837),
.Y(n_17540)
);

AND2x2_ASAP7_75t_L g17541 ( 
.A(n_16828),
.B(n_10898),
.Y(n_17541)
);

INVx2_ASAP7_75t_L g17542 ( 
.A(n_17244),
.Y(n_17542)
);

BUFx2_ASAP7_75t_L g17543 ( 
.A(n_16872),
.Y(n_17543)
);

OA21x2_ASAP7_75t_L g17544 ( 
.A1(n_17281),
.A2(n_10937),
.B(n_10935),
.Y(n_17544)
);

AND2x4_ASAP7_75t_L g17545 ( 
.A(n_16650),
.B(n_10898),
.Y(n_17545)
);

INVxp67_ASAP7_75t_SL g17546 ( 
.A(n_16834),
.Y(n_17546)
);

AOI21xp33_ASAP7_75t_L g17547 ( 
.A1(n_17135),
.A2(n_10897),
.B(n_11367),
.Y(n_17547)
);

AND2x2_ASAP7_75t_L g17548 ( 
.A(n_16772),
.B(n_10898),
.Y(n_17548)
);

INVx1_ASAP7_75t_SL g17549 ( 
.A(n_16762),
.Y(n_17549)
);

INVx1_ASAP7_75t_L g17550 ( 
.A(n_16941),
.Y(n_17550)
);

INVx2_ASAP7_75t_L g17551 ( 
.A(n_16765),
.Y(n_17551)
);

AND2x2_ASAP7_75t_L g17552 ( 
.A(n_16780),
.B(n_10898),
.Y(n_17552)
);

NAND3xp33_ASAP7_75t_L g17553 ( 
.A(n_17246),
.B(n_17218),
.C(n_16721),
.Y(n_17553)
);

INVx5_ASAP7_75t_L g17554 ( 
.A(n_16841),
.Y(n_17554)
);

NOR2x1p5_ASAP7_75t_L g17555 ( 
.A(n_16722),
.B(n_9092),
.Y(n_17555)
);

BUFx2_ASAP7_75t_L g17556 ( 
.A(n_16999),
.Y(n_17556)
);

INVx1_ASAP7_75t_L g17557 ( 
.A(n_16948),
.Y(n_17557)
);

INVx1_ASAP7_75t_L g17558 ( 
.A(n_16961),
.Y(n_17558)
);

INVx2_ASAP7_75t_L g17559 ( 
.A(n_17057),
.Y(n_17559)
);

BUFx2_ASAP7_75t_L g17560 ( 
.A(n_17073),
.Y(n_17560)
);

INVx3_ASAP7_75t_L g17561 ( 
.A(n_16932),
.Y(n_17561)
);

INVx1_ASAP7_75t_L g17562 ( 
.A(n_16967),
.Y(n_17562)
);

INVx2_ASAP7_75t_L g17563 ( 
.A(n_17076),
.Y(n_17563)
);

INVx1_ASAP7_75t_SL g17564 ( 
.A(n_17144),
.Y(n_17564)
);

INVx1_ASAP7_75t_L g17565 ( 
.A(n_16850),
.Y(n_17565)
);

OA21x2_ASAP7_75t_L g17566 ( 
.A1(n_16990),
.A2(n_10938),
.B(n_10937),
.Y(n_17566)
);

OA21x2_ASAP7_75t_L g17567 ( 
.A1(n_17271),
.A2(n_10941),
.B(n_10938),
.Y(n_17567)
);

OAI21xp5_ASAP7_75t_L g17568 ( 
.A1(n_17266),
.A2(n_10774),
.B(n_10771),
.Y(n_17568)
);

NAND2xp5_ASAP7_75t_SL g17569 ( 
.A(n_17146),
.B(n_10155),
.Y(n_17569)
);

INVx3_ASAP7_75t_L g17570 ( 
.A(n_16883),
.Y(n_17570)
);

NAND3xp33_ASAP7_75t_L g17571 ( 
.A(n_16742),
.B(n_10813),
.C(n_11860),
.Y(n_17571)
);

HB1xp67_ASAP7_75t_L g17572 ( 
.A(n_17233),
.Y(n_17572)
);

INVxp67_ASAP7_75t_L g17573 ( 
.A(n_16784),
.Y(n_17573)
);

INVxp67_ASAP7_75t_SL g17574 ( 
.A(n_17245),
.Y(n_17574)
);

INVx1_ASAP7_75t_L g17575 ( 
.A(n_16940),
.Y(n_17575)
);

INVx2_ASAP7_75t_L g17576 ( 
.A(n_17148),
.Y(n_17576)
);

INVx2_ASAP7_75t_L g17577 ( 
.A(n_17068),
.Y(n_17577)
);

OAI21xp5_ASAP7_75t_SL g17578 ( 
.A1(n_17171),
.A2(n_10038),
.B(n_10011),
.Y(n_17578)
);

INVx1_ASAP7_75t_L g17579 ( 
.A(n_16661),
.Y(n_17579)
);

INVx2_ASAP7_75t_L g17580 ( 
.A(n_17089),
.Y(n_17580)
);

HB1xp67_ASAP7_75t_L g17581 ( 
.A(n_17264),
.Y(n_17581)
);

INVx2_ASAP7_75t_L g17582 ( 
.A(n_16984),
.Y(n_17582)
);

AND2x2_ASAP7_75t_L g17583 ( 
.A(n_16823),
.B(n_11180),
.Y(n_17583)
);

OAI21x1_ASAP7_75t_L g17584 ( 
.A1(n_16824),
.A2(n_12082),
.B(n_12256),
.Y(n_17584)
);

INVxp67_ASAP7_75t_R g17585 ( 
.A(n_16819),
.Y(n_17585)
);

AND2x2_ASAP7_75t_L g17586 ( 
.A(n_17134),
.B(n_11180),
.Y(n_17586)
);

OR2x2_ASAP7_75t_L g17587 ( 
.A(n_16837),
.B(n_11202),
.Y(n_17587)
);

INVx2_ASAP7_75t_SL g17588 ( 
.A(n_17110),
.Y(n_17588)
);

INVx1_ASAP7_75t_L g17589 ( 
.A(n_17002),
.Y(n_17589)
);

INVx2_ASAP7_75t_L g17590 ( 
.A(n_17249),
.Y(n_17590)
);

AND2x4_ASAP7_75t_L g17591 ( 
.A(n_16985),
.B(n_10084),
.Y(n_17591)
);

INVx3_ASAP7_75t_L g17592 ( 
.A(n_16891),
.Y(n_17592)
);

INVx3_ASAP7_75t_L g17593 ( 
.A(n_16853),
.Y(n_17593)
);

INVx3_ASAP7_75t_L g17594 ( 
.A(n_16971),
.Y(n_17594)
);

INVx1_ASAP7_75t_SL g17595 ( 
.A(n_16818),
.Y(n_17595)
);

BUFx2_ASAP7_75t_L g17596 ( 
.A(n_17048),
.Y(n_17596)
);

INVx4_ASAP7_75t_L g17597 ( 
.A(n_16918),
.Y(n_17597)
);

INVx1_ASAP7_75t_L g17598 ( 
.A(n_16854),
.Y(n_17598)
);

AND2x2_ASAP7_75t_L g17599 ( 
.A(n_16978),
.B(n_11180),
.Y(n_17599)
);

OAI21x1_ASAP7_75t_L g17600 ( 
.A1(n_16943),
.A2(n_12336),
.B(n_12540),
.Y(n_17600)
);

INVxp67_ASAP7_75t_SL g17601 ( 
.A(n_17268),
.Y(n_17601)
);

INVx1_ASAP7_75t_L g17602 ( 
.A(n_16696),
.Y(n_17602)
);

BUFx2_ASAP7_75t_SL g17603 ( 
.A(n_16778),
.Y(n_17603)
);

INVx3_ASAP7_75t_L g17604 ( 
.A(n_16992),
.Y(n_17604)
);

INVx4_ASAP7_75t_SL g17605 ( 
.A(n_16795),
.Y(n_17605)
);

INVx2_ASAP7_75t_L g17606 ( 
.A(n_17256),
.Y(n_17606)
);

AOI21x1_ASAP7_75t_L g17607 ( 
.A1(n_16809),
.A2(n_13502),
.B(n_10956),
.Y(n_17607)
);

INVx2_ASAP7_75t_L g17608 ( 
.A(n_17156),
.Y(n_17608)
);

OAI21x1_ASAP7_75t_L g17609 ( 
.A1(n_17158),
.A2(n_12020),
.B(n_12016),
.Y(n_17609)
);

NAND2xp5_ASAP7_75t_SL g17610 ( 
.A(n_17288),
.B(n_10155),
.Y(n_17610)
);

NAND3xp33_ASAP7_75t_L g17611 ( 
.A(n_16793),
.B(n_10813),
.C(n_11860),
.Y(n_17611)
);

HB1xp67_ASAP7_75t_L g17612 ( 
.A(n_17203),
.Y(n_17612)
);

HB1xp67_ASAP7_75t_L g17613 ( 
.A(n_17172),
.Y(n_17613)
);

INVx1_ASAP7_75t_L g17614 ( 
.A(n_16697),
.Y(n_17614)
);

INVx1_ASAP7_75t_L g17615 ( 
.A(n_16812),
.Y(n_17615)
);

INVx1_ASAP7_75t_L g17616 ( 
.A(n_16729),
.Y(n_17616)
);

AND2x4_ASAP7_75t_L g17617 ( 
.A(n_16902),
.B(n_10084),
.Y(n_17617)
);

INVx1_ASAP7_75t_L g17618 ( 
.A(n_16735),
.Y(n_17618)
);

AOI21x1_ASAP7_75t_L g17619 ( 
.A1(n_16730),
.A2(n_13502),
.B(n_10956),
.Y(n_17619)
);

BUFx2_ASAP7_75t_L g17620 ( 
.A(n_17147),
.Y(n_17620)
);

INVxp67_ASAP7_75t_SL g17621 ( 
.A(n_16758),
.Y(n_17621)
);

BUFx12f_ASAP7_75t_L g17622 ( 
.A(n_16972),
.Y(n_17622)
);

INVx1_ASAP7_75t_L g17623 ( 
.A(n_16964),
.Y(n_17623)
);

OR2x2_ASAP7_75t_L g17624 ( 
.A(n_16744),
.B(n_11202),
.Y(n_17624)
);

INVx1_ASAP7_75t_L g17625 ( 
.A(n_17099),
.Y(n_17625)
);

HB1xp67_ASAP7_75t_L g17626 ( 
.A(n_17262),
.Y(n_17626)
);

INVx1_ASAP7_75t_L g17627 ( 
.A(n_17105),
.Y(n_17627)
);

OA21x2_ASAP7_75t_L g17628 ( 
.A1(n_17096),
.A2(n_10958),
.B(n_10941),
.Y(n_17628)
);

INVx1_ASAP7_75t_SL g17629 ( 
.A(n_17078),
.Y(n_17629)
);

INVx1_ASAP7_75t_L g17630 ( 
.A(n_17107),
.Y(n_17630)
);

NAND2xp5_ASAP7_75t_L g17631 ( 
.A(n_17252),
.B(n_10985),
.Y(n_17631)
);

INVx2_ASAP7_75t_SL g17632 ( 
.A(n_17093),
.Y(n_17632)
);

INVx1_ASAP7_75t_L g17633 ( 
.A(n_16847),
.Y(n_17633)
);

INVx1_ASAP7_75t_L g17634 ( 
.A(n_16849),
.Y(n_17634)
);

BUFx2_ASAP7_75t_L g17635 ( 
.A(n_17162),
.Y(n_17635)
);

INVx1_ASAP7_75t_L g17636 ( 
.A(n_16689),
.Y(n_17636)
);

INVx2_ASAP7_75t_L g17637 ( 
.A(n_17166),
.Y(n_17637)
);

AND2x2_ASAP7_75t_L g17638 ( 
.A(n_17282),
.B(n_11180),
.Y(n_17638)
);

OA21x2_ASAP7_75t_L g17639 ( 
.A1(n_17291),
.A2(n_10958),
.B(n_11158),
.Y(n_17639)
);

INVx6_ASAP7_75t_L g17640 ( 
.A(n_17285),
.Y(n_17640)
);

INVx1_ASAP7_75t_L g17641 ( 
.A(n_16871),
.Y(n_17641)
);

INVx1_ASAP7_75t_L g17642 ( 
.A(n_16800),
.Y(n_17642)
);

NAND3xp33_ASAP7_75t_L g17643 ( 
.A(n_17231),
.B(n_10813),
.C(n_11860),
.Y(n_17643)
);

OAI21x1_ASAP7_75t_L g17644 ( 
.A1(n_17070),
.A2(n_12054),
.B(n_11748),
.Y(n_17644)
);

OA21x2_ASAP7_75t_L g17645 ( 
.A1(n_17111),
.A2(n_11167),
.B(n_11162),
.Y(n_17645)
);

AND2x2_ASAP7_75t_L g17646 ( 
.A(n_17217),
.B(n_17036),
.Y(n_17646)
);

CKINVDCx20_ASAP7_75t_R g17647 ( 
.A(n_17157),
.Y(n_17647)
);

HB1xp67_ASAP7_75t_L g17648 ( 
.A(n_17119),
.Y(n_17648)
);

OR2x2_ASAP7_75t_L g17649 ( 
.A(n_16751),
.B(n_11202),
.Y(n_17649)
);

INVx2_ASAP7_75t_L g17650 ( 
.A(n_16973),
.Y(n_17650)
);

INVx2_ASAP7_75t_L g17651 ( 
.A(n_17170),
.Y(n_17651)
);

OA21x2_ASAP7_75t_L g17652 ( 
.A1(n_17200),
.A2(n_11168),
.B(n_11167),
.Y(n_17652)
);

INVx1_ASAP7_75t_L g17653 ( 
.A(n_16933),
.Y(n_17653)
);

INVxp67_ASAP7_75t_L g17654 ( 
.A(n_16791),
.Y(n_17654)
);

OA21x2_ASAP7_75t_L g17655 ( 
.A1(n_17259),
.A2(n_11173),
.B(n_11168),
.Y(n_17655)
);

INVx3_ASAP7_75t_R g17656 ( 
.A(n_17150),
.Y(n_17656)
);

BUFx2_ASAP7_75t_L g17657 ( 
.A(n_17153),
.Y(n_17657)
);

OAI21xp5_ASAP7_75t_L g17658 ( 
.A1(n_17173),
.A2(n_17269),
.B(n_16925),
.Y(n_17658)
);

NAND3xp33_ASAP7_75t_L g17659 ( 
.A(n_17240),
.B(n_17049),
.C(n_17260),
.Y(n_17659)
);

BUFx2_ASAP7_75t_L g17660 ( 
.A(n_17192),
.Y(n_17660)
);

INVx2_ASAP7_75t_L g17661 ( 
.A(n_17024),
.Y(n_17661)
);

NAND3xp33_ASAP7_75t_L g17662 ( 
.A(n_17265),
.B(n_11867),
.C(n_11837),
.Y(n_17662)
);

INVx1_ASAP7_75t_L g17663 ( 
.A(n_16934),
.Y(n_17663)
);

INVx1_ASAP7_75t_L g17664 ( 
.A(n_16935),
.Y(n_17664)
);

INVxp67_ASAP7_75t_L g17665 ( 
.A(n_17026),
.Y(n_17665)
);

INVx2_ASAP7_75t_L g17666 ( 
.A(n_17155),
.Y(n_17666)
);

INVx1_ASAP7_75t_L g17667 ( 
.A(n_16939),
.Y(n_17667)
);

INVxp67_ASAP7_75t_L g17668 ( 
.A(n_17196),
.Y(n_17668)
);

INVx2_ASAP7_75t_L g17669 ( 
.A(n_16903),
.Y(n_17669)
);

INVx1_ASAP7_75t_SL g17670 ( 
.A(n_17250),
.Y(n_17670)
);

NAND2xp5_ASAP7_75t_L g17671 ( 
.A(n_17013),
.B(n_10985),
.Y(n_17671)
);

BUFx3_ASAP7_75t_L g17672 ( 
.A(n_17003),
.Y(n_17672)
);

INVx1_ASAP7_75t_L g17673 ( 
.A(n_16949),
.Y(n_17673)
);

OR2x6_ASAP7_75t_L g17674 ( 
.A(n_16836),
.B(n_10027),
.Y(n_17674)
);

INVx1_ASAP7_75t_L g17675 ( 
.A(n_16950),
.Y(n_17675)
);

INVx1_ASAP7_75t_L g17676 ( 
.A(n_16750),
.Y(n_17676)
);

BUFx3_ASAP7_75t_L g17677 ( 
.A(n_17219),
.Y(n_17677)
);

NOR2x1p5_ASAP7_75t_L g17678 ( 
.A(n_16764),
.B(n_9092),
.Y(n_17678)
);

INVx1_ASAP7_75t_L g17679 ( 
.A(n_17204),
.Y(n_17679)
);

INVx4_ASAP7_75t_SL g17680 ( 
.A(n_16843),
.Y(n_17680)
);

BUFx3_ASAP7_75t_L g17681 ( 
.A(n_17021),
.Y(n_17681)
);

OA21x2_ASAP7_75t_L g17682 ( 
.A1(n_17270),
.A2(n_11186),
.B(n_11173),
.Y(n_17682)
);

INVxp67_ASAP7_75t_SL g17683 ( 
.A(n_16929),
.Y(n_17683)
);

AND2x2_ASAP7_75t_L g17684 ( 
.A(n_16805),
.B(n_11180),
.Y(n_17684)
);

AND2x2_ASAP7_75t_L g17685 ( 
.A(n_16858),
.B(n_11180),
.Y(n_17685)
);

INVxp67_ASAP7_75t_L g17686 ( 
.A(n_17176),
.Y(n_17686)
);

NAND2xp5_ASAP7_75t_L g17687 ( 
.A(n_17032),
.B(n_10985),
.Y(n_17687)
);

INVx2_ASAP7_75t_L g17688 ( 
.A(n_17124),
.Y(n_17688)
);

INVx2_ASAP7_75t_L g17689 ( 
.A(n_17169),
.Y(n_17689)
);

NAND2xp5_ASAP7_75t_SL g17690 ( 
.A(n_17186),
.B(n_10155),
.Y(n_17690)
);

INVx1_ASAP7_75t_L g17691 ( 
.A(n_17104),
.Y(n_17691)
);

INVx1_ASAP7_75t_L g17692 ( 
.A(n_16861),
.Y(n_17692)
);

INVx2_ASAP7_75t_L g17693 ( 
.A(n_17009),
.Y(n_17693)
);

AND2x2_ASAP7_75t_L g17694 ( 
.A(n_16862),
.B(n_16866),
.Y(n_17694)
);

INVx1_ASAP7_75t_L g17695 ( 
.A(n_16870),
.Y(n_17695)
);

AND2x2_ASAP7_75t_L g17696 ( 
.A(n_16869),
.B(n_11180),
.Y(n_17696)
);

INVx1_ASAP7_75t_L g17697 ( 
.A(n_16748),
.Y(n_17697)
);

INVx2_ASAP7_75t_L g17698 ( 
.A(n_17009),
.Y(n_17698)
);

INVx2_ASAP7_75t_L g17699 ( 
.A(n_17064),
.Y(n_17699)
);

INVx2_ASAP7_75t_L g17700 ( 
.A(n_17064),
.Y(n_17700)
);

NAND2xp5_ASAP7_75t_L g17701 ( 
.A(n_16887),
.B(n_10985),
.Y(n_17701)
);

INVx2_ASAP7_75t_L g17702 ( 
.A(n_17072),
.Y(n_17702)
);

HB1xp67_ASAP7_75t_L g17703 ( 
.A(n_17216),
.Y(n_17703)
);

INVx2_ASAP7_75t_L g17704 ( 
.A(n_17072),
.Y(n_17704)
);

AND2x2_ASAP7_75t_L g17705 ( 
.A(n_16894),
.B(n_11198),
.Y(n_17705)
);

INVx4_ASAP7_75t_L g17706 ( 
.A(n_16844),
.Y(n_17706)
);

INVx1_ASAP7_75t_L g17707 ( 
.A(n_17005),
.Y(n_17707)
);

INVx1_ASAP7_75t_L g17708 ( 
.A(n_17008),
.Y(n_17708)
);

BUFx2_ASAP7_75t_L g17709 ( 
.A(n_17230),
.Y(n_17709)
);

INVx1_ASAP7_75t_L g17710 ( 
.A(n_17010),
.Y(n_17710)
);

INVx1_ASAP7_75t_L g17711 ( 
.A(n_17012),
.Y(n_17711)
);

INVx2_ASAP7_75t_SL g17712 ( 
.A(n_17023),
.Y(n_17712)
);

AND2x2_ASAP7_75t_L g17713 ( 
.A(n_16897),
.B(n_11198),
.Y(n_17713)
);

AND2x4_ASAP7_75t_L g17714 ( 
.A(n_16889),
.B(n_10084),
.Y(n_17714)
);

INVx1_ASAP7_75t_L g17715 ( 
.A(n_17017),
.Y(n_17715)
);

NAND2xp5_ASAP7_75t_L g17716 ( 
.A(n_17019),
.B(n_10985),
.Y(n_17716)
);

INVx1_ASAP7_75t_L g17717 ( 
.A(n_16956),
.Y(n_17717)
);

AND2x2_ASAP7_75t_L g17718 ( 
.A(n_17278),
.B(n_11198),
.Y(n_17718)
);

INVx1_ASAP7_75t_L g17719 ( 
.A(n_16957),
.Y(n_17719)
);

BUFx2_ASAP7_75t_L g17720 ( 
.A(n_17242),
.Y(n_17720)
);

INVx2_ASAP7_75t_L g17721 ( 
.A(n_16898),
.Y(n_17721)
);

INVx2_ASAP7_75t_L g17722 ( 
.A(n_16899),
.Y(n_17722)
);

INVx1_ASAP7_75t_L g17723 ( 
.A(n_16962),
.Y(n_17723)
);

INVx1_ASAP7_75t_L g17724 ( 
.A(n_16963),
.Y(n_17724)
);

OR2x2_ASAP7_75t_L g17725 ( 
.A(n_16875),
.B(n_11202),
.Y(n_17725)
);

INVx2_ASAP7_75t_SL g17726 ( 
.A(n_17015),
.Y(n_17726)
);

HB1xp67_ASAP7_75t_L g17727 ( 
.A(n_17199),
.Y(n_17727)
);

INVx1_ASAP7_75t_L g17728 ( 
.A(n_16975),
.Y(n_17728)
);

INVx1_ASAP7_75t_L g17729 ( 
.A(n_17014),
.Y(n_17729)
);

HB1xp67_ASAP7_75t_L g17730 ( 
.A(n_17208),
.Y(n_17730)
);

INVx2_ASAP7_75t_L g17731 ( 
.A(n_16907),
.Y(n_17731)
);

HB1xp67_ASAP7_75t_L g17732 ( 
.A(n_16966),
.Y(n_17732)
);

INVxp67_ASAP7_75t_L g17733 ( 
.A(n_17225),
.Y(n_17733)
);

AND2x2_ASAP7_75t_L g17734 ( 
.A(n_17277),
.B(n_11198),
.Y(n_17734)
);

BUFx3_ASAP7_75t_L g17735 ( 
.A(n_16905),
.Y(n_17735)
);

OA21x2_ASAP7_75t_L g17736 ( 
.A1(n_17272),
.A2(n_11190),
.B(n_11186),
.Y(n_17736)
);

INVx2_ASAP7_75t_L g17737 ( 
.A(n_16908),
.Y(n_17737)
);

NAND2xp5_ASAP7_75t_L g17738 ( 
.A(n_17091),
.B(n_10985),
.Y(n_17738)
);

INVx2_ASAP7_75t_L g17739 ( 
.A(n_16910),
.Y(n_17739)
);

INVxp67_ASAP7_75t_SL g17740 ( 
.A(n_17234),
.Y(n_17740)
);

INVx1_ASAP7_75t_L g17741 ( 
.A(n_17092),
.Y(n_17741)
);

NAND3xp33_ASAP7_75t_L g17742 ( 
.A(n_16952),
.B(n_11867),
.C(n_11833),
.Y(n_17742)
);

AND2x2_ASAP7_75t_L g17743 ( 
.A(n_17201),
.B(n_11198),
.Y(n_17743)
);

INVx1_ASAP7_75t_L g17744 ( 
.A(n_17094),
.Y(n_17744)
);

NAND2xp5_ASAP7_75t_SL g17745 ( 
.A(n_17186),
.B(n_10155),
.Y(n_17745)
);

NAND3xp33_ASAP7_75t_L g17746 ( 
.A(n_16757),
.B(n_11867),
.C(n_11833),
.Y(n_17746)
);

AND2x2_ASAP7_75t_L g17747 ( 
.A(n_17054),
.B(n_11198),
.Y(n_17747)
);

BUFx2_ASAP7_75t_L g17748 ( 
.A(n_17000),
.Y(n_17748)
);

NOR2x1_ASAP7_75t_SL g17749 ( 
.A(n_17062),
.B(n_17065),
.Y(n_17749)
);

NOR2xp33_ASAP7_75t_L g17750 ( 
.A(n_16717),
.B(n_16912),
.Y(n_17750)
);

INVx2_ASAP7_75t_L g17751 ( 
.A(n_16913),
.Y(n_17751)
);

INVx1_ASAP7_75t_L g17752 ( 
.A(n_17095),
.Y(n_17752)
);

AND2x2_ASAP7_75t_L g17753 ( 
.A(n_17253),
.B(n_11198),
.Y(n_17753)
);

NAND2xp5_ASAP7_75t_L g17754 ( 
.A(n_17103),
.B(n_11176),
.Y(n_17754)
);

INVx1_ASAP7_75t_L g17755 ( 
.A(n_17130),
.Y(n_17755)
);

INVx2_ASAP7_75t_L g17756 ( 
.A(n_16920),
.Y(n_17756)
);

INVx1_ASAP7_75t_L g17757 ( 
.A(n_17131),
.Y(n_17757)
);

NAND3xp33_ASAP7_75t_SL g17758 ( 
.A(n_16877),
.B(n_10038),
.C(n_10011),
.Y(n_17758)
);

INVx1_ASAP7_75t_L g17759 ( 
.A(n_16915),
.Y(n_17759)
);

NAND2xp5_ASAP7_75t_L g17760 ( 
.A(n_16766),
.B(n_11176),
.Y(n_17760)
);

INVx1_ASAP7_75t_L g17761 ( 
.A(n_16922),
.Y(n_17761)
);

INVx2_ASAP7_75t_L g17762 ( 
.A(n_17149),
.Y(n_17762)
);

HB1xp67_ASAP7_75t_L g17763 ( 
.A(n_17187),
.Y(n_17763)
);

INVx2_ASAP7_75t_L g17764 ( 
.A(n_16860),
.Y(n_17764)
);

AND2x2_ASAP7_75t_L g17765 ( 
.A(n_17254),
.B(n_11337),
.Y(n_17765)
);

INVx2_ASAP7_75t_L g17766 ( 
.A(n_16863),
.Y(n_17766)
);

INVx4_ASAP7_75t_SL g17767 ( 
.A(n_16876),
.Y(n_17767)
);

INVx1_ASAP7_75t_L g17768 ( 
.A(n_17109),
.Y(n_17768)
);

OR2x2_ASAP7_75t_SL g17769 ( 
.A(n_17237),
.B(n_11833),
.Y(n_17769)
);

INVx2_ASAP7_75t_L g17770 ( 
.A(n_16865),
.Y(n_17770)
);

INVx1_ASAP7_75t_L g17771 ( 
.A(n_16880),
.Y(n_17771)
);

INVx1_ASAP7_75t_L g17772 ( 
.A(n_17112),
.Y(n_17772)
);

INVx3_ASAP7_75t_L g17773 ( 
.A(n_17006),
.Y(n_17773)
);

NAND3xp33_ASAP7_75t_L g17774 ( 
.A(n_16769),
.B(n_10026),
.C(n_10007),
.Y(n_17774)
);

INVx1_ASAP7_75t_L g17775 ( 
.A(n_17116),
.Y(n_17775)
);

INVx1_ASAP7_75t_L g17776 ( 
.A(n_17117),
.Y(n_17776)
);

NOR2xp33_ASAP7_75t_L g17777 ( 
.A(n_16773),
.B(n_10159),
.Y(n_17777)
);

INVx4_ASAP7_75t_SL g17778 ( 
.A(n_16774),
.Y(n_17778)
);

NAND3xp33_ASAP7_75t_L g17779 ( 
.A(n_16776),
.B(n_10026),
.C(n_10007),
.Y(n_17779)
);

OAI21xp5_ASAP7_75t_L g17780 ( 
.A1(n_16878),
.A2(n_16909),
.B(n_17235),
.Y(n_17780)
);

AND2x2_ASAP7_75t_L g17781 ( 
.A(n_17209),
.B(n_11337),
.Y(n_17781)
);

AND2x2_ASAP7_75t_L g17782 ( 
.A(n_17258),
.B(n_11337),
.Y(n_17782)
);

OAI21xp5_ASAP7_75t_L g17783 ( 
.A1(n_17284),
.A2(n_17177),
.B(n_17202),
.Y(n_17783)
);

INVx1_ASAP7_75t_L g17784 ( 
.A(n_17118),
.Y(n_17784)
);

NAND2xp5_ASAP7_75t_SL g17785 ( 
.A(n_17202),
.B(n_10155),
.Y(n_17785)
);

OR2x2_ASAP7_75t_SL g17786 ( 
.A(n_16995),
.B(n_10748),
.Y(n_17786)
);

NAND3xp33_ASAP7_75t_SL g17787 ( 
.A(n_16782),
.B(n_10038),
.C(n_10011),
.Y(n_17787)
);

INVx2_ASAP7_75t_SL g17788 ( 
.A(n_17034),
.Y(n_17788)
);

INVx2_ASAP7_75t_L g17789 ( 
.A(n_17043),
.Y(n_17789)
);

OAI21x1_ASAP7_75t_L g17790 ( 
.A1(n_17038),
.A2(n_11767),
.B(n_11765),
.Y(n_17790)
);

OA21x2_ASAP7_75t_L g17791 ( 
.A1(n_16955),
.A2(n_11204),
.B(n_11190),
.Y(n_17791)
);

INVx2_ASAP7_75t_SL g17792 ( 
.A(n_16997),
.Y(n_17792)
);

INVx2_ASAP7_75t_L g17793 ( 
.A(n_17128),
.Y(n_17793)
);

INVx1_ASAP7_75t_L g17794 ( 
.A(n_17123),
.Y(n_17794)
);

HB1xp67_ASAP7_75t_L g17795 ( 
.A(n_17177),
.Y(n_17795)
);

OR2x6_ASAP7_75t_L g17796 ( 
.A(n_16790),
.B(n_10027),
.Y(n_17796)
);

INVxp67_ASAP7_75t_L g17797 ( 
.A(n_17047),
.Y(n_17797)
);

AND2x2_ASAP7_75t_L g17798 ( 
.A(n_17138),
.B(n_11337),
.Y(n_17798)
);

INVx2_ASAP7_75t_L g17799 ( 
.A(n_17128),
.Y(n_17799)
);

INVx2_ASAP7_75t_L g17800 ( 
.A(n_16970),
.Y(n_17800)
);

INVx2_ASAP7_75t_L g17801 ( 
.A(n_17122),
.Y(n_17801)
);

BUFx2_ASAP7_75t_L g17802 ( 
.A(n_16873),
.Y(n_17802)
);

INVx2_ASAP7_75t_L g17803 ( 
.A(n_17175),
.Y(n_17803)
);

INVx2_ASAP7_75t_L g17804 ( 
.A(n_17178),
.Y(n_17804)
);

INVx2_ASAP7_75t_L g17805 ( 
.A(n_17165),
.Y(n_17805)
);

INVxp67_ASAP7_75t_SL g17806 ( 
.A(n_17181),
.Y(n_17806)
);

INVx4_ASAP7_75t_SL g17807 ( 
.A(n_17142),
.Y(n_17807)
);

NAND2xp5_ASAP7_75t_L g17808 ( 
.A(n_17132),
.B(n_11176),
.Y(n_17808)
);

NAND2xp5_ASAP7_75t_SL g17809 ( 
.A(n_17224),
.B(n_10155),
.Y(n_17809)
);

BUFx2_ASAP7_75t_SL g17810 ( 
.A(n_17159),
.Y(n_17810)
);

INVx1_ASAP7_75t_L g17811 ( 
.A(n_17125),
.Y(n_17811)
);

OAI21x1_ASAP7_75t_L g17812 ( 
.A1(n_17152),
.A2(n_11819),
.B(n_12599),
.Y(n_17812)
);

HB1xp67_ASAP7_75t_L g17813 ( 
.A(n_16958),
.Y(n_17813)
);

INVx5_ASAP7_75t_L g17814 ( 
.A(n_17179),
.Y(n_17814)
);

INVx4_ASAP7_75t_L g17815 ( 
.A(n_17145),
.Y(n_17815)
);

INVx2_ASAP7_75t_L g17816 ( 
.A(n_17167),
.Y(n_17816)
);

INVx2_ASAP7_75t_L g17817 ( 
.A(n_16945),
.Y(n_17817)
);

INVx3_ASAP7_75t_L g17818 ( 
.A(n_17007),
.Y(n_17818)
);

INVx4_ASAP7_75t_L g17819 ( 
.A(n_17154),
.Y(n_17819)
);

INVx2_ASAP7_75t_L g17820 ( 
.A(n_17031),
.Y(n_17820)
);

INVx2_ASAP7_75t_L g17821 ( 
.A(n_17247),
.Y(n_17821)
);

BUFx8_ASAP7_75t_L g17822 ( 
.A(n_17161),
.Y(n_17822)
);

AND2x2_ASAP7_75t_L g17823 ( 
.A(n_16988),
.B(n_11337),
.Y(n_17823)
);

INVx1_ASAP7_75t_L g17824 ( 
.A(n_16991),
.Y(n_17824)
);

INVx1_ASAP7_75t_L g17825 ( 
.A(n_16994),
.Y(n_17825)
);

INVx1_ASAP7_75t_L g17826 ( 
.A(n_16996),
.Y(n_17826)
);

AOI21xp5_ASAP7_75t_L g17827 ( 
.A1(n_17274),
.A2(n_11698),
.B(n_11679),
.Y(n_17827)
);

INVx1_ASAP7_75t_L g17828 ( 
.A(n_17001),
.Y(n_17828)
);

INVx2_ASAP7_75t_L g17829 ( 
.A(n_17214),
.Y(n_17829)
);

INVxp67_ASAP7_75t_SL g17830 ( 
.A(n_17004),
.Y(n_17830)
);

BUFx2_ASAP7_75t_L g17831 ( 
.A(n_17085),
.Y(n_17831)
);

INVx1_ASAP7_75t_SL g17832 ( 
.A(n_17221),
.Y(n_17832)
);

BUFx3_ASAP7_75t_L g17833 ( 
.A(n_17126),
.Y(n_17833)
);

INVx1_ASAP7_75t_L g17834 ( 
.A(n_17083),
.Y(n_17834)
);

INVx1_ASAP7_75t_SL g17835 ( 
.A(n_17211),
.Y(n_17835)
);

INVx2_ASAP7_75t_L g17836 ( 
.A(n_17033),
.Y(n_17836)
);

BUFx2_ASAP7_75t_L g17837 ( 
.A(n_17087),
.Y(n_17837)
);

INVx1_ASAP7_75t_L g17838 ( 
.A(n_17088),
.Y(n_17838)
);

INVx1_ASAP7_75t_L g17839 ( 
.A(n_17029),
.Y(n_17839)
);

BUFx3_ASAP7_75t_L g17840 ( 
.A(n_17030),
.Y(n_17840)
);

AND2x4_ASAP7_75t_L g17841 ( 
.A(n_17041),
.B(n_10084),
.Y(n_17841)
);

INVx2_ASAP7_75t_L g17842 ( 
.A(n_17229),
.Y(n_17842)
);

INVx1_ASAP7_75t_SL g17843 ( 
.A(n_16874),
.Y(n_17843)
);

HB1xp67_ASAP7_75t_L g17844 ( 
.A(n_16900),
.Y(n_17844)
);

OA21x2_ASAP7_75t_L g17845 ( 
.A1(n_17058),
.A2(n_11211),
.B(n_11204),
.Y(n_17845)
);

INVxp67_ASAP7_75t_L g17846 ( 
.A(n_17050),
.Y(n_17846)
);

INVx2_ASAP7_75t_L g17847 ( 
.A(n_16959),
.Y(n_17847)
);

AND2x4_ASAP7_75t_SL g17848 ( 
.A(n_16924),
.B(n_8124),
.Y(n_17848)
);

INVx1_ASAP7_75t_L g17849 ( 
.A(n_17055),
.Y(n_17849)
);

INVx2_ASAP7_75t_L g17850 ( 
.A(n_16960),
.Y(n_17850)
);

INVx1_ASAP7_75t_L g17851 ( 
.A(n_17059),
.Y(n_17851)
);

INVx4_ASAP7_75t_SL g17852 ( 
.A(n_17163),
.Y(n_17852)
);

INVx1_ASAP7_75t_L g17853 ( 
.A(n_17060),
.Y(n_17853)
);

OAI21x1_ASAP7_75t_L g17854 ( 
.A1(n_17239),
.A2(n_12638),
.B(n_12598),
.Y(n_17854)
);

INVx3_ASAP7_75t_L g17855 ( 
.A(n_16927),
.Y(n_17855)
);

NOR2xp33_ASAP7_75t_L g17856 ( 
.A(n_17061),
.B(n_10159),
.Y(n_17856)
);

OA21x2_ASAP7_75t_L g17857 ( 
.A1(n_17220),
.A2(n_11233),
.B(n_11211),
.Y(n_17857)
);

INVx2_ASAP7_75t_L g17858 ( 
.A(n_16965),
.Y(n_17858)
);

INVx2_ASAP7_75t_L g17859 ( 
.A(n_16968),
.Y(n_17859)
);

BUFx2_ASAP7_75t_L g17860 ( 
.A(n_17063),
.Y(n_17860)
);

INVx1_ASAP7_75t_L g17861 ( 
.A(n_17067),
.Y(n_17861)
);

INVx2_ASAP7_75t_L g17862 ( 
.A(n_17197),
.Y(n_17862)
);

AND2x4_ASAP7_75t_L g17863 ( 
.A(n_17071),
.B(n_17074),
.Y(n_17863)
);

INVx2_ASAP7_75t_L g17864 ( 
.A(n_16906),
.Y(n_17864)
);

AOI21xp5_ASAP7_75t_L g17865 ( 
.A1(n_16917),
.A2(n_11698),
.B(n_11679),
.Y(n_17865)
);

INVx1_ASAP7_75t_L g17866 ( 
.A(n_17080),
.Y(n_17866)
);

INVx1_ASAP7_75t_L g17867 ( 
.A(n_17082),
.Y(n_17867)
);

INVx1_ASAP7_75t_L g17868 ( 
.A(n_17174),
.Y(n_17868)
);

INVx2_ASAP7_75t_SL g17869 ( 
.A(n_16953),
.Y(n_17869)
);

OA21x2_ASAP7_75t_L g17870 ( 
.A1(n_17129),
.A2(n_11244),
.B(n_11233),
.Y(n_17870)
);

INVx1_ASAP7_75t_L g17871 ( 
.A(n_17182),
.Y(n_17871)
);

BUFx2_ASAP7_75t_L g17872 ( 
.A(n_17267),
.Y(n_17872)
);

OR2x6_ASAP7_75t_L g17873 ( 
.A(n_17185),
.B(n_10027),
.Y(n_17873)
);

INVx2_ASAP7_75t_L g17874 ( 
.A(n_17180),
.Y(n_17874)
);

NAND2xp5_ASAP7_75t_L g17875 ( 
.A(n_17188),
.B(n_11176),
.Y(n_17875)
);

AND2x2_ASAP7_75t_L g17876 ( 
.A(n_17011),
.B(n_11337),
.Y(n_17876)
);

HB1xp67_ASAP7_75t_L g17877 ( 
.A(n_17207),
.Y(n_17877)
);

INVx2_ASAP7_75t_L g17878 ( 
.A(n_17018),
.Y(n_17878)
);

AND2x2_ASAP7_75t_L g17879 ( 
.A(n_17275),
.B(n_16937),
.Y(n_17879)
);

INVx2_ASAP7_75t_L g17880 ( 
.A(n_17039),
.Y(n_17880)
);

BUFx2_ASAP7_75t_L g17881 ( 
.A(n_16923),
.Y(n_17881)
);

INVx1_ASAP7_75t_L g17882 ( 
.A(n_16986),
.Y(n_17882)
);

OR2x2_ASAP7_75t_L g17883 ( 
.A(n_17127),
.B(n_10754),
.Y(n_17883)
);

HB1xp67_ASAP7_75t_L g17884 ( 
.A(n_17183),
.Y(n_17884)
);

INVx1_ASAP7_75t_L g17885 ( 
.A(n_16993),
.Y(n_17885)
);

NAND2xp5_ASAP7_75t_L g17886 ( 
.A(n_16983),
.B(n_17193),
.Y(n_17886)
);

NOR3xp33_ASAP7_75t_L g17887 ( 
.A(n_17136),
.B(n_10023),
.C(n_9993),
.Y(n_17887)
);

INVx1_ASAP7_75t_L g17888 ( 
.A(n_16938),
.Y(n_17888)
);

AND2x2_ASAP7_75t_L g17889 ( 
.A(n_17016),
.B(n_17086),
.Y(n_17889)
);

INVx1_ASAP7_75t_L g17890 ( 
.A(n_16944),
.Y(n_17890)
);

OR2x2_ASAP7_75t_L g17891 ( 
.A(n_17301),
.B(n_16946),
.Y(n_17891)
);

AND2x4_ASAP7_75t_L g17892 ( 
.A(n_17338),
.B(n_17098),
.Y(n_17892)
);

AND2x2_ASAP7_75t_L g17893 ( 
.A(n_17293),
.B(n_17100),
.Y(n_17893)
);

INVx1_ASAP7_75t_L g17894 ( 
.A(n_17352),
.Y(n_17894)
);

INVx1_ASAP7_75t_L g17895 ( 
.A(n_17321),
.Y(n_17895)
);

INVx1_ASAP7_75t_L g17896 ( 
.A(n_17404),
.Y(n_17896)
);

AND2x2_ASAP7_75t_L g17897 ( 
.A(n_17585),
.B(n_17101),
.Y(n_17897)
);

INVx1_ASAP7_75t_L g17898 ( 
.A(n_17294),
.Y(n_17898)
);

INVx1_ASAP7_75t_L g17899 ( 
.A(n_17295),
.Y(n_17899)
);

INVx2_ASAP7_75t_L g17900 ( 
.A(n_17434),
.Y(n_17900)
);

NOR2xp33_ASAP7_75t_L g17901 ( 
.A(n_17367),
.B(n_17191),
.Y(n_17901)
);

OR2x2_ASAP7_75t_L g17902 ( 
.A(n_17436),
.B(n_17028),
.Y(n_17902)
);

AND2x2_ASAP7_75t_L g17903 ( 
.A(n_17396),
.B(n_17279),
.Y(n_17903)
);

NOR2xp67_ASAP7_75t_R g17904 ( 
.A(n_17538),
.B(n_17554),
.Y(n_17904)
);

NAND2xp5_ASAP7_75t_L g17905 ( 
.A(n_17371),
.B(n_17133),
.Y(n_17905)
);

AND2x2_ASAP7_75t_L g17906 ( 
.A(n_17395),
.B(n_17044),
.Y(n_17906)
);

INVx2_ASAP7_75t_L g17907 ( 
.A(n_17434),
.Y(n_17907)
);

AOI22xp5_ASAP7_75t_L g17908 ( 
.A1(n_17344),
.A2(n_17263),
.B1(n_17280),
.B2(n_17273),
.Y(n_17908)
);

OR2x2_ASAP7_75t_L g17909 ( 
.A(n_17336),
.B(n_17337),
.Y(n_17909)
);

INVx1_ASAP7_75t_L g17910 ( 
.A(n_17300),
.Y(n_17910)
);

INVx1_ASAP7_75t_L g17911 ( 
.A(n_17363),
.Y(n_17911)
);

INVx1_ASAP7_75t_L g17912 ( 
.A(n_17323),
.Y(n_17912)
);

NAND3xp33_ASAP7_75t_L g17913 ( 
.A(n_17359),
.B(n_17195),
.C(n_17184),
.Y(n_17913)
);

BUFx2_ASAP7_75t_L g17914 ( 
.A(n_17647),
.Y(n_17914)
);

AND2x2_ASAP7_75t_L g17915 ( 
.A(n_17322),
.B(n_17066),
.Y(n_17915)
);

AND3x2_ASAP7_75t_L g17916 ( 
.A(n_17474),
.B(n_17133),
.C(n_17283),
.Y(n_17916)
);

INVx1_ASAP7_75t_L g17917 ( 
.A(n_17319),
.Y(n_17917)
);

BUFx3_ASAP7_75t_L g17918 ( 
.A(n_17358),
.Y(n_17918)
);

INVx2_ASAP7_75t_L g17919 ( 
.A(n_17749),
.Y(n_17919)
);

AND2x2_ASAP7_75t_L g17920 ( 
.A(n_17298),
.B(n_17075),
.Y(n_17920)
);

INVx2_ASAP7_75t_L g17921 ( 
.A(n_17538),
.Y(n_17921)
);

AND2x2_ASAP7_75t_L g17922 ( 
.A(n_17426),
.B(n_17079),
.Y(n_17922)
);

INVx1_ASAP7_75t_SL g17923 ( 
.A(n_17428),
.Y(n_17923)
);

INVx2_ASAP7_75t_L g17924 ( 
.A(n_17554),
.Y(n_17924)
);

AND2x2_ASAP7_75t_L g17925 ( 
.A(n_17385),
.B(n_17362),
.Y(n_17925)
);

INVx1_ASAP7_75t_L g17926 ( 
.A(n_17430),
.Y(n_17926)
);

NAND2xp5_ASAP7_75t_L g17927 ( 
.A(n_17500),
.B(n_17084),
.Y(n_17927)
);

NAND2x1p5_ASAP7_75t_L g17928 ( 
.A(n_17390),
.B(n_17261),
.Y(n_17928)
);

AOI22xp5_ASAP7_75t_L g17929 ( 
.A1(n_17335),
.A2(n_17361),
.B1(n_17553),
.B2(n_17621),
.Y(n_17929)
);

INVx1_ASAP7_75t_L g17930 ( 
.A(n_17406),
.Y(n_17930)
);

INVx1_ASAP7_75t_L g17931 ( 
.A(n_17406),
.Y(n_17931)
);

NAND2xp5_ASAP7_75t_L g17932 ( 
.A(n_17564),
.B(n_17106),
.Y(n_17932)
);

INVx1_ASAP7_75t_L g17933 ( 
.A(n_17424),
.Y(n_17933)
);

INVx2_ASAP7_75t_L g17934 ( 
.A(n_17309),
.Y(n_17934)
);

INVx1_ASAP7_75t_L g17935 ( 
.A(n_17424),
.Y(n_17935)
);

INVx1_ASAP7_75t_SL g17936 ( 
.A(n_17469),
.Y(n_17936)
);

AND2x2_ASAP7_75t_L g17937 ( 
.A(n_17429),
.B(n_17386),
.Y(n_17937)
);

NAND2xp5_ASAP7_75t_L g17938 ( 
.A(n_17310),
.B(n_17108),
.Y(n_17938)
);

HB1xp67_ASAP7_75t_L g17939 ( 
.A(n_17341),
.Y(n_17939)
);

INVx1_ASAP7_75t_L g17940 ( 
.A(n_17497),
.Y(n_17940)
);

OR2x2_ASAP7_75t_L g17941 ( 
.A(n_17376),
.B(n_17276),
.Y(n_17941)
);

OR2x2_ASAP7_75t_L g17942 ( 
.A(n_17377),
.B(n_17241),
.Y(n_17942)
);

NAND2xp5_ASAP7_75t_L g17943 ( 
.A(n_17473),
.B(n_17492),
.Y(n_17943)
);

AND2x2_ASAP7_75t_L g17944 ( 
.A(n_17346),
.B(n_17115),
.Y(n_17944)
);

INVx1_ASAP7_75t_L g17945 ( 
.A(n_17504),
.Y(n_17945)
);

INVx1_ASAP7_75t_L g17946 ( 
.A(n_17505),
.Y(n_17946)
);

INVx2_ASAP7_75t_L g17947 ( 
.A(n_17334),
.Y(n_17947)
);

OR2x6_ASAP7_75t_L g17948 ( 
.A(n_17603),
.B(n_16981),
.Y(n_17948)
);

AND2x2_ASAP7_75t_L g17949 ( 
.A(n_17560),
.B(n_17139),
.Y(n_17949)
);

INVx1_ASAP7_75t_L g17950 ( 
.A(n_17535),
.Y(n_17950)
);

OR2x2_ASAP7_75t_L g17951 ( 
.A(n_17399),
.B(n_17232),
.Y(n_17951)
);

AND2x2_ASAP7_75t_L g17952 ( 
.A(n_17366),
.B(n_17140),
.Y(n_17952)
);

OR2x2_ASAP7_75t_L g17953 ( 
.A(n_17479),
.B(n_17287),
.Y(n_17953)
);

INVx1_ASAP7_75t_SL g17954 ( 
.A(n_17491),
.Y(n_17954)
);

AND2x2_ASAP7_75t_L g17955 ( 
.A(n_17357),
.B(n_17190),
.Y(n_17955)
);

INVx1_ASAP7_75t_L g17956 ( 
.A(n_17454),
.Y(n_17956)
);

AND2x2_ASAP7_75t_L g17957 ( 
.A(n_17379),
.B(n_17222),
.Y(n_17957)
);

OR2x2_ASAP7_75t_L g17958 ( 
.A(n_17484),
.B(n_17081),
.Y(n_17958)
);

AND2x4_ASAP7_75t_L g17959 ( 
.A(n_17476),
.B(n_17226),
.Y(n_17959)
);

INVx2_ASAP7_75t_L g17960 ( 
.A(n_17380),
.Y(n_17960)
);

OR2x2_ASAP7_75t_L g17961 ( 
.A(n_17432),
.B(n_17206),
.Y(n_17961)
);

AOI21xp33_ASAP7_75t_L g17962 ( 
.A1(n_17549),
.A2(n_17248),
.B(n_17210),
.Y(n_17962)
);

INVx2_ASAP7_75t_L g17963 ( 
.A(n_17393),
.Y(n_17963)
);

HB1xp67_ASAP7_75t_L g17964 ( 
.A(n_17356),
.Y(n_17964)
);

INVx1_ASAP7_75t_L g17965 ( 
.A(n_17454),
.Y(n_17965)
);

INVxp67_ASAP7_75t_L g17966 ( 
.A(n_17763),
.Y(n_17966)
);

AND2x2_ASAP7_75t_L g17967 ( 
.A(n_17884),
.B(n_17223),
.Y(n_17967)
);

AND2x4_ASAP7_75t_L g17968 ( 
.A(n_17476),
.B(n_17212),
.Y(n_17968)
);

OR2x2_ASAP7_75t_L g17969 ( 
.A(n_17330),
.B(n_17143),
.Y(n_17969)
);

INVx1_ASAP7_75t_L g17970 ( 
.A(n_17464),
.Y(n_17970)
);

HB1xp67_ASAP7_75t_L g17971 ( 
.A(n_17542),
.Y(n_17971)
);

OR2x2_ASAP7_75t_L g17972 ( 
.A(n_17410),
.B(n_17035),
.Y(n_17972)
);

AND2x4_ASAP7_75t_SL g17973 ( 
.A(n_17597),
.B(n_17213),
.Y(n_17973)
);

INVx1_ASAP7_75t_L g17974 ( 
.A(n_17464),
.Y(n_17974)
);

AND2x2_ASAP7_75t_L g17975 ( 
.A(n_17407),
.B(n_17228),
.Y(n_17975)
);

AND2x2_ASAP7_75t_L g17976 ( 
.A(n_17407),
.B(n_17215),
.Y(n_17976)
);

OR2x2_ASAP7_75t_L g17977 ( 
.A(n_17418),
.B(n_17042),
.Y(n_17977)
);

INVx2_ASAP7_75t_SL g17978 ( 
.A(n_17814),
.Y(n_17978)
);

INVx2_ASAP7_75t_L g17979 ( 
.A(n_17786),
.Y(n_17979)
);

AND2x2_ASAP7_75t_L g17980 ( 
.A(n_17551),
.B(n_17227),
.Y(n_17980)
);

HB1xp67_ASAP7_75t_L g17981 ( 
.A(n_17506),
.Y(n_17981)
);

INVx1_ASAP7_75t_L g17982 ( 
.A(n_17364),
.Y(n_17982)
);

INVx1_ASAP7_75t_L g17983 ( 
.A(n_17409),
.Y(n_17983)
);

AND2x2_ASAP7_75t_L g17984 ( 
.A(n_17382),
.B(n_17243),
.Y(n_17984)
);

BUFx2_ASAP7_75t_L g17985 ( 
.A(n_17450),
.Y(n_17985)
);

AND2x2_ASAP7_75t_L g17986 ( 
.A(n_17381),
.B(n_17045),
.Y(n_17986)
);

AND2x2_ASAP7_75t_L g17987 ( 
.A(n_17398),
.B(n_17052),
.Y(n_17987)
);

AND2x2_ASAP7_75t_L g17988 ( 
.A(n_17405),
.B(n_17053),
.Y(n_17988)
);

OR2x2_ASAP7_75t_L g17989 ( 
.A(n_17365),
.B(n_17090),
.Y(n_17989)
);

AND2x2_ASAP7_75t_L g17990 ( 
.A(n_17408),
.B(n_17137),
.Y(n_17990)
);

INVx3_ASAP7_75t_L g17991 ( 
.A(n_17368),
.Y(n_17991)
);

OR2x2_ASAP7_75t_L g17992 ( 
.A(n_17369),
.B(n_17370),
.Y(n_17992)
);

INVx1_ASAP7_75t_L g17993 ( 
.A(n_17703),
.Y(n_17993)
);

INVx1_ASAP7_75t_L g17994 ( 
.A(n_17354),
.Y(n_17994)
);

AND2x2_ASAP7_75t_L g17995 ( 
.A(n_17488),
.B(n_17517),
.Y(n_17995)
);

AND2x2_ASAP7_75t_L g17996 ( 
.A(n_17438),
.B(n_17141),
.Y(n_17996)
);

AND2x4_ASAP7_75t_L g17997 ( 
.A(n_17439),
.B(n_17168),
.Y(n_17997)
);

NAND2xp5_ASAP7_75t_L g17998 ( 
.A(n_17595),
.B(n_11176),
.Y(n_17998)
);

AND2x4_ASAP7_75t_L g17999 ( 
.A(n_17452),
.B(n_11337),
.Y(n_17999)
);

INVx1_ASAP7_75t_L g18000 ( 
.A(n_17355),
.Y(n_18000)
);

AND2x2_ASAP7_75t_L g18001 ( 
.A(n_17709),
.B(n_11433),
.Y(n_18001)
);

NOR2xp33_ASAP7_75t_L g18002 ( 
.A(n_17573),
.B(n_10159),
.Y(n_18002)
);

INVx2_ASAP7_75t_L g18003 ( 
.A(n_17502),
.Y(n_18003)
);

INVx2_ASAP7_75t_L g18004 ( 
.A(n_17421),
.Y(n_18004)
);

NAND2xp5_ASAP7_75t_L g18005 ( 
.A(n_17372),
.B(n_11184),
.Y(n_18005)
);

NOR2x1p5_ASAP7_75t_L g18006 ( 
.A(n_17546),
.B(n_9174),
.Y(n_18006)
);

INVx1_ASAP7_75t_L g18007 ( 
.A(n_17730),
.Y(n_18007)
);

NAND2xp5_ASAP7_75t_L g18008 ( 
.A(n_17574),
.B(n_11184),
.Y(n_18008)
);

AND2x2_ASAP7_75t_L g18009 ( 
.A(n_17720),
.B(n_17556),
.Y(n_18009)
);

INVx1_ASAP7_75t_L g18010 ( 
.A(n_17727),
.Y(n_18010)
);

INVx2_ASAP7_75t_L g18011 ( 
.A(n_17814),
.Y(n_18011)
);

INVx1_ASAP7_75t_L g18012 ( 
.A(n_17331),
.Y(n_18012)
);

AND2x2_ASAP7_75t_L g18013 ( 
.A(n_17459),
.B(n_11433),
.Y(n_18013)
);

NAND2xp5_ASAP7_75t_L g18014 ( 
.A(n_17601),
.B(n_17392),
.Y(n_18014)
);

AND2x2_ASAP7_75t_L g18015 ( 
.A(n_17466),
.B(n_11433),
.Y(n_18015)
);

INVx2_ASAP7_75t_L g18016 ( 
.A(n_17383),
.Y(n_18016)
);

INVx1_ASAP7_75t_L g18017 ( 
.A(n_17306),
.Y(n_18017)
);

AND2x2_ASAP7_75t_L g18018 ( 
.A(n_17444),
.B(n_17612),
.Y(n_18018)
);

AND2x2_ASAP7_75t_L g18019 ( 
.A(n_17411),
.B(n_11433),
.Y(n_18019)
);

AND2x2_ASAP7_75t_L g18020 ( 
.A(n_17590),
.B(n_11433),
.Y(n_18020)
);

AND2x2_ASAP7_75t_L g18021 ( 
.A(n_17559),
.B(n_11433),
.Y(n_18021)
);

INVx1_ASAP7_75t_L g18022 ( 
.A(n_17307),
.Y(n_18022)
);

AND2x2_ASAP7_75t_L g18023 ( 
.A(n_17563),
.B(n_11433),
.Y(n_18023)
);

NAND2xp5_ASAP7_75t_L g18024 ( 
.A(n_17455),
.B(n_17333),
.Y(n_18024)
);

OR2x2_ASAP7_75t_L g18025 ( 
.A(n_17329),
.B(n_10754),
.Y(n_18025)
);

INVx2_ASAP7_75t_L g18026 ( 
.A(n_17807),
.Y(n_18026)
);

AND2x2_ASAP7_75t_L g18027 ( 
.A(n_17543),
.B(n_17460),
.Y(n_18027)
);

AND2x2_ASAP7_75t_L g18028 ( 
.A(n_17565),
.B(n_10754),
.Y(n_18028)
);

INVx1_ASAP7_75t_L g18029 ( 
.A(n_17318),
.Y(n_18029)
);

NAND2xp5_ASAP7_75t_SL g18030 ( 
.A(n_17431),
.B(n_10036),
.Y(n_18030)
);

INVx2_ASAP7_75t_SL g18031 ( 
.A(n_17431),
.Y(n_18031)
);

NAND2xp5_ASAP7_75t_L g18032 ( 
.A(n_17332),
.B(n_11184),
.Y(n_18032)
);

HB1xp67_ASAP7_75t_L g18033 ( 
.A(n_17645),
.Y(n_18033)
);

INVx2_ASAP7_75t_L g18034 ( 
.A(n_17807),
.Y(n_18034)
);

NAND2x1p5_ASAP7_75t_L g18035 ( 
.A(n_17596),
.B(n_10169),
.Y(n_18035)
);

INVx2_ASAP7_75t_L g18036 ( 
.A(n_17487),
.Y(n_18036)
);

AND2x2_ASAP7_75t_L g18037 ( 
.A(n_17494),
.B(n_17495),
.Y(n_18037)
);

AND2x2_ASAP7_75t_L g18038 ( 
.A(n_17657),
.B(n_10754),
.Y(n_18038)
);

AND2x2_ASAP7_75t_L g18039 ( 
.A(n_17496),
.B(n_10782),
.Y(n_18039)
);

AND2x2_ASAP7_75t_L g18040 ( 
.A(n_17456),
.B(n_10782),
.Y(n_18040)
);

INVx2_ASAP7_75t_L g18041 ( 
.A(n_17516),
.Y(n_18041)
);

INVx1_ASAP7_75t_L g18042 ( 
.A(n_17320),
.Y(n_18042)
);

AND2x4_ASAP7_75t_L g18043 ( 
.A(n_17570),
.B(n_9461),
.Y(n_18043)
);

OR2x2_ASAP7_75t_L g18044 ( 
.A(n_17412),
.B(n_10782),
.Y(n_18044)
);

AND2x2_ASAP7_75t_SL g18045 ( 
.A(n_17831),
.B(n_9775),
.Y(n_18045)
);

INVx1_ASAP7_75t_L g18046 ( 
.A(n_17475),
.Y(n_18046)
);

INVx1_ASAP7_75t_L g18047 ( 
.A(n_17475),
.Y(n_18047)
);

NAND2x1_ASAP7_75t_L g18048 ( 
.A(n_17527),
.B(n_17561),
.Y(n_18048)
);

INVx1_ASAP7_75t_L g18049 ( 
.A(n_17342),
.Y(n_18049)
);

INVx2_ASAP7_75t_L g18050 ( 
.A(n_17767),
.Y(n_18050)
);

NAND2xp5_ASAP7_75t_SL g18051 ( 
.A(n_17458),
.B(n_10036),
.Y(n_18051)
);

INVx2_ASAP7_75t_L g18052 ( 
.A(n_17767),
.Y(n_18052)
);

INVx2_ASAP7_75t_L g18053 ( 
.A(n_17778),
.Y(n_18053)
);

OR2x2_ASAP7_75t_L g18054 ( 
.A(n_17348),
.B(n_17350),
.Y(n_18054)
);

INVx2_ASAP7_75t_L g18055 ( 
.A(n_17778),
.Y(n_18055)
);

NAND2xp5_ASAP7_75t_L g18056 ( 
.A(n_17480),
.B(n_11184),
.Y(n_18056)
);

INVx2_ASAP7_75t_L g18057 ( 
.A(n_17672),
.Y(n_18057)
);

INVx2_ASAP7_75t_SL g18058 ( 
.A(n_17848),
.Y(n_18058)
);

NAND2xp5_ASAP7_75t_SL g18059 ( 
.A(n_17447),
.B(n_10036),
.Y(n_18059)
);

INVx2_ASAP7_75t_L g18060 ( 
.A(n_17681),
.Y(n_18060)
);

OR2x2_ASAP7_75t_L g18061 ( 
.A(n_17613),
.B(n_10782),
.Y(n_18061)
);

INVx1_ASAP7_75t_L g18062 ( 
.A(n_17483),
.Y(n_18062)
);

INVx1_ASAP7_75t_L g18063 ( 
.A(n_17483),
.Y(n_18063)
);

HB1xp67_ASAP7_75t_L g18064 ( 
.A(n_17533),
.Y(n_18064)
);

NAND2xp5_ASAP7_75t_L g18065 ( 
.A(n_17534),
.B(n_11184),
.Y(n_18065)
);

AND2x2_ASAP7_75t_L g18066 ( 
.A(n_17635),
.B(n_10782),
.Y(n_18066)
);

AND2x2_ASAP7_75t_L g18067 ( 
.A(n_17493),
.B(n_10782),
.Y(n_18067)
);

INVx1_ASAP7_75t_L g18068 ( 
.A(n_17533),
.Y(n_18068)
);

INVxp67_ASAP7_75t_L g18069 ( 
.A(n_17351),
.Y(n_18069)
);

AND2x2_ASAP7_75t_L g18070 ( 
.A(n_17577),
.B(n_10782),
.Y(n_18070)
);

OR2x2_ASAP7_75t_L g18071 ( 
.A(n_17877),
.B(n_17810),
.Y(n_18071)
);

INVx1_ASAP7_75t_L g18072 ( 
.A(n_17605),
.Y(n_18072)
);

INVx1_ASAP7_75t_L g18073 ( 
.A(n_17605),
.Y(n_18073)
);

INVx2_ASAP7_75t_L g18074 ( 
.A(n_17651),
.Y(n_18074)
);

INVx2_ASAP7_75t_L g18075 ( 
.A(n_17693),
.Y(n_18075)
);

AND2x2_ASAP7_75t_L g18076 ( 
.A(n_17580),
.B(n_10782),
.Y(n_18076)
);

INVx1_ASAP7_75t_L g18077 ( 
.A(n_17303),
.Y(n_18077)
);

AND2x2_ASAP7_75t_L g18078 ( 
.A(n_17530),
.B(n_11148),
.Y(n_18078)
);

OR2x2_ASAP7_75t_L g18079 ( 
.A(n_17394),
.B(n_11284),
.Y(n_18079)
);

AND2x2_ASAP7_75t_L g18080 ( 
.A(n_17442),
.B(n_11148),
.Y(n_18080)
);

INVx1_ASAP7_75t_L g18081 ( 
.A(n_17305),
.Y(n_18081)
);

NAND2xp5_ASAP7_75t_L g18082 ( 
.A(n_17572),
.B(n_11034),
.Y(n_18082)
);

INVx1_ASAP7_75t_L g18083 ( 
.A(n_17626),
.Y(n_18083)
);

INVx2_ASAP7_75t_L g18084 ( 
.A(n_17698),
.Y(n_18084)
);

NAND2xp5_ASAP7_75t_L g18085 ( 
.A(n_17581),
.B(n_11034),
.Y(n_18085)
);

AND2x2_ASAP7_75t_L g18086 ( 
.A(n_17523),
.B(n_11148),
.Y(n_18086)
);

INVx1_ASAP7_75t_L g18087 ( 
.A(n_17748),
.Y(n_18087)
);

INVx2_ASAP7_75t_L g18088 ( 
.A(n_17699),
.Y(n_18088)
);

NAND2xp5_ASAP7_75t_L g18089 ( 
.A(n_17391),
.B(n_11034),
.Y(n_18089)
);

INVxp67_ASAP7_75t_L g18090 ( 
.A(n_17360),
.Y(n_18090)
);

INVxp67_ASAP7_75t_L g18091 ( 
.A(n_17648),
.Y(n_18091)
);

INVx2_ASAP7_75t_SL g18092 ( 
.A(n_17591),
.Y(n_18092)
);

AND2x2_ASAP7_75t_L g18093 ( 
.A(n_17531),
.B(n_11148),
.Y(n_18093)
);

INVx1_ASAP7_75t_L g18094 ( 
.A(n_17680),
.Y(n_18094)
);

INVx1_ASAP7_75t_L g18095 ( 
.A(n_17680),
.Y(n_18095)
);

AND2x2_ASAP7_75t_L g18096 ( 
.A(n_17463),
.B(n_11148),
.Y(n_18096)
);

INVx2_ASAP7_75t_L g18097 ( 
.A(n_17700),
.Y(n_18097)
);

NOR2xp33_ASAP7_75t_L g18098 ( 
.A(n_17510),
.B(n_10159),
.Y(n_18098)
);

AND2x2_ASAP7_75t_L g18099 ( 
.A(n_17471),
.B(n_11148),
.Y(n_18099)
);

NAND2xp5_ASAP7_75t_L g18100 ( 
.A(n_17437),
.B(n_11034),
.Y(n_18100)
);

AND2x2_ASAP7_75t_L g18101 ( 
.A(n_17529),
.B(n_11148),
.Y(n_18101)
);

HB1xp67_ASAP7_75t_L g18102 ( 
.A(n_17732),
.Y(n_18102)
);

OR2x6_ASAP7_75t_L g18103 ( 
.A(n_17622),
.B(n_10027),
.Y(n_18103)
);

INVx2_ASAP7_75t_SL g18104 ( 
.A(n_17555),
.Y(n_18104)
);

AND2x4_ASAP7_75t_L g18105 ( 
.A(n_17521),
.B(n_9461),
.Y(n_18105)
);

INVx1_ASAP7_75t_L g18106 ( 
.A(n_17813),
.Y(n_18106)
);

OR2x6_ASAP7_75t_L g18107 ( 
.A(n_17422),
.B(n_10027),
.Y(n_18107)
);

INVx1_ASAP7_75t_L g18108 ( 
.A(n_17296),
.Y(n_18108)
);

INVx1_ASAP7_75t_L g18109 ( 
.A(n_17302),
.Y(n_18109)
);

AND2x2_ASAP7_75t_L g18110 ( 
.A(n_17660),
.B(n_17694),
.Y(n_18110)
);

OR2x2_ASAP7_75t_L g18111 ( 
.A(n_17441),
.B(n_11284),
.Y(n_18111)
);

OR2x2_ASAP7_75t_L g18112 ( 
.A(n_17378),
.B(n_11284),
.Y(n_18112)
);

OR2x2_ASAP7_75t_L g18113 ( 
.A(n_17594),
.B(n_11284),
.Y(n_18113)
);

AND2x2_ASAP7_75t_L g18114 ( 
.A(n_17889),
.B(n_11148),
.Y(n_18114)
);

OR2x2_ASAP7_75t_L g18115 ( 
.A(n_17604),
.B(n_11284),
.Y(n_18115)
);

NAND2xp5_ASAP7_75t_L g18116 ( 
.A(n_17773),
.B(n_11034),
.Y(n_18116)
);

INVx2_ASAP7_75t_L g18117 ( 
.A(n_17702),
.Y(n_18117)
);

BUFx2_ASAP7_75t_L g18118 ( 
.A(n_17489),
.Y(n_18118)
);

NAND2xp5_ASAP7_75t_L g18119 ( 
.A(n_17795),
.B(n_11034),
.Y(n_18119)
);

AND2x2_ASAP7_75t_L g18120 ( 
.A(n_17679),
.B(n_10084),
.Y(n_18120)
);

AND2x4_ASAP7_75t_L g18121 ( 
.A(n_17726),
.B(n_9472),
.Y(n_18121)
);

AND3x2_ASAP7_75t_L g18122 ( 
.A(n_17837),
.B(n_10173),
.C(n_10172),
.Y(n_18122)
);

NAND2xp5_ASAP7_75t_L g18123 ( 
.A(n_17670),
.B(n_11034),
.Y(n_18123)
);

NOR3xp33_ASAP7_75t_L g18124 ( 
.A(n_17659),
.B(n_10795),
.C(n_10741),
.Y(n_18124)
);

AND2x2_ASAP7_75t_L g18125 ( 
.A(n_17802),
.B(n_10084),
.Y(n_18125)
);

INVx2_ASAP7_75t_SL g18126 ( 
.A(n_17308),
.Y(n_18126)
);

AND2x2_ASAP7_75t_L g18127 ( 
.A(n_17740),
.B(n_10084),
.Y(n_18127)
);

AND2x2_ASAP7_75t_L g18128 ( 
.A(n_17579),
.B(n_10084),
.Y(n_18128)
);

NAND2xp5_ASAP7_75t_L g18129 ( 
.A(n_17686),
.B(n_11034),
.Y(n_18129)
);

INVx1_ASAP7_75t_L g18130 ( 
.A(n_17704),
.Y(n_18130)
);

INVx1_ASAP7_75t_L g18131 ( 
.A(n_17793),
.Y(n_18131)
);

INVxp67_ASAP7_75t_L g18132 ( 
.A(n_17340),
.Y(n_18132)
);

BUFx2_ASAP7_75t_L g18133 ( 
.A(n_17860),
.Y(n_18133)
);

AND2x2_ASAP7_75t_L g18134 ( 
.A(n_17526),
.B(n_10084),
.Y(n_18134)
);

NAND2xp5_ASAP7_75t_L g18135 ( 
.A(n_17733),
.B(n_10173),
.Y(n_18135)
);

AND2x2_ASAP7_75t_L g18136 ( 
.A(n_17606),
.B(n_10102),
.Y(n_18136)
);

NAND2xp5_ASAP7_75t_L g18137 ( 
.A(n_17427),
.B(n_10173),
.Y(n_18137)
);

NAND2xp5_ASAP7_75t_L g18138 ( 
.A(n_17435),
.B(n_10190),
.Y(n_18138)
);

INVx1_ASAP7_75t_L g18139 ( 
.A(n_17799),
.Y(n_18139)
);

INVx2_ASAP7_75t_L g18140 ( 
.A(n_17862),
.Y(n_18140)
);

INVx2_ASAP7_75t_L g18141 ( 
.A(n_17874),
.Y(n_18141)
);

NAND2x1p5_ASAP7_75t_L g18142 ( 
.A(n_17706),
.B(n_17453),
.Y(n_18142)
);

AND2x2_ASAP7_75t_L g18143 ( 
.A(n_17576),
.B(n_10102),
.Y(n_18143)
);

INVx1_ASAP7_75t_L g18144 ( 
.A(n_17852),
.Y(n_18144)
);

NAND2xp5_ASAP7_75t_L g18145 ( 
.A(n_17443),
.B(n_10190),
.Y(n_18145)
);

INVx1_ASAP7_75t_L g18146 ( 
.A(n_17852),
.Y(n_18146)
);

INVxp67_ASAP7_75t_SL g18147 ( 
.A(n_17518),
.Y(n_18147)
);

AND2x2_ASAP7_75t_L g18148 ( 
.A(n_17384),
.B(n_10102),
.Y(n_18148)
);

AND2x2_ASAP7_75t_L g18149 ( 
.A(n_17637),
.B(n_10102),
.Y(n_18149)
);

INVx1_ASAP7_75t_L g18150 ( 
.A(n_17446),
.Y(n_18150)
);

AND3x2_ASAP7_75t_L g18151 ( 
.A(n_17665),
.B(n_17806),
.C(n_17654),
.Y(n_18151)
);

NAND2xp5_ASAP7_75t_L g18152 ( 
.A(n_17470),
.B(n_10190),
.Y(n_18152)
);

INVx5_ASAP7_75t_L g18153 ( 
.A(n_17640),
.Y(n_18153)
);

NAND2xp5_ASAP7_75t_L g18154 ( 
.A(n_17712),
.B(n_10362),
.Y(n_18154)
);

INVx2_ASAP7_75t_L g18155 ( 
.A(n_17292),
.Y(n_18155)
);

OR2x2_ASAP7_75t_L g18156 ( 
.A(n_17315),
.B(n_11284),
.Y(n_18156)
);

INVx1_ASAP7_75t_L g18157 ( 
.A(n_17375),
.Y(n_18157)
);

INVx1_ASAP7_75t_L g18158 ( 
.A(n_17598),
.Y(n_18158)
);

INVx1_ASAP7_75t_L g18159 ( 
.A(n_17515),
.Y(n_18159)
);

NAND2x1p5_ASAP7_75t_L g18160 ( 
.A(n_17499),
.B(n_10169),
.Y(n_18160)
);

AND2x2_ASAP7_75t_L g18161 ( 
.A(n_17879),
.B(n_10102),
.Y(n_18161)
);

INVx1_ASAP7_75t_L g18162 ( 
.A(n_17830),
.Y(n_18162)
);

AND2x2_ASAP7_75t_L g18163 ( 
.A(n_17666),
.B(n_17661),
.Y(n_18163)
);

INVx1_ASAP7_75t_L g18164 ( 
.A(n_17794),
.Y(n_18164)
);

INVx2_ASAP7_75t_L g18165 ( 
.A(n_17433),
.Y(n_18165)
);

INVx2_ASAP7_75t_L g18166 ( 
.A(n_17818),
.Y(n_18166)
);

AND2x2_ASAP7_75t_L g18167 ( 
.A(n_17688),
.B(n_10102),
.Y(n_18167)
);

INVx2_ASAP7_75t_L g18168 ( 
.A(n_17833),
.Y(n_18168)
);

AND2x2_ASAP7_75t_L g18169 ( 
.A(n_17820),
.B(n_10102),
.Y(n_18169)
);

AND2x2_ASAP7_75t_L g18170 ( 
.A(n_17620),
.B(n_10102),
.Y(n_18170)
);

INVx1_ASAP7_75t_L g18171 ( 
.A(n_17537),
.Y(n_18171)
);

INVx3_ASAP7_75t_L g18172 ( 
.A(n_17617),
.Y(n_18172)
);

OR2x2_ASAP7_75t_L g18173 ( 
.A(n_17343),
.B(n_11284),
.Y(n_18173)
);

INVx1_ASAP7_75t_L g18174 ( 
.A(n_17539),
.Y(n_18174)
);

INVx1_ASAP7_75t_L g18175 ( 
.A(n_17550),
.Y(n_18175)
);

AND2x4_ASAP7_75t_L g18176 ( 
.A(n_17788),
.B(n_9472),
.Y(n_18176)
);

INVx1_ASAP7_75t_L g18177 ( 
.A(n_17557),
.Y(n_18177)
);

INVx1_ASAP7_75t_L g18178 ( 
.A(n_17558),
.Y(n_18178)
);

NAND2xp5_ASAP7_75t_L g18179 ( 
.A(n_17328),
.B(n_17562),
.Y(n_18179)
);

NAND2xp5_ASAP7_75t_L g18180 ( 
.A(n_17509),
.B(n_10362),
.Y(n_18180)
);

NAND2xp5_ASAP7_75t_L g18181 ( 
.A(n_17503),
.B(n_10362),
.Y(n_18181)
);

NAND2xp5_ASAP7_75t_SL g18182 ( 
.A(n_17482),
.B(n_10036),
.Y(n_18182)
);

AND2x2_ASAP7_75t_L g18183 ( 
.A(n_17592),
.B(n_10102),
.Y(n_18183)
);

NAND2xp5_ASAP7_75t_L g18184 ( 
.A(n_17522),
.B(n_10362),
.Y(n_18184)
);

AND2x2_ASAP7_75t_L g18185 ( 
.A(n_17805),
.B(n_8253),
.Y(n_18185)
);

OR2x2_ASAP7_75t_L g18186 ( 
.A(n_17789),
.B(n_11284),
.Y(n_18186)
);

AND2x2_ASAP7_75t_L g18187 ( 
.A(n_17816),
.B(n_8253),
.Y(n_18187)
);

INVx2_ASAP7_75t_L g18188 ( 
.A(n_17840),
.Y(n_18188)
);

INVx1_ASAP7_75t_L g18189 ( 
.A(n_17525),
.Y(n_18189)
);

OR2x2_ASAP7_75t_L g18190 ( 
.A(n_17801),
.B(n_11349),
.Y(n_18190)
);

INVx1_ASAP7_75t_L g18191 ( 
.A(n_17589),
.Y(n_18191)
);

INVx1_ASAP7_75t_L g18192 ( 
.A(n_17511),
.Y(n_18192)
);

INVx2_ASAP7_75t_L g18193 ( 
.A(n_17735),
.Y(n_18193)
);

INVx2_ASAP7_75t_L g18194 ( 
.A(n_17593),
.Y(n_18194)
);

OR2x2_ASAP7_75t_L g18195 ( 
.A(n_17513),
.B(n_11349),
.Y(n_18195)
);

NAND2x1p5_ASAP7_75t_L g18196 ( 
.A(n_17575),
.B(n_17588),
.Y(n_18196)
);

NOR2xp33_ASAP7_75t_L g18197 ( 
.A(n_17629),
.B(n_10169),
.Y(n_18197)
);

NAND2xp5_ASAP7_75t_L g18198 ( 
.A(n_17792),
.B(n_10362),
.Y(n_18198)
);

OR2x2_ASAP7_75t_L g18199 ( 
.A(n_17514),
.B(n_11349),
.Y(n_18199)
);

AND2x2_ASAP7_75t_L g18200 ( 
.A(n_17689),
.B(n_8253),
.Y(n_18200)
);

OR2x2_ASAP7_75t_L g18201 ( 
.A(n_17477),
.B(n_11349),
.Y(n_18201)
);

AND2x2_ASAP7_75t_L g18202 ( 
.A(n_17803),
.B(n_8253),
.Y(n_18202)
);

AND2x2_ASAP7_75t_L g18203 ( 
.A(n_17804),
.B(n_8286),
.Y(n_18203)
);

INVx1_ASAP7_75t_L g18204 ( 
.A(n_17478),
.Y(n_18204)
);

NAND2xp5_ASAP7_75t_L g18205 ( 
.A(n_17608),
.B(n_10362),
.Y(n_18205)
);

NAND2xp5_ASAP7_75t_L g18206 ( 
.A(n_17797),
.B(n_10362),
.Y(n_18206)
);

AND2x4_ASAP7_75t_L g18207 ( 
.A(n_17847),
.B(n_9472),
.Y(n_18207)
);

NAND2xp5_ASAP7_75t_L g18208 ( 
.A(n_17481),
.B(n_10362),
.Y(n_18208)
);

AND2x2_ASAP7_75t_L g18209 ( 
.A(n_17850),
.B(n_8286),
.Y(n_18209)
);

INVx1_ASAP7_75t_L g18210 ( 
.A(n_17486),
.Y(n_18210)
);

INVx1_ASAP7_75t_L g18211 ( 
.A(n_17844),
.Y(n_18211)
);

AND2x2_ASAP7_75t_L g18212 ( 
.A(n_17858),
.B(n_8286),
.Y(n_18212)
);

OR2x2_ASAP7_75t_L g18213 ( 
.A(n_17623),
.B(n_11349),
.Y(n_18213)
);

INVx1_ASAP7_75t_L g18214 ( 
.A(n_17650),
.Y(n_18214)
);

INVx3_ASAP7_75t_SL g18215 ( 
.A(n_17863),
.Y(n_18215)
);

INVx2_ASAP7_75t_L g18216 ( 
.A(n_17829),
.Y(n_18216)
);

OAI21xp5_ASAP7_75t_L g18217 ( 
.A1(n_17299),
.A2(n_10774),
.B(n_10771),
.Y(n_18217)
);

NAND2xp5_ASAP7_75t_L g18218 ( 
.A(n_17462),
.B(n_10571),
.Y(n_18218)
);

AND2x2_ASAP7_75t_SL g18219 ( 
.A(n_17313),
.B(n_9775),
.Y(n_18219)
);

INVx2_ASAP7_75t_L g18220 ( 
.A(n_17677),
.Y(n_18220)
);

NAND2x1p5_ASAP7_75t_L g18221 ( 
.A(n_17855),
.B(n_10169),
.Y(n_18221)
);

OR2x2_ASAP7_75t_L g18222 ( 
.A(n_17836),
.B(n_11349),
.Y(n_18222)
);

AND2x2_ASAP7_75t_L g18223 ( 
.A(n_17859),
.B(n_8286),
.Y(n_18223)
);

OR2x2_ASAP7_75t_L g18224 ( 
.A(n_17532),
.B(n_11349),
.Y(n_18224)
);

NOR2xp33_ASAP7_75t_L g18225 ( 
.A(n_17762),
.B(n_10169),
.Y(n_18225)
);

NAND2x1_ASAP7_75t_L g18226 ( 
.A(n_17308),
.B(n_10169),
.Y(n_18226)
);

NAND2xp5_ASAP7_75t_L g18227 ( 
.A(n_17869),
.B(n_10571),
.Y(n_18227)
);

AND2x2_ASAP7_75t_L g18228 ( 
.A(n_17817),
.B(n_8291),
.Y(n_18228)
);

NOR2xp33_ASAP7_75t_L g18229 ( 
.A(n_17656),
.B(n_17878),
.Y(n_18229)
);

OR2x2_ASAP7_75t_L g18230 ( 
.A(n_17536),
.B(n_11349),
.Y(n_18230)
);

NAND2xp5_ASAP7_75t_L g18231 ( 
.A(n_17414),
.B(n_10571),
.Y(n_18231)
);

INVx1_ASAP7_75t_L g18232 ( 
.A(n_17881),
.Y(n_18232)
);

INVx1_ASAP7_75t_L g18233 ( 
.A(n_17683),
.Y(n_18233)
);

AND2x2_ASAP7_75t_L g18234 ( 
.A(n_17880),
.B(n_8291),
.Y(n_18234)
);

AND2x2_ASAP7_75t_L g18235 ( 
.A(n_17842),
.B(n_8291),
.Y(n_18235)
);

OR2x2_ASAP7_75t_L g18236 ( 
.A(n_17413),
.B(n_11354),
.Y(n_18236)
);

NOR2x1_ASAP7_75t_L g18237 ( 
.A(n_17387),
.B(n_10169),
.Y(n_18237)
);

HB1xp67_ASAP7_75t_L g18238 ( 
.A(n_17655),
.Y(n_18238)
);

INVx4_ASAP7_75t_L g18239 ( 
.A(n_17815),
.Y(n_18239)
);

NAND2xp5_ASAP7_75t_L g18240 ( 
.A(n_17417),
.B(n_10571),
.Y(n_18240)
);

INVx2_ASAP7_75t_L g18241 ( 
.A(n_17841),
.Y(n_18241)
);

INVx1_ASAP7_75t_L g18242 ( 
.A(n_17800),
.Y(n_18242)
);

INVx1_ASAP7_75t_L g18243 ( 
.A(n_17419),
.Y(n_18243)
);

AND2x4_ASAP7_75t_L g18244 ( 
.A(n_17632),
.B(n_17625),
.Y(n_18244)
);

NAND2x1_ASAP7_75t_L g18245 ( 
.A(n_17682),
.B(n_10169),
.Y(n_18245)
);

AND2x2_ASAP7_75t_L g18246 ( 
.A(n_17498),
.B(n_8291),
.Y(n_18246)
);

INVx2_ASAP7_75t_L g18247 ( 
.A(n_17457),
.Y(n_18247)
);

OR2x2_ASAP7_75t_L g18248 ( 
.A(n_17627),
.B(n_11354),
.Y(n_18248)
);

AND2x2_ASAP7_75t_L g18249 ( 
.A(n_17501),
.B(n_8363),
.Y(n_18249)
);

OAI21xp5_ASAP7_75t_L g18250 ( 
.A1(n_17304),
.A2(n_10922),
.B(n_10915),
.Y(n_18250)
);

INVx2_ASAP7_75t_SL g18251 ( 
.A(n_17714),
.Y(n_18251)
);

NAND2xp5_ASAP7_75t_L g18252 ( 
.A(n_17420),
.B(n_10571),
.Y(n_18252)
);

INVx1_ASAP7_75t_L g18253 ( 
.A(n_17582),
.Y(n_18253)
);

NAND2xp5_ASAP7_75t_L g18254 ( 
.A(n_17821),
.B(n_10571),
.Y(n_18254)
);

INVx1_ASAP7_75t_L g18255 ( 
.A(n_17630),
.Y(n_18255)
);

AND2x2_ASAP7_75t_L g18256 ( 
.A(n_17552),
.B(n_8363),
.Y(n_18256)
);

AND2x2_ASAP7_75t_L g18257 ( 
.A(n_17646),
.B(n_8363),
.Y(n_18257)
);

NAND2xp5_ASAP7_75t_L g18258 ( 
.A(n_17832),
.B(n_10571),
.Y(n_18258)
);

INVx1_ASAP7_75t_L g18259 ( 
.A(n_17402),
.Y(n_18259)
);

INVx1_ASAP7_75t_L g18260 ( 
.A(n_17822),
.Y(n_18260)
);

OR2x2_ASAP7_75t_L g18261 ( 
.A(n_17835),
.B(n_11354),
.Y(n_18261)
);

AND2x2_ASAP7_75t_L g18262 ( 
.A(n_17314),
.B(n_8363),
.Y(n_18262)
);

NAND5xp2_ASAP7_75t_L g18263 ( 
.A(n_17324),
.B(n_10047),
.C(n_10104),
.D(n_10038),
.E(n_10011),
.Y(n_18263)
);

OR2x2_ASAP7_75t_L g18264 ( 
.A(n_17347),
.B(n_11354),
.Y(n_18264)
);

AND2x2_ASAP7_75t_L g18265 ( 
.A(n_17314),
.B(n_8382),
.Y(n_18265)
);

AND2x2_ASAP7_75t_L g18266 ( 
.A(n_17541),
.B(n_8382),
.Y(n_18266)
);

OR2x2_ASAP7_75t_L g18267 ( 
.A(n_17448),
.B(n_11354),
.Y(n_18267)
);

INVx2_ASAP7_75t_SL g18268 ( 
.A(n_17312),
.Y(n_18268)
);

INVx2_ASAP7_75t_L g18269 ( 
.A(n_17678),
.Y(n_18269)
);

NAND2x1_ASAP7_75t_L g18270 ( 
.A(n_17736),
.B(n_11679),
.Y(n_18270)
);

INVx1_ASAP7_75t_L g18271 ( 
.A(n_17886),
.Y(n_18271)
);

OR2x2_ASAP7_75t_L g18272 ( 
.A(n_17783),
.B(n_11354),
.Y(n_18272)
);

OR2x2_ASAP7_75t_L g18273 ( 
.A(n_17524),
.B(n_11354),
.Y(n_18273)
);

AND2x2_ASAP7_75t_L g18274 ( 
.A(n_17764),
.B(n_8382),
.Y(n_18274)
);

NAND2xp5_ASAP7_75t_SL g18275 ( 
.A(n_17317),
.B(n_10036),
.Y(n_18275)
);

INVx1_ASAP7_75t_L g18276 ( 
.A(n_17472),
.Y(n_18276)
);

AND2x2_ASAP7_75t_L g18277 ( 
.A(n_17766),
.B(n_8382),
.Y(n_18277)
);

INVx2_ASAP7_75t_L g18278 ( 
.A(n_17544),
.Y(n_18278)
);

OR2x2_ASAP7_75t_L g18279 ( 
.A(n_17653),
.B(n_11354),
.Y(n_18279)
);

OR2x2_ASAP7_75t_L g18280 ( 
.A(n_17663),
.B(n_17664),
.Y(n_18280)
);

INVx1_ASAP7_75t_L g18281 ( 
.A(n_17633),
.Y(n_18281)
);

NAND2xp5_ASAP7_75t_SL g18282 ( 
.A(n_17345),
.B(n_10048),
.Y(n_18282)
);

INVx2_ASAP7_75t_SL g18283 ( 
.A(n_17312),
.Y(n_18283)
);

HB1xp67_ASAP7_75t_L g18284 ( 
.A(n_17639),
.Y(n_18284)
);

OR2x2_ASAP7_75t_L g18285 ( 
.A(n_17667),
.B(n_11499),
.Y(n_18285)
);

INVx1_ASAP7_75t_L g18286 ( 
.A(n_17634),
.Y(n_18286)
);

INVx1_ASAP7_75t_SL g18287 ( 
.A(n_17624),
.Y(n_18287)
);

INVx2_ASAP7_75t_SL g18288 ( 
.A(n_17311),
.Y(n_18288)
);

AND2x2_ASAP7_75t_L g18289 ( 
.A(n_17770),
.B(n_8394),
.Y(n_18289)
);

AND2x2_ASAP7_75t_L g18290 ( 
.A(n_17403),
.B(n_8394),
.Y(n_18290)
);

INVx1_ASAP7_75t_L g18291 ( 
.A(n_17641),
.Y(n_18291)
);

OR2x6_ASAP7_75t_L g18292 ( 
.A(n_17449),
.B(n_10027),
.Y(n_18292)
);

NAND2xp5_ASAP7_75t_L g18293 ( 
.A(n_17658),
.B(n_17721),
.Y(n_18293)
);

INVx2_ASAP7_75t_L g18294 ( 
.A(n_17423),
.Y(n_18294)
);

AND2x2_ASAP7_75t_L g18295 ( 
.A(n_17403),
.B(n_8394),
.Y(n_18295)
);

INVx1_ASAP7_75t_SL g18296 ( 
.A(n_17649),
.Y(n_18296)
);

NOR2xp33_ASAP7_75t_L g18297 ( 
.A(n_17819),
.B(n_10741),
.Y(n_18297)
);

INVx2_ASAP7_75t_L g18298 ( 
.A(n_17425),
.Y(n_18298)
);

OR2x2_ASAP7_75t_L g18299 ( 
.A(n_17673),
.B(n_11499),
.Y(n_18299)
);

INVx2_ASAP7_75t_L g18300 ( 
.A(n_17567),
.Y(n_18300)
);

INVx1_ASAP7_75t_L g18301 ( 
.A(n_17691),
.Y(n_18301)
);

INVxp67_ASAP7_75t_L g18302 ( 
.A(n_17400),
.Y(n_18302)
);

NAND2xp5_ASAP7_75t_L g18303 ( 
.A(n_17722),
.B(n_10571),
.Y(n_18303)
);

AND2x4_ASAP7_75t_L g18304 ( 
.A(n_17669),
.B(n_9472),
.Y(n_18304)
);

INVx2_ASAP7_75t_L g18305 ( 
.A(n_17769),
.Y(n_18305)
);

INVx1_ASAP7_75t_L g18306 ( 
.A(n_17675),
.Y(n_18306)
);

AND2x2_ASAP7_75t_L g18307 ( 
.A(n_17548),
.B(n_8394),
.Y(n_18307)
);

AND2x4_ASAP7_75t_L g18308 ( 
.A(n_17614),
.B(n_9472),
.Y(n_18308)
);

AND2x2_ASAP7_75t_L g18309 ( 
.A(n_17586),
.B(n_8443),
.Y(n_18309)
);

NOR2xp33_ASAP7_75t_L g18310 ( 
.A(n_17846),
.B(n_10741),
.Y(n_18310)
);

AND2x4_ASAP7_75t_L g18311 ( 
.A(n_17731),
.B(n_9526),
.Y(n_18311)
);

OR2x2_ASAP7_75t_L g18312 ( 
.A(n_17451),
.B(n_11499),
.Y(n_18312)
);

NAND2xp5_ASAP7_75t_L g18313 ( 
.A(n_17737),
.B(n_10654),
.Y(n_18313)
);

INVx1_ASAP7_75t_L g18314 ( 
.A(n_17768),
.Y(n_18314)
);

NAND2xp5_ASAP7_75t_L g18315 ( 
.A(n_17739),
.B(n_10654),
.Y(n_18315)
);

AND2x4_ASAP7_75t_L g18316 ( 
.A(n_17751),
.B(n_9526),
.Y(n_18316)
);

INVx1_ASAP7_75t_L g18317 ( 
.A(n_17729),
.Y(n_18317)
);

INVx1_ASAP7_75t_L g18318 ( 
.A(n_17755),
.Y(n_18318)
);

AND2x2_ASAP7_75t_L g18319 ( 
.A(n_17583),
.B(n_8443),
.Y(n_18319)
);

NAND2xp5_ASAP7_75t_L g18320 ( 
.A(n_17756),
.B(n_10654),
.Y(n_18320)
);

INVx2_ASAP7_75t_L g18321 ( 
.A(n_17508),
.Y(n_18321)
);

NAND2xp5_ASAP7_75t_L g18322 ( 
.A(n_17864),
.B(n_10654),
.Y(n_18322)
);

NAND2xp5_ASAP7_75t_SL g18323 ( 
.A(n_17611),
.B(n_10048),
.Y(n_18323)
);

NAND2xp5_ASAP7_75t_L g18324 ( 
.A(n_17297),
.B(n_10654),
.Y(n_18324)
);

NAND2xp5_ASAP7_75t_L g18325 ( 
.A(n_17872),
.B(n_10654),
.Y(n_18325)
);

OR2x2_ASAP7_75t_L g18326 ( 
.A(n_17757),
.B(n_11499),
.Y(n_18326)
);

INVxp67_ASAP7_75t_L g18327 ( 
.A(n_17750),
.Y(n_18327)
);

AND2x2_ASAP7_75t_L g18328 ( 
.A(n_17743),
.B(n_8443),
.Y(n_18328)
);

OAI21xp5_ASAP7_75t_L g18329 ( 
.A1(n_17326),
.A2(n_10922),
.B(n_10915),
.Y(n_18329)
);

INVx1_ASAP7_75t_L g18330 ( 
.A(n_17772),
.Y(n_18330)
);

OR2x2_ASAP7_75t_L g18331 ( 
.A(n_17809),
.B(n_11499),
.Y(n_18331)
);

INVx1_ASAP7_75t_L g18332 ( 
.A(n_17775),
.Y(n_18332)
);

INVx2_ASAP7_75t_SL g18333 ( 
.A(n_17325),
.Y(n_18333)
);

INVx1_ASAP7_75t_L g18334 ( 
.A(n_17776),
.Y(n_18334)
);

OR2x2_ASAP7_75t_L g18335 ( 
.A(n_17587),
.B(n_11499),
.Y(n_18335)
);

NAND2xp5_ASAP7_75t_L g18336 ( 
.A(n_17784),
.B(n_10654),
.Y(n_18336)
);

INVx1_ASAP7_75t_L g18337 ( 
.A(n_17811),
.Y(n_18337)
);

INVx1_ASAP7_75t_L g18338 ( 
.A(n_17824),
.Y(n_18338)
);

INVx2_ASAP7_75t_L g18339 ( 
.A(n_17467),
.Y(n_18339)
);

INVx1_ASAP7_75t_L g18340 ( 
.A(n_17825),
.Y(n_18340)
);

OAI21xp5_ASAP7_75t_L g18341 ( 
.A1(n_17349),
.A2(n_10922),
.B(n_10915),
.Y(n_18341)
);

INVx1_ASAP7_75t_L g18342 ( 
.A(n_17826),
.Y(n_18342)
);

AND2x2_ASAP7_75t_L g18343 ( 
.A(n_17638),
.B(n_17781),
.Y(n_18343)
);

INVx5_ASAP7_75t_SL g18344 ( 
.A(n_17325),
.Y(n_18344)
);

AND2x2_ASAP7_75t_L g18345 ( 
.A(n_17753),
.B(n_8443),
.Y(n_18345)
);

OR3x2_ASAP7_75t_L g18346 ( 
.A(n_17697),
.B(n_10795),
.C(n_10815),
.Y(n_18346)
);

AND2x2_ASAP7_75t_L g18347 ( 
.A(n_17765),
.B(n_8478),
.Y(n_18347)
);

INVx1_ASAP7_75t_SL g18348 ( 
.A(n_17690),
.Y(n_18348)
);

OR2x2_ASAP7_75t_L g18349 ( 
.A(n_17759),
.B(n_11499),
.Y(n_18349)
);

AND2x2_ASAP7_75t_L g18350 ( 
.A(n_17782),
.B(n_8478),
.Y(n_18350)
);

INVx1_ASAP7_75t_L g18351 ( 
.A(n_17828),
.Y(n_18351)
);

INVx1_ASAP7_75t_L g18352 ( 
.A(n_17834),
.Y(n_18352)
);

OR2x2_ASAP7_75t_L g18353 ( 
.A(n_17761),
.B(n_11499),
.Y(n_18353)
);

INVx1_ASAP7_75t_L g18354 ( 
.A(n_17838),
.Y(n_18354)
);

INVx1_ASAP7_75t_L g18355 ( 
.A(n_17839),
.Y(n_18355)
);

OR2x2_ASAP7_75t_L g18356 ( 
.A(n_17771),
.B(n_11514),
.Y(n_18356)
);

NAND2xp5_ASAP7_75t_L g18357 ( 
.A(n_17849),
.B(n_10654),
.Y(n_18357)
);

AND2x4_ASAP7_75t_L g18358 ( 
.A(n_17615),
.B(n_9526),
.Y(n_18358)
);

INVx2_ASAP7_75t_L g18359 ( 
.A(n_17468),
.Y(n_18359)
);

AND2x2_ASAP7_75t_L g18360 ( 
.A(n_17668),
.B(n_8478),
.Y(n_18360)
);

INVxp67_ASAP7_75t_SL g18361 ( 
.A(n_17610),
.Y(n_18361)
);

INVx2_ASAP7_75t_L g18362 ( 
.A(n_17512),
.Y(n_18362)
);

NOR3x1_ASAP7_75t_L g18363 ( 
.A(n_17780),
.B(n_9174),
.C(n_9008),
.Y(n_18363)
);

NAND2xp5_ASAP7_75t_L g18364 ( 
.A(n_17851),
.B(n_11244),
.Y(n_18364)
);

OR2x2_ASAP7_75t_L g18365 ( 
.A(n_17636),
.B(n_11514),
.Y(n_18365)
);

INVx1_ASAP7_75t_L g18366 ( 
.A(n_17853),
.Y(n_18366)
);

NAND2xp5_ASAP7_75t_L g18367 ( 
.A(n_17861),
.B(n_11247),
.Y(n_18367)
);

AND2x2_ASAP7_75t_L g18368 ( 
.A(n_17718),
.B(n_8478),
.Y(n_18368)
);

NAND2xp5_ASAP7_75t_L g18369 ( 
.A(n_17866),
.B(n_11247),
.Y(n_18369)
);

INVx1_ASAP7_75t_L g18370 ( 
.A(n_17867),
.Y(n_18370)
);

AND2x2_ASAP7_75t_L g18371 ( 
.A(n_17734),
.B(n_17545),
.Y(n_18371)
);

AND2x2_ASAP7_75t_L g18372 ( 
.A(n_17684),
.B(n_9526),
.Y(n_18372)
);

HB1xp67_ASAP7_75t_L g18373 ( 
.A(n_17339),
.Y(n_18373)
);

INVx1_ASAP7_75t_L g18374 ( 
.A(n_17616),
.Y(n_18374)
);

AND2x4_ASAP7_75t_SL g18375 ( 
.A(n_17674),
.B(n_8124),
.Y(n_18375)
);

INVx1_ASAP7_75t_L g18376 ( 
.A(n_17618),
.Y(n_18376)
);

OR2x2_ASAP7_75t_L g18377 ( 
.A(n_17642),
.B(n_11514),
.Y(n_18377)
);

INVx1_ASAP7_75t_L g18378 ( 
.A(n_17602),
.Y(n_18378)
);

AND2x2_ASAP7_75t_L g18379 ( 
.A(n_17796),
.B(n_9526),
.Y(n_18379)
);

AND2x4_ASAP7_75t_L g18380 ( 
.A(n_17692),
.B(n_9529),
.Y(n_18380)
);

AND2x2_ASAP7_75t_L g18381 ( 
.A(n_17796),
.B(n_9529),
.Y(n_18381)
);

AND2x2_ASAP7_75t_L g18382 ( 
.A(n_17823),
.B(n_9529),
.Y(n_18382)
);

INVx1_ASAP7_75t_L g18383 ( 
.A(n_17888),
.Y(n_18383)
);

NAND2x1p5_ASAP7_75t_L g18384 ( 
.A(n_17695),
.B(n_9587),
.Y(n_18384)
);

AND2x2_ASAP7_75t_L g18385 ( 
.A(n_17440),
.B(n_9529),
.Y(n_18385)
);

NAND2xp5_ASAP7_75t_L g18386 ( 
.A(n_17843),
.B(n_17707),
.Y(n_18386)
);

AND2x2_ASAP7_75t_L g18387 ( 
.A(n_17599),
.B(n_9529),
.Y(n_18387)
);

AND2x2_ASAP7_75t_L g18388 ( 
.A(n_17674),
.B(n_9529),
.Y(n_18388)
);

NAND2xp5_ASAP7_75t_L g18389 ( 
.A(n_17708),
.B(n_17710),
.Y(n_18389)
);

CKINVDCx16_ASAP7_75t_R g18390 ( 
.A(n_17711),
.Y(n_18390)
);

OR2x2_ASAP7_75t_L g18391 ( 
.A(n_17416),
.B(n_11514),
.Y(n_18391)
);

OR2x2_ASAP7_75t_L g18392 ( 
.A(n_17715),
.B(n_11514),
.Y(n_18392)
);

OR2x2_ASAP7_75t_L g18393 ( 
.A(n_17676),
.B(n_11514),
.Y(n_18393)
);

AND2x2_ASAP7_75t_L g18394 ( 
.A(n_17485),
.B(n_9550),
.Y(n_18394)
);

AND2x2_ASAP7_75t_L g18395 ( 
.A(n_17685),
.B(n_9550),
.Y(n_18395)
);

INVx2_ASAP7_75t_L g18396 ( 
.A(n_17619),
.Y(n_18396)
);

INVx1_ASAP7_75t_L g18397 ( 
.A(n_17890),
.Y(n_18397)
);

AND2x2_ASAP7_75t_L g18398 ( 
.A(n_17696),
.B(n_9550),
.Y(n_18398)
);

INVx3_ASAP7_75t_SL g18399 ( 
.A(n_17741),
.Y(n_18399)
);

NAND2xp5_ASAP7_75t_SL g18400 ( 
.A(n_17569),
.B(n_10048),
.Y(n_18400)
);

INVx2_ASAP7_75t_L g18401 ( 
.A(n_17798),
.Y(n_18401)
);

NOR2xp33_ASAP7_75t_L g18402 ( 
.A(n_17744),
.B(n_10795),
.Y(n_18402)
);

INVx1_ASAP7_75t_L g18403 ( 
.A(n_17882),
.Y(n_18403)
);

OR2x2_ASAP7_75t_L g18404 ( 
.A(n_17745),
.B(n_11514),
.Y(n_18404)
);

INVx1_ASAP7_75t_L g18405 ( 
.A(n_17885),
.Y(n_18405)
);

AND2x2_ASAP7_75t_L g18406 ( 
.A(n_17705),
.B(n_9550),
.Y(n_18406)
);

OR2x2_ASAP7_75t_L g18407 ( 
.A(n_17785),
.B(n_11514),
.Y(n_18407)
);

NAND2xp5_ASAP7_75t_L g18408 ( 
.A(n_17752),
.B(n_11256),
.Y(n_18408)
);

INVx1_ASAP7_75t_L g18409 ( 
.A(n_17717),
.Y(n_18409)
);

AOI21xp5_ASAP7_75t_L g18410 ( 
.A1(n_17445),
.A2(n_11766),
.B(n_11698),
.Y(n_18410)
);

INVx2_ASAP7_75t_L g18411 ( 
.A(n_17607),
.Y(n_18411)
);

AND2x2_ASAP7_75t_L g18412 ( 
.A(n_17713),
.B(n_9550),
.Y(n_18412)
);

INVx1_ASAP7_75t_L g18413 ( 
.A(n_17719),
.Y(n_18413)
);

AND2x4_ASAP7_75t_L g18414 ( 
.A(n_17723),
.B(n_9550),
.Y(n_18414)
);

AND2x2_ASAP7_75t_L g18415 ( 
.A(n_17747),
.B(n_9442),
.Y(n_18415)
);

NAND2xp5_ASAP7_75t_L g18416 ( 
.A(n_17724),
.B(n_11256),
.Y(n_18416)
);

NAND2xp5_ASAP7_75t_L g18417 ( 
.A(n_17728),
.B(n_11283),
.Y(n_18417)
);

INVx1_ASAP7_75t_L g18418 ( 
.A(n_17868),
.Y(n_18418)
);

AND2x2_ASAP7_75t_L g18419 ( 
.A(n_17876),
.B(n_9442),
.Y(n_18419)
);

AND2x4_ASAP7_75t_L g18420 ( 
.A(n_17871),
.B(n_9442),
.Y(n_18420)
);

INVx1_ASAP7_75t_L g18421 ( 
.A(n_17628),
.Y(n_18421)
);

INVx1_ASAP7_75t_L g18422 ( 
.A(n_17566),
.Y(n_18422)
);

AND2x2_ASAP7_75t_L g18423 ( 
.A(n_17519),
.B(n_9442),
.Y(n_18423)
);

OR2x2_ASAP7_75t_L g18424 ( 
.A(n_17465),
.B(n_11522),
.Y(n_18424)
);

INVx1_ASAP7_75t_L g18425 ( 
.A(n_17507),
.Y(n_18425)
);

INVx2_ASAP7_75t_L g18426 ( 
.A(n_17609),
.Y(n_18426)
);

AND2x2_ASAP7_75t_L g18427 ( 
.A(n_17873),
.B(n_9442),
.Y(n_18427)
);

INVx1_ASAP7_75t_L g18428 ( 
.A(n_17845),
.Y(n_18428)
);

NAND2xp5_ASAP7_75t_L g18429 ( 
.A(n_17777),
.B(n_11283),
.Y(n_18429)
);

NAND2xp5_ASAP7_75t_L g18430 ( 
.A(n_17856),
.B(n_11286),
.Y(n_18430)
);

AND2x2_ASAP7_75t_L g18431 ( 
.A(n_17873),
.B(n_9442),
.Y(n_18431)
);

NAND2xp5_ASAP7_75t_L g18432 ( 
.A(n_17401),
.B(n_11286),
.Y(n_18432)
);

AND2x2_ASAP7_75t_L g18433 ( 
.A(n_17528),
.B(n_9442),
.Y(n_18433)
);

INVx1_ASAP7_75t_L g18434 ( 
.A(n_17701),
.Y(n_18434)
);

NAND2xp5_ASAP7_75t_L g18435 ( 
.A(n_17373),
.B(n_11289),
.Y(n_18435)
);

AND2x2_ASAP7_75t_L g18436 ( 
.A(n_17415),
.B(n_9442),
.Y(n_18436)
);

INVx1_ASAP7_75t_L g18437 ( 
.A(n_17870),
.Y(n_18437)
);

INVx1_ASAP7_75t_L g18438 ( 
.A(n_17671),
.Y(n_18438)
);

NAND2xp5_ASAP7_75t_L g18439 ( 
.A(n_17887),
.B(n_11289),
.Y(n_18439)
);

INVx1_ASAP7_75t_L g18440 ( 
.A(n_17687),
.Y(n_18440)
);

NAND2xp5_ASAP7_75t_L g18441 ( 
.A(n_17316),
.B(n_17490),
.Y(n_18441)
);

HB1xp67_ASAP7_75t_L g18442 ( 
.A(n_17389),
.Y(n_18442)
);

NAND2xp5_ASAP7_75t_L g18443 ( 
.A(n_17857),
.B(n_11297),
.Y(n_18443)
);

INVx3_ASAP7_75t_SL g18444 ( 
.A(n_17883),
.Y(n_18444)
);

BUFx3_ASAP7_75t_L g18445 ( 
.A(n_18048),
.Y(n_18445)
);

NAND2xp5_ASAP7_75t_L g18446 ( 
.A(n_17978),
.B(n_17914),
.Y(n_18446)
);

AND2x4_ASAP7_75t_SL g18447 ( 
.A(n_18009),
.B(n_17327),
.Y(n_18447)
);

INVxp67_ASAP7_75t_SL g18448 ( 
.A(n_17964),
.Y(n_18448)
);

AO22x1_ASAP7_75t_L g18449 ( 
.A1(n_18147),
.A2(n_17631),
.B1(n_17716),
.B2(n_17738),
.Y(n_18449)
);

INVx1_ASAP7_75t_L g18450 ( 
.A(n_18238),
.Y(n_18450)
);

NAND2xp5_ASAP7_75t_L g18451 ( 
.A(n_18215),
.B(n_17397),
.Y(n_18451)
);

AND2x4_ASAP7_75t_L g18452 ( 
.A(n_17947),
.B(n_18018),
.Y(n_18452)
);

HB1xp67_ASAP7_75t_L g18453 ( 
.A(n_18373),
.Y(n_18453)
);

INVx1_ASAP7_75t_L g18454 ( 
.A(n_18284),
.Y(n_18454)
);

OR2x2_ASAP7_75t_L g18455 ( 
.A(n_18071),
.B(n_17725),
.Y(n_18455)
);

INVx1_ASAP7_75t_L g18456 ( 
.A(n_18033),
.Y(n_18456)
);

NAND2xp5_ASAP7_75t_L g18457 ( 
.A(n_17919),
.B(n_17584),
.Y(n_18457)
);

INVx1_ASAP7_75t_L g18458 ( 
.A(n_17911),
.Y(n_18458)
);

INVx1_ASAP7_75t_L g18459 ( 
.A(n_18247),
.Y(n_18459)
);

INVx1_ASAP7_75t_L g18460 ( 
.A(n_18278),
.Y(n_18460)
);

NAND2xp5_ASAP7_75t_L g18461 ( 
.A(n_18011),
.B(n_17388),
.Y(n_18461)
);

AND2x2_ASAP7_75t_L g18462 ( 
.A(n_17985),
.B(n_18110),
.Y(n_18462)
);

OAI31xp33_ASAP7_75t_L g18463 ( 
.A1(n_18442),
.A2(n_17643),
.A3(n_17571),
.B(n_17547),
.Y(n_18463)
);

NAND2xp5_ASAP7_75t_L g18464 ( 
.A(n_17923),
.B(n_17374),
.Y(n_18464)
);

INVx1_ASAP7_75t_L g18465 ( 
.A(n_18339),
.Y(n_18465)
);

AOI22xp33_ASAP7_75t_L g18466 ( 
.A1(n_18282),
.A2(n_17353),
.B1(n_17461),
.B2(n_17742),
.Y(n_18466)
);

INVx1_ASAP7_75t_L g18467 ( 
.A(n_18321),
.Y(n_18467)
);

INVx1_ASAP7_75t_L g18468 ( 
.A(n_18133),
.Y(n_18468)
);

OR2x2_ASAP7_75t_L g18469 ( 
.A(n_17936),
.B(n_17791),
.Y(n_18469)
);

AND2x2_ASAP7_75t_L g18470 ( 
.A(n_17906),
.B(n_17925),
.Y(n_18470)
);

OR2x2_ASAP7_75t_L g18471 ( 
.A(n_17943),
.B(n_17812),
.Y(n_18471)
);

BUFx2_ASAP7_75t_L g18472 ( 
.A(n_18064),
.Y(n_18472)
);

NAND2xp5_ASAP7_75t_L g18473 ( 
.A(n_17900),
.B(n_17600),
.Y(n_18473)
);

NAND2xp5_ASAP7_75t_L g18474 ( 
.A(n_17907),
.B(n_17540),
.Y(n_18474)
);

INVx1_ASAP7_75t_L g18475 ( 
.A(n_18300),
.Y(n_18475)
);

HB1xp67_ASAP7_75t_L g18476 ( 
.A(n_18245),
.Y(n_18476)
);

AND2x4_ASAP7_75t_L g18477 ( 
.A(n_18153),
.B(n_17790),
.Y(n_18477)
);

OR2x2_ASAP7_75t_L g18478 ( 
.A(n_17909),
.B(n_17652),
.Y(n_18478)
);

AND2x2_ASAP7_75t_L g18479 ( 
.A(n_18027),
.B(n_17854),
.Y(n_18479)
);

AOI21x1_ASAP7_75t_SL g18480 ( 
.A1(n_18441),
.A2(n_17760),
.B(n_17754),
.Y(n_18480)
);

OR2x2_ASAP7_75t_L g18481 ( 
.A(n_17896),
.B(n_17808),
.Y(n_18481)
);

NAND2xp5_ASAP7_75t_L g18482 ( 
.A(n_17981),
.B(n_17520),
.Y(n_18482)
);

AOI221xp5_ASAP7_75t_L g18483 ( 
.A1(n_18132),
.A2(n_17662),
.B1(n_17827),
.B2(n_17746),
.C(n_17779),
.Y(n_18483)
);

OR2x2_ASAP7_75t_L g18484 ( 
.A(n_18024),
.B(n_17644),
.Y(n_18484)
);

OR2x2_ASAP7_75t_L g18485 ( 
.A(n_17954),
.B(n_17875),
.Y(n_18485)
);

BUFx3_ASAP7_75t_L g18486 ( 
.A(n_18196),
.Y(n_18486)
);

NAND2xp5_ASAP7_75t_L g18487 ( 
.A(n_18026),
.B(n_18034),
.Y(n_18487)
);

HB1xp67_ASAP7_75t_L g18488 ( 
.A(n_18153),
.Y(n_18488)
);

INVx2_ASAP7_75t_L g18489 ( 
.A(n_17918),
.Y(n_18489)
);

HB1xp67_ASAP7_75t_L g18490 ( 
.A(n_18428),
.Y(n_18490)
);

OR2x2_ASAP7_75t_L g18491 ( 
.A(n_18390),
.B(n_17758),
.Y(n_18491)
);

INVxp67_ASAP7_75t_L g18492 ( 
.A(n_17904),
.Y(n_18492)
);

NAND2xp5_ASAP7_75t_L g18493 ( 
.A(n_18046),
.B(n_17578),
.Y(n_18493)
);

AND2x2_ASAP7_75t_L g18494 ( 
.A(n_17937),
.B(n_17568),
.Y(n_18494)
);

INVx1_ASAP7_75t_L g18495 ( 
.A(n_18437),
.Y(n_18495)
);

AND2x2_ASAP7_75t_L g18496 ( 
.A(n_17949),
.B(n_17774),
.Y(n_18496)
);

OR2x2_ASAP7_75t_L g18497 ( 
.A(n_17910),
.B(n_17895),
.Y(n_18497)
);

INVx1_ASAP7_75t_L g18498 ( 
.A(n_18118),
.Y(n_18498)
);

AND2x2_ASAP7_75t_L g18499 ( 
.A(n_18037),
.B(n_17865),
.Y(n_18499)
);

INVx2_ASAP7_75t_L g18500 ( 
.A(n_18050),
.Y(n_18500)
);

OAI221xp5_ASAP7_75t_SL g18501 ( 
.A1(n_17929),
.A2(n_18302),
.B1(n_17908),
.B2(n_18090),
.C(n_18091),
.Y(n_18501)
);

INVx1_ASAP7_75t_SL g18502 ( 
.A(n_18399),
.Y(n_18502)
);

OR2x2_ASAP7_75t_L g18503 ( 
.A(n_17926),
.B(n_17787),
.Y(n_18503)
);

INVx1_ASAP7_75t_L g18504 ( 
.A(n_18102),
.Y(n_18504)
);

INVx2_ASAP7_75t_L g18505 ( 
.A(n_18052),
.Y(n_18505)
);

NOR2xp33_ASAP7_75t_L g18506 ( 
.A(n_18239),
.B(n_11297),
.Y(n_18506)
);

NAND2xp5_ASAP7_75t_L g18507 ( 
.A(n_18047),
.B(n_11301),
.Y(n_18507)
);

OR2x2_ASAP7_75t_L g18508 ( 
.A(n_18142),
.B(n_18036),
.Y(n_18508)
);

INVx2_ASAP7_75t_L g18509 ( 
.A(n_18053),
.Y(n_18509)
);

INVx2_ASAP7_75t_L g18510 ( 
.A(n_18055),
.Y(n_18510)
);

INVx1_ASAP7_75t_SL g18511 ( 
.A(n_17973),
.Y(n_18511)
);

INVx1_ASAP7_75t_L g18512 ( 
.A(n_17995),
.Y(n_18512)
);

INVx1_ASAP7_75t_L g18513 ( 
.A(n_18421),
.Y(n_18513)
);

INVx1_ASAP7_75t_L g18514 ( 
.A(n_18422),
.Y(n_18514)
);

AND2x2_ASAP7_75t_L g18515 ( 
.A(n_17976),
.B(n_9442),
.Y(n_18515)
);

OAI31xp67_ASAP7_75t_L g18516 ( 
.A1(n_17960),
.A2(n_9212),
.A3(n_9058),
.B(n_9787),
.Y(n_18516)
);

AND2x2_ASAP7_75t_L g18517 ( 
.A(n_17893),
.B(n_10704),
.Y(n_18517)
);

NOR2x1_ASAP7_75t_L g18518 ( 
.A(n_18062),
.B(n_11766),
.Y(n_18518)
);

INVx1_ASAP7_75t_L g18519 ( 
.A(n_17894),
.Y(n_18519)
);

AND2x2_ASAP7_75t_L g18520 ( 
.A(n_17920),
.B(n_10704),
.Y(n_18520)
);

AND2x2_ASAP7_75t_L g18521 ( 
.A(n_18260),
.B(n_10704),
.Y(n_18521)
);

NAND2x1_ASAP7_75t_L g18522 ( 
.A(n_17968),
.B(n_17959),
.Y(n_18522)
);

OR2x2_ASAP7_75t_L g18523 ( 
.A(n_18041),
.B(n_11301),
.Y(n_18523)
);

NAND2xp5_ASAP7_75t_L g18524 ( 
.A(n_17921),
.B(n_11306),
.Y(n_18524)
);

OR2x2_ASAP7_75t_L g18525 ( 
.A(n_17950),
.B(n_11306),
.Y(n_18525)
);

AND2x2_ASAP7_75t_L g18526 ( 
.A(n_17967),
.B(n_10704),
.Y(n_18526)
);

INVx1_ASAP7_75t_L g18527 ( 
.A(n_17940),
.Y(n_18527)
);

NAND2xp5_ASAP7_75t_L g18528 ( 
.A(n_17924),
.B(n_18229),
.Y(n_18528)
);

INVx1_ASAP7_75t_L g18529 ( 
.A(n_17945),
.Y(n_18529)
);

INVx1_ASAP7_75t_L g18530 ( 
.A(n_17946),
.Y(n_18530)
);

AND2x2_ASAP7_75t_L g18531 ( 
.A(n_17903),
.B(n_17897),
.Y(n_18531)
);

INVx1_ASAP7_75t_L g18532 ( 
.A(n_17971),
.Y(n_18532)
);

AND2x2_ASAP7_75t_L g18533 ( 
.A(n_17915),
.B(n_10704),
.Y(n_18533)
);

HB1xp67_ASAP7_75t_L g18534 ( 
.A(n_18063),
.Y(n_18534)
);

NAND2x1_ASAP7_75t_L g18535 ( 
.A(n_17991),
.B(n_11766),
.Y(n_18535)
);

AND2x2_ASAP7_75t_L g18536 ( 
.A(n_17892),
.B(n_10704),
.Y(n_18536)
);

INVx1_ASAP7_75t_L g18537 ( 
.A(n_18014),
.Y(n_18537)
);

AND2x2_ASAP7_75t_L g18538 ( 
.A(n_17975),
.B(n_10704),
.Y(n_18538)
);

INVx1_ASAP7_75t_L g18539 ( 
.A(n_18087),
.Y(n_18539)
);

AND2x4_ASAP7_75t_L g18540 ( 
.A(n_17934),
.B(n_9186),
.Y(n_18540)
);

NOR2xp33_ASAP7_75t_L g18541 ( 
.A(n_17966),
.B(n_11313),
.Y(n_18541)
);

INVx1_ASAP7_75t_L g18542 ( 
.A(n_18163),
.Y(n_18542)
);

AND2x2_ASAP7_75t_L g18543 ( 
.A(n_18016),
.B(n_10704),
.Y(n_18543)
);

INVx2_ASAP7_75t_L g18544 ( 
.A(n_18035),
.Y(n_18544)
);

INVx1_ASAP7_75t_L g18545 ( 
.A(n_17992),
.Y(n_18545)
);

NAND2xp5_ASAP7_75t_L g18546 ( 
.A(n_17930),
.B(n_11313),
.Y(n_18546)
);

NAND2xp5_ASAP7_75t_L g18547 ( 
.A(n_17931),
.B(n_11328),
.Y(n_18547)
);

INVx1_ASAP7_75t_L g18548 ( 
.A(n_18054),
.Y(n_18548)
);

NOR2xp33_ASAP7_75t_L g18549 ( 
.A(n_18083),
.B(n_11328),
.Y(n_18549)
);

NAND2xp5_ASAP7_75t_L g18550 ( 
.A(n_17933),
.B(n_11331),
.Y(n_18550)
);

INVx2_ASAP7_75t_L g18551 ( 
.A(n_18221),
.Y(n_18551)
);

OR2x2_ASAP7_75t_L g18552 ( 
.A(n_18003),
.B(n_11331),
.Y(n_18552)
);

INVx1_ASAP7_75t_L g18553 ( 
.A(n_17982),
.Y(n_18553)
);

NAND2xp5_ASAP7_75t_L g18554 ( 
.A(n_17935),
.B(n_11332),
.Y(n_18554)
);

NAND2xp5_ASAP7_75t_L g18555 ( 
.A(n_17956),
.B(n_11332),
.Y(n_18555)
);

HB1xp67_ASAP7_75t_L g18556 ( 
.A(n_18068),
.Y(n_18556)
);

NAND2xp5_ASAP7_75t_L g18557 ( 
.A(n_17965),
.B(n_11339),
.Y(n_18557)
);

AOI211xp5_ASAP7_75t_L g18558 ( 
.A1(n_17962),
.A2(n_9211),
.B(n_9386),
.C(n_9159),
.Y(n_18558)
);

INVx1_ASAP7_75t_L g18559 ( 
.A(n_17983),
.Y(n_18559)
);

AND2x2_ASAP7_75t_L g18560 ( 
.A(n_18060),
.B(n_8503),
.Y(n_18560)
);

NAND2xp5_ASAP7_75t_L g18561 ( 
.A(n_17970),
.B(n_11339),
.Y(n_18561)
);

INVx1_ASAP7_75t_SL g18562 ( 
.A(n_18348),
.Y(n_18562)
);

OR2x2_ASAP7_75t_L g18563 ( 
.A(n_18179),
.B(n_11346),
.Y(n_18563)
);

AND2x2_ASAP7_75t_L g18564 ( 
.A(n_17952),
.B(n_8503),
.Y(n_18564)
);

HB1xp67_ASAP7_75t_L g18565 ( 
.A(n_18072),
.Y(n_18565)
);

OAI21xp5_ASAP7_75t_L g18566 ( 
.A1(n_18069),
.A2(n_10699),
.B(n_10748),
.Y(n_18566)
);

INVx1_ASAP7_75t_L g18567 ( 
.A(n_18305),
.Y(n_18567)
);

INVx2_ASAP7_75t_L g18568 ( 
.A(n_18160),
.Y(n_18568)
);

INVx1_ASAP7_75t_L g18569 ( 
.A(n_17993),
.Y(n_18569)
);

OR2x2_ASAP7_75t_L g18570 ( 
.A(n_18194),
.B(n_11346),
.Y(n_18570)
);

INVx1_ASAP7_75t_L g18571 ( 
.A(n_18007),
.Y(n_18571)
);

AND2x2_ASAP7_75t_L g18572 ( 
.A(n_17963),
.B(n_8503),
.Y(n_18572)
);

INVx1_ASAP7_75t_L g18573 ( 
.A(n_18010),
.Y(n_18573)
);

AND2x4_ASAP7_75t_L g18574 ( 
.A(n_18004),
.B(n_9186),
.Y(n_18574)
);

AND2x2_ASAP7_75t_L g18575 ( 
.A(n_17922),
.B(n_8503),
.Y(n_18575)
);

OR2x2_ASAP7_75t_L g18576 ( 
.A(n_18031),
.B(n_11353),
.Y(n_18576)
);

INVx2_ASAP7_75t_L g18577 ( 
.A(n_17974),
.Y(n_18577)
);

NAND2xp5_ASAP7_75t_L g18578 ( 
.A(n_18073),
.B(n_11353),
.Y(n_18578)
);

INVx1_ASAP7_75t_L g18579 ( 
.A(n_17898),
.Y(n_18579)
);

NAND2x2_ASAP7_75t_L g18580 ( 
.A(n_18288),
.B(n_9993),
.Y(n_18580)
);

INVx1_ASAP7_75t_L g18581 ( 
.A(n_17899),
.Y(n_18581)
);

INVxp33_ASAP7_75t_SL g18582 ( 
.A(n_17901),
.Y(n_18582)
);

INVx1_ASAP7_75t_L g18583 ( 
.A(n_18012),
.Y(n_18583)
);

INVxp67_ASAP7_75t_SL g18584 ( 
.A(n_17939),
.Y(n_18584)
);

AND2x2_ASAP7_75t_L g18585 ( 
.A(n_17944),
.B(n_8534),
.Y(n_18585)
);

INVx1_ASAP7_75t_L g18586 ( 
.A(n_17927),
.Y(n_18586)
);

AND2x2_ASAP7_75t_L g18587 ( 
.A(n_18057),
.B(n_8534),
.Y(n_18587)
);

INVx1_ASAP7_75t_L g18588 ( 
.A(n_18094),
.Y(n_18588)
);

NAND2xp5_ASAP7_75t_L g18589 ( 
.A(n_18095),
.B(n_11366),
.Y(n_18589)
);

NOR2x1_ASAP7_75t_L g18590 ( 
.A(n_18144),
.B(n_11366),
.Y(n_18590)
);

AND2x2_ASAP7_75t_L g18591 ( 
.A(n_17984),
.B(n_17980),
.Y(n_18591)
);

AND2x2_ASAP7_75t_L g18592 ( 
.A(n_18166),
.B(n_8534),
.Y(n_18592)
);

OR2x2_ASAP7_75t_L g18593 ( 
.A(n_18293),
.B(n_11375),
.Y(n_18593)
);

INVx2_ASAP7_75t_L g18594 ( 
.A(n_18146),
.Y(n_18594)
);

INVx1_ASAP7_75t_L g18595 ( 
.A(n_18106),
.Y(n_18595)
);

INVxp67_ASAP7_75t_L g18596 ( 
.A(n_17932),
.Y(n_18596)
);

INVx1_ASAP7_75t_L g18597 ( 
.A(n_17917),
.Y(n_18597)
);

AND2x2_ASAP7_75t_L g18598 ( 
.A(n_18074),
.B(n_8534),
.Y(n_18598)
);

OR2x2_ASAP7_75t_L g18599 ( 
.A(n_17961),
.B(n_11375),
.Y(n_18599)
);

INVx2_ASAP7_75t_L g18600 ( 
.A(n_17928),
.Y(n_18600)
);

AND2x2_ASAP7_75t_L g18601 ( 
.A(n_17957),
.B(n_9698),
.Y(n_18601)
);

OR2x6_ASAP7_75t_L g18602 ( 
.A(n_18168),
.B(n_10027),
.Y(n_18602)
);

INVx1_ASAP7_75t_SL g18603 ( 
.A(n_18151),
.Y(n_18603)
);

INVx1_ASAP7_75t_L g18604 ( 
.A(n_18232),
.Y(n_18604)
);

HB1xp67_ASAP7_75t_L g18605 ( 
.A(n_17979),
.Y(n_18605)
);

INVx3_ASAP7_75t_L g18606 ( 
.A(n_18226),
.Y(n_18606)
);

NAND2xp67_ASAP7_75t_L g18607 ( 
.A(n_18155),
.B(n_11277),
.Y(n_18607)
);

AND2x2_ASAP7_75t_L g18608 ( 
.A(n_18220),
.B(n_9698),
.Y(n_18608)
);

INVx1_ASAP7_75t_L g18609 ( 
.A(n_17912),
.Y(n_18609)
);

AOI31xp33_ASAP7_75t_L g18610 ( 
.A1(n_18162),
.A2(n_10038),
.A3(n_10047),
.B(n_10011),
.Y(n_18610)
);

INVx1_ASAP7_75t_L g18611 ( 
.A(n_17938),
.Y(n_18611)
);

INVx1_ASAP7_75t_L g18612 ( 
.A(n_18211),
.Y(n_18612)
);

INVx2_ASAP7_75t_L g18613 ( 
.A(n_18172),
.Y(n_18613)
);

INVx1_ASAP7_75t_L g18614 ( 
.A(n_18361),
.Y(n_18614)
);

AND2x2_ASAP7_75t_L g18615 ( 
.A(n_17955),
.B(n_9698),
.Y(n_18615)
);

INVx1_ASAP7_75t_L g18616 ( 
.A(n_18075),
.Y(n_18616)
);

INVx2_ASAP7_75t_SL g18617 ( 
.A(n_18423),
.Y(n_18617)
);

INVx1_ASAP7_75t_L g18618 ( 
.A(n_18084),
.Y(n_18618)
);

INVxp67_ASAP7_75t_L g18619 ( 
.A(n_18237),
.Y(n_18619)
);

INVx1_ASAP7_75t_L g18620 ( 
.A(n_18088),
.Y(n_18620)
);

INVx1_ASAP7_75t_L g18621 ( 
.A(n_18097),
.Y(n_18621)
);

NAND3xp33_ASAP7_75t_L g18622 ( 
.A(n_17913),
.B(n_10026),
.C(n_10007),
.Y(n_18622)
);

HB1xp67_ASAP7_75t_L g18623 ( 
.A(n_18251),
.Y(n_18623)
);

INVx4_ASAP7_75t_L g18624 ( 
.A(n_18244),
.Y(n_18624)
);

AND2x2_ASAP7_75t_SL g18625 ( 
.A(n_18188),
.B(n_9060),
.Y(n_18625)
);

INVx2_ASAP7_75t_L g18626 ( 
.A(n_18092),
.Y(n_18626)
);

INVx2_ASAP7_75t_L g18627 ( 
.A(n_18346),
.Y(n_18627)
);

OR2x2_ASAP7_75t_L g18628 ( 
.A(n_17953),
.B(n_11378),
.Y(n_18628)
);

NAND2xp5_ASAP7_75t_L g18629 ( 
.A(n_17916),
.B(n_11378),
.Y(n_18629)
);

INVx1_ASAP7_75t_L g18630 ( 
.A(n_18117),
.Y(n_18630)
);

OR2x2_ASAP7_75t_L g18631 ( 
.A(n_17951),
.B(n_11382),
.Y(n_18631)
);

NOR2x1_ASAP7_75t_L g18632 ( 
.A(n_18411),
.B(n_11382),
.Y(n_18632)
);

NAND2xp5_ASAP7_75t_L g18633 ( 
.A(n_18193),
.B(n_11402),
.Y(n_18633)
);

INVx1_ASAP7_75t_SL g18634 ( 
.A(n_17902),
.Y(n_18634)
);

OR2x2_ASAP7_75t_L g18635 ( 
.A(n_17941),
.B(n_11402),
.Y(n_18635)
);

NAND2xp5_ASAP7_75t_L g18636 ( 
.A(n_18077),
.B(n_11407),
.Y(n_18636)
);

NAND2xp5_ASAP7_75t_L g18637 ( 
.A(n_18081),
.B(n_11407),
.Y(n_18637)
);

AND2x4_ASAP7_75t_L g18638 ( 
.A(n_18140),
.B(n_9186),
.Y(n_18638)
);

BUFx2_ASAP7_75t_SL g18639 ( 
.A(n_18141),
.Y(n_18639)
);

OR2x2_ASAP7_75t_L g18640 ( 
.A(n_17942),
.B(n_11422),
.Y(n_18640)
);

INVx1_ASAP7_75t_L g18641 ( 
.A(n_18108),
.Y(n_18641)
);

OR2x2_ASAP7_75t_L g18642 ( 
.A(n_17969),
.B(n_11422),
.Y(n_18642)
);

INVx2_ASAP7_75t_L g18643 ( 
.A(n_18170),
.Y(n_18643)
);

OR2x2_ASAP7_75t_L g18644 ( 
.A(n_17905),
.B(n_10748),
.Y(n_18644)
);

INVx1_ASAP7_75t_L g18645 ( 
.A(n_18109),
.Y(n_18645)
);

NAND2xp5_ASAP7_75t_L g18646 ( 
.A(n_18130),
.B(n_11231),
.Y(n_18646)
);

AND2x2_ASAP7_75t_L g18647 ( 
.A(n_18343),
.B(n_9698),
.Y(n_18647)
);

NAND2xp5_ASAP7_75t_L g18648 ( 
.A(n_18131),
.B(n_11231),
.Y(n_18648)
);

INVx1_ASAP7_75t_L g18649 ( 
.A(n_18139),
.Y(n_18649)
);

OR2x6_ASAP7_75t_L g18650 ( 
.A(n_18386),
.B(n_10027),
.Y(n_18650)
);

NAND2xp67_ASAP7_75t_L g18651 ( 
.A(n_18426),
.B(n_11277),
.Y(n_18651)
);

OR2x2_ASAP7_75t_L g18652 ( 
.A(n_18216),
.B(n_10748),
.Y(n_18652)
);

AND2x2_ASAP7_75t_L g18653 ( 
.A(n_18043),
.B(n_9698),
.Y(n_18653)
);

NAND3xp33_ASAP7_75t_L g18654 ( 
.A(n_18218),
.B(n_10026),
.C(n_10007),
.Y(n_18654)
);

INVx1_ASAP7_75t_L g18655 ( 
.A(n_17891),
.Y(n_18655)
);

OR2x2_ASAP7_75t_L g18656 ( 
.A(n_17972),
.B(n_10748),
.Y(n_18656)
);

INVx1_ASAP7_75t_L g18657 ( 
.A(n_18253),
.Y(n_18657)
);

OR2x2_ASAP7_75t_L g18658 ( 
.A(n_18049),
.B(n_10748),
.Y(n_18658)
);

OAI21xp5_ASAP7_75t_L g18659 ( 
.A1(n_18327),
.A2(n_18197),
.B(n_18182),
.Y(n_18659)
);

OAI31xp33_ASAP7_75t_L g18660 ( 
.A1(n_18275),
.A2(n_9001),
.A3(n_9294),
.B(n_9108),
.Y(n_18660)
);

INVxp67_ASAP7_75t_SL g18661 ( 
.A(n_18396),
.Y(n_18661)
);

INVx1_ASAP7_75t_L g18662 ( 
.A(n_18029),
.Y(n_18662)
);

OR2x2_ASAP7_75t_L g18663 ( 
.A(n_18214),
.B(n_11522),
.Y(n_18663)
);

AND2x2_ASAP7_75t_L g18664 ( 
.A(n_18241),
.B(n_9698),
.Y(n_18664)
);

HB1xp67_ASAP7_75t_L g18665 ( 
.A(n_17948),
.Y(n_18665)
);

INVx1_ASAP7_75t_L g18666 ( 
.A(n_18042),
.Y(n_18666)
);

AOI32xp33_ASAP7_75t_L g18667 ( 
.A1(n_18001),
.A2(n_9013),
.A3(n_9075),
.B1(n_9008),
.B2(n_8977),
.Y(n_18667)
);

AND2x2_ASAP7_75t_L g18668 ( 
.A(n_18371),
.B(n_9698),
.Y(n_18668)
);

INVx1_ASAP7_75t_L g18669 ( 
.A(n_18158),
.Y(n_18669)
);

AND2x2_ASAP7_75t_L g18670 ( 
.A(n_18165),
.B(n_9698),
.Y(n_18670)
);

INVx2_ASAP7_75t_L g18671 ( 
.A(n_18127),
.Y(n_18671)
);

OR2x2_ASAP7_75t_L g18672 ( 
.A(n_18242),
.B(n_11522),
.Y(n_18672)
);

NAND2xp5_ASAP7_75t_SL g18673 ( 
.A(n_18121),
.B(n_10048),
.Y(n_18673)
);

INVx1_ASAP7_75t_L g18674 ( 
.A(n_18189),
.Y(n_18674)
);

OR2x2_ASAP7_75t_L g18675 ( 
.A(n_18164),
.B(n_11522),
.Y(n_18675)
);

INVx1_ASAP7_75t_L g18676 ( 
.A(n_17994),
.Y(n_18676)
);

AND2x2_ASAP7_75t_L g18677 ( 
.A(n_18058),
.B(n_9698),
.Y(n_18677)
);

INVx1_ASAP7_75t_L g18678 ( 
.A(n_18000),
.Y(n_18678)
);

INVxp67_ASAP7_75t_L g18679 ( 
.A(n_18098),
.Y(n_18679)
);

NAND2xp5_ASAP7_75t_L g18680 ( 
.A(n_18176),
.B(n_11231),
.Y(n_18680)
);

INVx1_ASAP7_75t_L g18681 ( 
.A(n_18017),
.Y(n_18681)
);

NAND2xp33_ASAP7_75t_L g18682 ( 
.A(n_18233),
.B(n_9060),
.Y(n_18682)
);

NAND2xp5_ASAP7_75t_L g18683 ( 
.A(n_18344),
.B(n_11231),
.Y(n_18683)
);

INVx2_ASAP7_75t_SL g18684 ( 
.A(n_18433),
.Y(n_18684)
);

AND2x2_ASAP7_75t_L g18685 ( 
.A(n_18020),
.B(n_9731),
.Y(n_18685)
);

AND2x2_ASAP7_75t_L g18686 ( 
.A(n_18362),
.B(n_9731),
.Y(n_18686)
);

INVx1_ASAP7_75t_L g18687 ( 
.A(n_18022),
.Y(n_18687)
);

INVxp67_ASAP7_75t_L g18688 ( 
.A(n_18002),
.Y(n_18688)
);

OAI21xp5_ASAP7_75t_L g18689 ( 
.A1(n_18089),
.A2(n_10699),
.B(n_10668),
.Y(n_18689)
);

INVx1_ASAP7_75t_L g18690 ( 
.A(n_18280),
.Y(n_18690)
);

INVx1_ASAP7_75t_L g18691 ( 
.A(n_17958),
.Y(n_18691)
);

AND2x2_ASAP7_75t_L g18692 ( 
.A(n_18294),
.B(n_9731),
.Y(n_18692)
);

INVx1_ASAP7_75t_L g18693 ( 
.A(n_17977),
.Y(n_18693)
);

AOI22xp5_ASAP7_75t_L g18694 ( 
.A1(n_18183),
.A2(n_11367),
.B1(n_10048),
.B2(n_10181),
.Y(n_18694)
);

OR2x2_ASAP7_75t_L g18695 ( 
.A(n_18191),
.B(n_11522),
.Y(n_18695)
);

NOR2xp67_ASAP7_75t_L g18696 ( 
.A(n_18425),
.B(n_9587),
.Y(n_18696)
);

INVx2_ASAP7_75t_L g18697 ( 
.A(n_18122),
.Y(n_18697)
);

NAND2xp5_ASAP7_75t_L g18698 ( 
.A(n_18344),
.B(n_11231),
.Y(n_18698)
);

AOI22xp5_ASAP7_75t_L g18699 ( 
.A1(n_18148),
.A2(n_11367),
.B1(n_10048),
.B2(n_10181),
.Y(n_18699)
);

AND2x2_ASAP7_75t_L g18700 ( 
.A(n_18298),
.B(n_9731),
.Y(n_18700)
);

OAI22xp5_ASAP7_75t_L g18701 ( 
.A1(n_18044),
.A2(n_10110),
.B1(n_10181),
.B2(n_10048),
.Y(n_18701)
);

INVx1_ASAP7_75t_L g18702 ( 
.A(n_17986),
.Y(n_18702)
);

NOR2xp33_ASAP7_75t_L g18703 ( 
.A(n_18150),
.B(n_7996),
.Y(n_18703)
);

INVx2_ASAP7_75t_SL g18704 ( 
.A(n_18436),
.Y(n_18704)
);

INVx2_ASAP7_75t_L g18705 ( 
.A(n_18125),
.Y(n_18705)
);

NAND2x1p5_ASAP7_75t_L g18706 ( 
.A(n_18259),
.B(n_9587),
.Y(n_18706)
);

NOR2xp33_ASAP7_75t_L g18707 ( 
.A(n_18159),
.B(n_7996),
.Y(n_18707)
);

INVx1_ASAP7_75t_L g18708 ( 
.A(n_17987),
.Y(n_18708)
);

INVx2_ASAP7_75t_L g18709 ( 
.A(n_18161),
.Y(n_18709)
);

AND2x2_ASAP7_75t_L g18710 ( 
.A(n_18359),
.B(n_9731),
.Y(n_18710)
);

INVx1_ASAP7_75t_L g18711 ( 
.A(n_17988),
.Y(n_18711)
);

INVx1_ASAP7_75t_SL g18712 ( 
.A(n_18105),
.Y(n_18712)
);

NAND2x1_ASAP7_75t_L g18713 ( 
.A(n_17948),
.B(n_10191),
.Y(n_18713)
);

INVx1_ASAP7_75t_L g18714 ( 
.A(n_17990),
.Y(n_18714)
);

NAND2xp5_ASAP7_75t_L g18715 ( 
.A(n_18420),
.B(n_11236),
.Y(n_18715)
);

OAI21xp33_ASAP7_75t_L g18716 ( 
.A1(n_18135),
.A2(n_10081),
.B(n_9993),
.Y(n_18716)
);

INVx2_ASAP7_75t_L g18717 ( 
.A(n_18207),
.Y(n_18717)
);

AND2x4_ASAP7_75t_SL g18718 ( 
.A(n_18103),
.B(n_7782),
.Y(n_18718)
);

AND2x2_ASAP7_75t_L g18719 ( 
.A(n_18401),
.B(n_9731),
.Y(n_18719)
);

OR2x2_ASAP7_75t_L g18720 ( 
.A(n_18171),
.B(n_11522),
.Y(n_18720)
);

OR2x2_ASAP7_75t_L g18721 ( 
.A(n_18174),
.B(n_11522),
.Y(n_18721)
);

INVx1_ASAP7_75t_L g18722 ( 
.A(n_18175),
.Y(n_18722)
);

NAND2xp5_ASAP7_75t_L g18723 ( 
.A(n_18308),
.B(n_11236),
.Y(n_18723)
);

NAND2xp5_ASAP7_75t_L g18724 ( 
.A(n_18358),
.B(n_11236),
.Y(n_18724)
);

INVx1_ASAP7_75t_L g18725 ( 
.A(n_18177),
.Y(n_18725)
);

BUFx2_ASAP7_75t_L g18726 ( 
.A(n_18103),
.Y(n_18726)
);

AND2x2_ASAP7_75t_L g18727 ( 
.A(n_18021),
.B(n_9731),
.Y(n_18727)
);

INVx1_ASAP7_75t_L g18728 ( 
.A(n_18178),
.Y(n_18728)
);

INVx1_ASAP7_75t_L g18729 ( 
.A(n_18192),
.Y(n_18729)
);

INVxp67_ASAP7_75t_L g18730 ( 
.A(n_17996),
.Y(n_18730)
);

INVx1_ASAP7_75t_L g18731 ( 
.A(n_18204),
.Y(n_18731)
);

OR2x2_ASAP7_75t_L g18732 ( 
.A(n_18210),
.B(n_11522),
.Y(n_18732)
);

OR2x2_ASAP7_75t_L g18733 ( 
.A(n_18137),
.B(n_11619),
.Y(n_18733)
);

INVx2_ASAP7_75t_SL g18734 ( 
.A(n_18375),
.Y(n_18734)
);

OR2x6_ASAP7_75t_L g18735 ( 
.A(n_18389),
.B(n_10191),
.Y(n_18735)
);

BUFx6f_ASAP7_75t_L g18736 ( 
.A(n_18255),
.Y(n_18736)
);

NAND2xp5_ASAP7_75t_L g18737 ( 
.A(n_18380),
.B(n_11236),
.Y(n_18737)
);

AND2x2_ASAP7_75t_L g18738 ( 
.A(n_18023),
.B(n_9731),
.Y(n_18738)
);

OR2x2_ASAP7_75t_L g18739 ( 
.A(n_18138),
.B(n_11619),
.Y(n_18739)
);

AND2x2_ASAP7_75t_L g18740 ( 
.A(n_18126),
.B(n_9731),
.Y(n_18740)
);

INVx1_ASAP7_75t_L g18741 ( 
.A(n_18257),
.Y(n_18741)
);

INVx2_ASAP7_75t_L g18742 ( 
.A(n_18143),
.Y(n_18742)
);

AND2x4_ASAP7_75t_L g18743 ( 
.A(n_18268),
.B(n_9186),
.Y(n_18743)
);

INVx1_ASAP7_75t_L g18744 ( 
.A(n_17989),
.Y(n_18744)
);

INVx2_ASAP7_75t_L g18745 ( 
.A(n_18149),
.Y(n_18745)
);

INVx1_ASAP7_75t_L g18746 ( 
.A(n_18157),
.Y(n_18746)
);

OAI21xp5_ASAP7_75t_L g18747 ( 
.A1(n_18225),
.A2(n_10699),
.B(n_10668),
.Y(n_18747)
);

INVx1_ASAP7_75t_L g18748 ( 
.A(n_18383),
.Y(n_18748)
);

HB1xp67_ASAP7_75t_L g18749 ( 
.A(n_18273),
.Y(n_18749)
);

INVx1_ASAP7_75t_L g18750 ( 
.A(n_18397),
.Y(n_18750)
);

NAND2xp5_ASAP7_75t_SL g18751 ( 
.A(n_18304),
.B(n_10110),
.Y(n_18751)
);

NAND2xp5_ASAP7_75t_L g18752 ( 
.A(n_18414),
.B(n_11236),
.Y(n_18752)
);

INVx1_ASAP7_75t_L g18753 ( 
.A(n_18403),
.Y(n_18753)
);

AND2x2_ASAP7_75t_L g18754 ( 
.A(n_18283),
.B(n_9768),
.Y(n_18754)
);

NAND2xp5_ASAP7_75t_L g18755 ( 
.A(n_18405),
.B(n_11311),
.Y(n_18755)
);

AND2x2_ASAP7_75t_L g18756 ( 
.A(n_18269),
.B(n_9768),
.Y(n_18756)
);

INVx2_ASAP7_75t_SL g18757 ( 
.A(n_18128),
.Y(n_18757)
);

NOR2xp67_ASAP7_75t_L g18758 ( 
.A(n_18297),
.B(n_9587),
.Y(n_18758)
);

AND2x4_ASAP7_75t_L g18759 ( 
.A(n_18333),
.B(n_9186),
.Y(n_18759)
);

INVx1_ASAP7_75t_L g18760 ( 
.A(n_18360),
.Y(n_18760)
);

INVx2_ASAP7_75t_L g18761 ( 
.A(n_18136),
.Y(n_18761)
);

OR2x2_ASAP7_75t_L g18762 ( 
.A(n_18145),
.B(n_11619),
.Y(n_18762)
);

INVx1_ASAP7_75t_L g18763 ( 
.A(n_18271),
.Y(n_18763)
);

AND2x2_ASAP7_75t_L g18764 ( 
.A(n_18019),
.B(n_9768),
.Y(n_18764)
);

AND2x2_ASAP7_75t_L g18765 ( 
.A(n_18013),
.B(n_9768),
.Y(n_18765)
);

INVx1_ASAP7_75t_L g18766 ( 
.A(n_18243),
.Y(n_18766)
);

NAND2xp5_ASAP7_75t_L g18767 ( 
.A(n_18104),
.B(n_11311),
.Y(n_18767)
);

INVx1_ASAP7_75t_L g18768 ( 
.A(n_18281),
.Y(n_18768)
);

INVx1_ASAP7_75t_L g18769 ( 
.A(n_18286),
.Y(n_18769)
);

HB1xp67_ASAP7_75t_L g18770 ( 
.A(n_18311),
.Y(n_18770)
);

INVx2_ASAP7_75t_L g18771 ( 
.A(n_18169),
.Y(n_18771)
);

OR2x2_ASAP7_75t_L g18772 ( 
.A(n_18152),
.B(n_18112),
.Y(n_18772)
);

INVx1_ASAP7_75t_L g18773 ( 
.A(n_18291),
.Y(n_18773)
);

AND2x2_ASAP7_75t_L g18774 ( 
.A(n_18015),
.B(n_9768),
.Y(n_18774)
);

NAND2xp5_ASAP7_75t_L g18775 ( 
.A(n_17997),
.B(n_11311),
.Y(n_18775)
);

NAND2xp5_ASAP7_75t_L g18776 ( 
.A(n_18316),
.B(n_11311),
.Y(n_18776)
);

NAND2xp5_ASAP7_75t_L g18777 ( 
.A(n_18301),
.B(n_11311),
.Y(n_18777)
);

AND2x4_ASAP7_75t_L g18778 ( 
.A(n_18276),
.B(n_9186),
.Y(n_18778)
);

OR2x2_ASAP7_75t_L g18779 ( 
.A(n_18079),
.B(n_11619),
.Y(n_18779)
);

INVx1_ASAP7_75t_L g18780 ( 
.A(n_18306),
.Y(n_18780)
);

AND2x2_ASAP7_75t_L g18781 ( 
.A(n_18120),
.B(n_9768),
.Y(n_18781)
);

NAND2x1_ASAP7_75t_SL g18782 ( 
.A(n_18444),
.B(n_9787),
.Y(n_18782)
);

AND2x2_ASAP7_75t_L g18783 ( 
.A(n_18167),
.B(n_9768),
.Y(n_18783)
);

NAND2xp5_ASAP7_75t_L g18784 ( 
.A(n_18314),
.B(n_11563),
.Y(n_18784)
);

NAND2xp5_ASAP7_75t_L g18785 ( 
.A(n_18317),
.B(n_11563),
.Y(n_18785)
);

AND2x2_ASAP7_75t_L g18786 ( 
.A(n_18234),
.B(n_9768),
.Y(n_18786)
);

INVx2_ASAP7_75t_L g18787 ( 
.A(n_18209),
.Y(n_18787)
);

OR2x2_ASAP7_75t_L g18788 ( 
.A(n_18061),
.B(n_11619),
.Y(n_18788)
);

INVx1_ASAP7_75t_L g18789 ( 
.A(n_18318),
.Y(n_18789)
);

NOR2xp33_ASAP7_75t_L g18790 ( 
.A(n_18330),
.B(n_7996),
.Y(n_18790)
);

INVx1_ASAP7_75t_L g18791 ( 
.A(n_18332),
.Y(n_18791)
);

NAND2xp5_ASAP7_75t_L g18792 ( 
.A(n_18334),
.B(n_18337),
.Y(n_18792)
);

BUFx2_ASAP7_75t_L g18793 ( 
.A(n_18107),
.Y(n_18793)
);

INVx1_ASAP7_75t_L g18794 ( 
.A(n_18338),
.Y(n_18794)
);

AND2x2_ASAP7_75t_L g18795 ( 
.A(n_18212),
.B(n_9768),
.Y(n_18795)
);

AOI21xp33_ASAP7_75t_L g18796 ( 
.A1(n_18287),
.A2(n_11367),
.B(n_10897),
.Y(n_18796)
);

AND2x2_ASAP7_75t_L g18797 ( 
.A(n_18223),
.B(n_18228),
.Y(n_18797)
);

INVx1_ASAP7_75t_L g18798 ( 
.A(n_18340),
.Y(n_18798)
);

NAND2xp5_ASAP7_75t_L g18799 ( 
.A(n_18342),
.B(n_11563),
.Y(n_18799)
);

NAND2x1_ASAP7_75t_L g18800 ( 
.A(n_18107),
.B(n_10191),
.Y(n_18800)
);

INVx2_ASAP7_75t_L g18801 ( 
.A(n_18134),
.Y(n_18801)
);

OR2x2_ASAP7_75t_L g18802 ( 
.A(n_18111),
.B(n_11619),
.Y(n_18802)
);

NOR2xp67_ASAP7_75t_L g18803 ( 
.A(n_18113),
.B(n_9636),
.Y(n_18803)
);

INVx1_ASAP7_75t_L g18804 ( 
.A(n_18351),
.Y(n_18804)
);

INVx1_ASAP7_75t_L g18805 ( 
.A(n_18352),
.Y(n_18805)
);

NAND2xp5_ASAP7_75t_L g18806 ( 
.A(n_18354),
.B(n_11563),
.Y(n_18806)
);

INVx1_ASAP7_75t_L g18807 ( 
.A(n_18355),
.Y(n_18807)
);

AND2x4_ASAP7_75t_L g18808 ( 
.A(n_17999),
.B(n_9186),
.Y(n_18808)
);

INVx1_ASAP7_75t_L g18809 ( 
.A(n_18366),
.Y(n_18809)
);

AND2x2_ASAP7_75t_L g18810 ( 
.A(n_18185),
.B(n_9777),
.Y(n_18810)
);

NAND2xp5_ASAP7_75t_L g18811 ( 
.A(n_18370),
.B(n_11563),
.Y(n_18811)
);

AND2x2_ASAP7_75t_L g18812 ( 
.A(n_18187),
.B(n_9777),
.Y(n_18812)
);

AND2x2_ASAP7_75t_L g18813 ( 
.A(n_18235),
.B(n_9777),
.Y(n_18813)
);

NAND2xp5_ASAP7_75t_SL g18814 ( 
.A(n_18038),
.B(n_18051),
.Y(n_18814)
);

HB1xp67_ASAP7_75t_L g18815 ( 
.A(n_18435),
.Y(n_18815)
);

NAND2x1p5_ASAP7_75t_L g18816 ( 
.A(n_18374),
.B(n_9636),
.Y(n_18816)
);

INVx1_ASAP7_75t_L g18817 ( 
.A(n_18376),
.Y(n_18817)
);

NOR2xp33_ASAP7_75t_L g18818 ( 
.A(n_18378),
.B(n_7996),
.Y(n_18818)
);

INVx1_ASAP7_75t_L g18819 ( 
.A(n_18409),
.Y(n_18819)
);

AND2x2_ASAP7_75t_L g18820 ( 
.A(n_18200),
.B(n_9777),
.Y(n_18820)
);

OR2x2_ASAP7_75t_L g18821 ( 
.A(n_18272),
.B(n_11619),
.Y(n_18821)
);

AND2x2_ASAP7_75t_L g18822 ( 
.A(n_18202),
.B(n_9777),
.Y(n_18822)
);

INVx2_ASAP7_75t_L g18823 ( 
.A(n_18203),
.Y(n_18823)
);

OR2x2_ASAP7_75t_SL g18824 ( 
.A(n_18213),
.B(n_10007),
.Y(n_18824)
);

AND2x2_ASAP7_75t_L g18825 ( 
.A(n_18394),
.B(n_9777),
.Y(n_18825)
);

INVx1_ASAP7_75t_L g18826 ( 
.A(n_18413),
.Y(n_18826)
);

INVx1_ASAP7_75t_L g18827 ( 
.A(n_18418),
.Y(n_18827)
);

AND2x2_ASAP7_75t_L g18828 ( 
.A(n_18372),
.B(n_18382),
.Y(n_18828)
);

INVx1_ASAP7_75t_L g18829 ( 
.A(n_18364),
.Y(n_18829)
);

NAND2xp5_ASAP7_75t_L g18830 ( 
.A(n_18296),
.B(n_11563),
.Y(n_18830)
);

AND2x2_ASAP7_75t_L g18831 ( 
.A(n_18395),
.B(n_9777),
.Y(n_18831)
);

AND3x1_ASAP7_75t_L g18832 ( 
.A(n_18325),
.B(n_9659),
.C(n_9620),
.Y(n_18832)
);

NAND2xp5_ASAP7_75t_L g18833 ( 
.A(n_18274),
.B(n_11563),
.Y(n_18833)
);

INVx1_ASAP7_75t_L g18834 ( 
.A(n_18367),
.Y(n_18834)
);

INVx1_ASAP7_75t_L g18835 ( 
.A(n_18369),
.Y(n_18835)
);

INVx2_ASAP7_75t_L g18836 ( 
.A(n_18266),
.Y(n_18836)
);

INVx1_ASAP7_75t_L g18837 ( 
.A(n_18408),
.Y(n_18837)
);

INVx1_ASAP7_75t_L g18838 ( 
.A(n_18416),
.Y(n_18838)
);

AND2x2_ASAP7_75t_L g18839 ( 
.A(n_18398),
.B(n_9777),
.Y(n_18839)
);

INVxp67_ASAP7_75t_L g18840 ( 
.A(n_18432),
.Y(n_18840)
);

INVx2_ASAP7_75t_L g18841 ( 
.A(n_18419),
.Y(n_18841)
);

INVx2_ASAP7_75t_L g18842 ( 
.A(n_18270),
.Y(n_18842)
);

AND2x2_ASAP7_75t_L g18843 ( 
.A(n_18406),
.B(n_18412),
.Y(n_18843)
);

INVx1_ASAP7_75t_L g18844 ( 
.A(n_18417),
.Y(n_18844)
);

INVx1_ASAP7_75t_L g18845 ( 
.A(n_18224),
.Y(n_18845)
);

AND2x2_ASAP7_75t_L g18846 ( 
.A(n_18277),
.B(n_9777),
.Y(n_18846)
);

NOR2xp33_ASAP7_75t_L g18847 ( 
.A(n_18434),
.B(n_7996),
.Y(n_18847)
);

AND2x2_ASAP7_75t_L g18848 ( 
.A(n_18289),
.B(n_9785),
.Y(n_18848)
);

INVxp67_ASAP7_75t_L g18849 ( 
.A(n_18082),
.Y(n_18849)
);

OR2x2_ASAP7_75t_L g18850 ( 
.A(n_18264),
.B(n_11619),
.Y(n_18850)
);

NAND2xp5_ASAP7_75t_L g18851 ( 
.A(n_18438),
.B(n_11563),
.Y(n_18851)
);

INVx2_ASAP7_75t_L g18852 ( 
.A(n_18328),
.Y(n_18852)
);

NAND2xp5_ASAP7_75t_L g18853 ( 
.A(n_18440),
.B(n_10473),
.Y(n_18853)
);

INVxp67_ASAP7_75t_L g18854 ( 
.A(n_18085),
.Y(n_18854)
);

AOI21xp5_ASAP7_75t_SL g18855 ( 
.A1(n_18008),
.A2(n_11904),
.B(n_10180),
.Y(n_18855)
);

NAND2xp67_ASAP7_75t_L g18856 ( 
.A(n_18066),
.B(n_11277),
.Y(n_18856)
);

INVx1_ASAP7_75t_L g18857 ( 
.A(n_18230),
.Y(n_18857)
);

NAND2xp5_ASAP7_75t_L g18858 ( 
.A(n_18028),
.B(n_18246),
.Y(n_18858)
);

INVx1_ASAP7_75t_L g18859 ( 
.A(n_18181),
.Y(n_18859)
);

OR2x2_ASAP7_75t_L g18860 ( 
.A(n_18156),
.B(n_11617),
.Y(n_18860)
);

NAND2xp5_ASAP7_75t_L g18861 ( 
.A(n_18249),
.B(n_10473),
.Y(n_18861)
);

INVx2_ASAP7_75t_SL g18862 ( 
.A(n_18379),
.Y(n_18862)
);

INVx3_ASAP7_75t_SL g18863 ( 
.A(n_18292),
.Y(n_18863)
);

INVx2_ASAP7_75t_L g18864 ( 
.A(n_18345),
.Y(n_18864)
);

OR2x2_ASAP7_75t_L g18865 ( 
.A(n_18236),
.B(n_18324),
.Y(n_18865)
);

INVx1_ASAP7_75t_L g18866 ( 
.A(n_18184),
.Y(n_18866)
);

INVx2_ASAP7_75t_L g18867 ( 
.A(n_18347),
.Y(n_18867)
);

INVx1_ASAP7_75t_L g18868 ( 
.A(n_18279),
.Y(n_18868)
);

HB1xp67_ASAP7_75t_L g18869 ( 
.A(n_18261),
.Y(n_18869)
);

INVxp67_ASAP7_75t_L g18870 ( 
.A(n_18123),
.Y(n_18870)
);

AOI22xp5_ASAP7_75t_L g18871 ( 
.A1(n_18385),
.A2(n_11367),
.B1(n_10110),
.B2(n_10181),
.Y(n_18871)
);

INVx1_ASAP7_75t_L g18872 ( 
.A(n_18285),
.Y(n_18872)
);

INVx1_ASAP7_75t_L g18873 ( 
.A(n_18299),
.Y(n_18873)
);

INVx1_ASAP7_75t_L g18874 ( 
.A(n_18326),
.Y(n_18874)
);

OR2x2_ASAP7_75t_L g18875 ( 
.A(n_18222),
.B(n_11617),
.Y(n_18875)
);

NAND2xp5_ASAP7_75t_L g18876 ( 
.A(n_18350),
.B(n_10473),
.Y(n_18876)
);

INVx1_ASAP7_75t_L g18877 ( 
.A(n_18349),
.Y(n_18877)
);

INVx2_ASAP7_75t_SL g18878 ( 
.A(n_18381),
.Y(n_18878)
);

INVx1_ASAP7_75t_L g18879 ( 
.A(n_18353),
.Y(n_18879)
);

NAND2xp5_ASAP7_75t_L g18880 ( 
.A(n_18368),
.B(n_10473),
.Y(n_18880)
);

INVx2_ASAP7_75t_L g18881 ( 
.A(n_18415),
.Y(n_18881)
);

AND2x2_ASAP7_75t_L g18882 ( 
.A(n_18387),
.B(n_9785),
.Y(n_18882)
);

INVxp67_ASAP7_75t_SL g18883 ( 
.A(n_18258),
.Y(n_18883)
);

INVx1_ASAP7_75t_SL g18884 ( 
.A(n_18186),
.Y(n_18884)
);

NAND2xp5_ASAP7_75t_L g18885 ( 
.A(n_18039),
.B(n_10473),
.Y(n_18885)
);

INVxp67_ASAP7_75t_L g18886 ( 
.A(n_18100),
.Y(n_18886)
);

AND2x2_ASAP7_75t_L g18887 ( 
.A(n_18388),
.B(n_9785),
.Y(n_18887)
);

AND2x2_ASAP7_75t_L g18888 ( 
.A(n_18292),
.B(n_9785),
.Y(n_18888)
);

INVx1_ASAP7_75t_L g18889 ( 
.A(n_18356),
.Y(n_18889)
);

NAND2xp5_ASAP7_75t_L g18890 ( 
.A(n_18080),
.B(n_10473),
.Y(n_18890)
);

INVx1_ASAP7_75t_L g18891 ( 
.A(n_18365),
.Y(n_18891)
);

AND2x2_ASAP7_75t_L g18892 ( 
.A(n_18427),
.B(n_9785),
.Y(n_18892)
);

NAND2xp5_ASAP7_75t_L g18893 ( 
.A(n_18096),
.B(n_10473),
.Y(n_18893)
);

A2O1A1Ixp33_ASAP7_75t_L g18894 ( 
.A1(n_18310),
.A2(n_10868),
.B(n_10871),
.C(n_11607),
.Y(n_18894)
);

AND2x2_ASAP7_75t_L g18895 ( 
.A(n_18431),
.B(n_9785),
.Y(n_18895)
);

INVx2_ASAP7_75t_L g18896 ( 
.A(n_18256),
.Y(n_18896)
);

NAND2xp5_ASAP7_75t_L g18897 ( 
.A(n_18099),
.B(n_10473),
.Y(n_18897)
);

AND2x2_ASAP7_75t_L g18898 ( 
.A(n_18309),
.B(n_18290),
.Y(n_18898)
);

NAND2xp5_ASAP7_75t_L g18899 ( 
.A(n_18180),
.B(n_10531),
.Y(n_18899)
);

OR2x6_ASAP7_75t_L g18900 ( 
.A(n_18227),
.B(n_10191),
.Y(n_18900)
);

BUFx2_ASAP7_75t_L g18901 ( 
.A(n_18201),
.Y(n_18901)
);

INVx2_ASAP7_75t_L g18902 ( 
.A(n_18404),
.Y(n_18902)
);

INVx1_ASAP7_75t_L g18903 ( 
.A(n_18377),
.Y(n_18903)
);

INVxp33_ASAP7_75t_L g18904 ( 
.A(n_18254),
.Y(n_18904)
);

NAND2xp5_ASAP7_75t_L g18905 ( 
.A(n_18488),
.B(n_18295),
.Y(n_18905)
);

OAI21xp5_ASAP7_75t_L g18906 ( 
.A1(n_18492),
.A2(n_18129),
.B(n_18402),
.Y(n_18906)
);

NAND2xp5_ASAP7_75t_L g18907 ( 
.A(n_18462),
.B(n_18040),
.Y(n_18907)
);

NAND2xp5_ASAP7_75t_L g18908 ( 
.A(n_18470),
.B(n_18070),
.Y(n_18908)
);

NAND2xp5_ASAP7_75t_L g18909 ( 
.A(n_18531),
.B(n_18076),
.Y(n_18909)
);

O2A1O1Ixp5_ASAP7_75t_R g18910 ( 
.A1(n_18451),
.A2(n_18205),
.B(n_18154),
.C(n_18206),
.Y(n_18910)
);

INVx2_ASAP7_75t_L g18911 ( 
.A(n_18445),
.Y(n_18911)
);

NAND2xp5_ASAP7_75t_L g18912 ( 
.A(n_18472),
.B(n_18319),
.Y(n_18912)
);

NAND2xp5_ASAP7_75t_L g18913 ( 
.A(n_18624),
.B(n_18262),
.Y(n_18913)
);

INVx1_ASAP7_75t_L g18914 ( 
.A(n_18476),
.Y(n_18914)
);

INVx1_ASAP7_75t_L g18915 ( 
.A(n_18534),
.Y(n_18915)
);

INVx1_ASAP7_75t_L g18916 ( 
.A(n_18556),
.Y(n_18916)
);

INVx1_ASAP7_75t_L g18917 ( 
.A(n_18565),
.Y(n_18917)
);

OR2x2_ASAP7_75t_L g18918 ( 
.A(n_18446),
.B(n_18173),
.Y(n_18918)
);

AND2x2_ASAP7_75t_L g18919 ( 
.A(n_18591),
.B(n_18265),
.Y(n_18919)
);

AND2x4_ASAP7_75t_L g18920 ( 
.A(n_18486),
.B(n_18006),
.Y(n_18920)
);

NOR2x1_ASAP7_75t_L g18921 ( 
.A(n_18522),
.B(n_18065),
.Y(n_18921)
);

NAND2xp5_ASAP7_75t_L g18922 ( 
.A(n_18511),
.B(n_18067),
.Y(n_18922)
);

AND2x2_ASAP7_75t_L g18923 ( 
.A(n_18452),
.B(n_18307),
.Y(n_18923)
);

HB1xp67_ASAP7_75t_L g18924 ( 
.A(n_18453),
.Y(n_18924)
);

HB1xp67_ASAP7_75t_L g18925 ( 
.A(n_18606),
.Y(n_18925)
);

NAND2xp5_ASAP7_75t_L g18926 ( 
.A(n_18623),
.B(n_18336),
.Y(n_18926)
);

INVx1_ASAP7_75t_L g18927 ( 
.A(n_18478),
.Y(n_18927)
);

AND2x2_ASAP7_75t_SL g18928 ( 
.A(n_18447),
.B(n_18198),
.Y(n_18928)
);

INVx3_ASAP7_75t_L g18929 ( 
.A(n_18477),
.Y(n_18929)
);

INVx1_ASAP7_75t_L g18930 ( 
.A(n_18665),
.Y(n_18930)
);

HB1xp67_ASAP7_75t_L g18931 ( 
.A(n_18450),
.Y(n_18931)
);

AND2x2_ASAP7_75t_L g18932 ( 
.A(n_18600),
.B(n_18078),
.Y(n_18932)
);

HB1xp67_ASAP7_75t_L g18933 ( 
.A(n_18454),
.Y(n_18933)
);

NAND2xp5_ASAP7_75t_L g18934 ( 
.A(n_18603),
.B(n_18357),
.Y(n_18934)
);

INVx1_ASAP7_75t_L g18935 ( 
.A(n_18590),
.Y(n_18935)
);

INVx1_ASAP7_75t_SL g18936 ( 
.A(n_18639),
.Y(n_18936)
);

NOR2xp33_ASAP7_75t_L g18937 ( 
.A(n_18582),
.B(n_18025),
.Y(n_18937)
);

INVx1_ASAP7_75t_L g18938 ( 
.A(n_18632),
.Y(n_18938)
);

NAND2xp5_ASAP7_75t_L g18939 ( 
.A(n_18502),
.B(n_18086),
.Y(n_18939)
);

INVx1_ASAP7_75t_L g18940 ( 
.A(n_18490),
.Y(n_18940)
);

OAI21xp33_ASAP7_75t_L g18941 ( 
.A1(n_18562),
.A2(n_18263),
.B(n_18101),
.Y(n_18941)
);

AND2x2_ASAP7_75t_L g18942 ( 
.A(n_18626),
.B(n_18114),
.Y(n_18942)
);

OR2x2_ASAP7_75t_L g18943 ( 
.A(n_18487),
.B(n_18195),
.Y(n_18943)
);

NAND2xp5_ASAP7_75t_L g18944 ( 
.A(n_18468),
.B(n_18231),
.Y(n_18944)
);

AND2x2_ASAP7_75t_L g18945 ( 
.A(n_18613),
.B(n_18643),
.Y(n_18945)
);

AND2x2_ASAP7_75t_L g18946 ( 
.A(n_18489),
.B(n_18363),
.Y(n_18946)
);

NAND4xp75_ASAP7_75t_L g18947 ( 
.A(n_18464),
.B(n_18056),
.C(n_18119),
.D(n_18208),
.Y(n_18947)
);

INVx2_ASAP7_75t_L g18948 ( 
.A(n_18782),
.Y(n_18948)
);

OAI21xp33_ASAP7_75t_L g18949 ( 
.A1(n_18501),
.A2(n_18528),
.B(n_18634),
.Y(n_18949)
);

INVx1_ASAP7_75t_SL g18950 ( 
.A(n_18508),
.Y(n_18950)
);

INVxp67_ASAP7_75t_L g18951 ( 
.A(n_18605),
.Y(n_18951)
);

INVx2_ASAP7_75t_SL g18952 ( 
.A(n_18713),
.Y(n_18952)
);

NAND2xp5_ASAP7_75t_L g18953 ( 
.A(n_18500),
.B(n_18505),
.Y(n_18953)
);

AND2x4_ASAP7_75t_L g18954 ( 
.A(n_18617),
.B(n_18248),
.Y(n_18954)
);

OR2x2_ASAP7_75t_L g18955 ( 
.A(n_18497),
.B(n_18199),
.Y(n_18955)
);

HB1xp67_ASAP7_75t_L g18956 ( 
.A(n_18456),
.Y(n_18956)
);

HB1xp67_ASAP7_75t_L g18957 ( 
.A(n_18619),
.Y(n_18957)
);

INVx1_ASAP7_75t_L g18958 ( 
.A(n_18842),
.Y(n_18958)
);

OAI22xp33_ASAP7_75t_L g18959 ( 
.A1(n_18448),
.A2(n_18331),
.B1(n_18407),
.B2(n_18303),
.Y(n_18959)
);

INVxp67_ASAP7_75t_L g18960 ( 
.A(n_18770),
.Y(n_18960)
);

NAND2x1p5_ASAP7_75t_L g18961 ( 
.A(n_18504),
.B(n_18115),
.Y(n_18961)
);

AND2x2_ASAP7_75t_L g18962 ( 
.A(n_18479),
.B(n_18093),
.Y(n_18962)
);

INVx1_ASAP7_75t_L g18963 ( 
.A(n_18651),
.Y(n_18963)
);

INVx1_ASAP7_75t_L g18964 ( 
.A(n_18461),
.Y(n_18964)
);

OR2x2_ASAP7_75t_L g18965 ( 
.A(n_18509),
.B(n_18510),
.Y(n_18965)
);

OAI22xp5_ASAP7_75t_L g18966 ( 
.A1(n_18466),
.A2(n_18313),
.B1(n_18320),
.B2(n_18315),
.Y(n_18966)
);

AND2x2_ASAP7_75t_L g18967 ( 
.A(n_18671),
.B(n_18240),
.Y(n_18967)
);

NAND3xp33_ASAP7_75t_SL g18968 ( 
.A(n_18469),
.B(n_17998),
.C(n_18384),
.Y(n_18968)
);

INVx1_ASAP7_75t_L g18969 ( 
.A(n_18584),
.Y(n_18969)
);

NAND3xp33_ASAP7_75t_SL g18970 ( 
.A(n_18659),
.B(n_18124),
.C(n_18252),
.Y(n_18970)
);

AND2x2_ASAP7_75t_L g18971 ( 
.A(n_18512),
.B(n_18322),
.Y(n_18971)
);

INVx1_ASAP7_75t_L g18972 ( 
.A(n_18498),
.Y(n_18972)
);

AND2x2_ASAP7_75t_L g18973 ( 
.A(n_18542),
.B(n_18312),
.Y(n_18973)
);

INVx1_ASAP7_75t_L g18974 ( 
.A(n_18749),
.Y(n_18974)
);

INVx1_ASAP7_75t_L g18975 ( 
.A(n_18459),
.Y(n_18975)
);

AND2x2_ASAP7_75t_L g18976 ( 
.A(n_18572),
.B(n_18392),
.Y(n_18976)
);

OR2x2_ASAP7_75t_L g18977 ( 
.A(n_18577),
.B(n_18190),
.Y(n_18977)
);

NAND2xp5_ASAP7_75t_L g18978 ( 
.A(n_18594),
.B(n_18059),
.Y(n_18978)
);

INVx2_ASAP7_75t_L g18979 ( 
.A(n_18697),
.Y(n_18979)
);

NAND2xp5_ASAP7_75t_L g18980 ( 
.A(n_18704),
.B(n_18393),
.Y(n_18980)
);

INVx1_ASAP7_75t_L g18981 ( 
.A(n_18460),
.Y(n_18981)
);

OR2x2_ASAP7_75t_L g18982 ( 
.A(n_18532),
.B(n_18429),
.Y(n_18982)
);

INVx1_ASAP7_75t_L g18983 ( 
.A(n_18465),
.Y(n_18983)
);

NAND2xp5_ASAP7_75t_L g18984 ( 
.A(n_18684),
.B(n_18116),
.Y(n_18984)
);

AND2x2_ASAP7_75t_L g18985 ( 
.A(n_18705),
.B(n_18219),
.Y(n_18985)
);

AND2x2_ASAP7_75t_L g18986 ( 
.A(n_18828),
.B(n_18430),
.Y(n_18986)
);

AND2x2_ASAP7_75t_L g18987 ( 
.A(n_18898),
.B(n_18391),
.Y(n_18987)
);

AND2x4_ASAP7_75t_L g18988 ( 
.A(n_18545),
.B(n_18548),
.Y(n_18988)
);

INVx1_ASAP7_75t_SL g18989 ( 
.A(n_18499),
.Y(n_18989)
);

NOR2xp33_ASAP7_75t_L g18990 ( 
.A(n_18588),
.B(n_18439),
.Y(n_18990)
);

INVx1_ASAP7_75t_L g18991 ( 
.A(n_18607),
.Y(n_18991)
);

INVx1_ASAP7_75t_L g18992 ( 
.A(n_18467),
.Y(n_18992)
);

NAND2x1p5_ASAP7_75t_L g18993 ( 
.A(n_18712),
.B(n_18267),
.Y(n_18993)
);

INVx2_ASAP7_75t_L g18994 ( 
.A(n_18515),
.Y(n_18994)
);

OR2x2_ASAP7_75t_L g18995 ( 
.A(n_18655),
.B(n_18424),
.Y(n_18995)
);

INVx1_ASAP7_75t_L g18996 ( 
.A(n_18856),
.Y(n_18996)
);

AND2x2_ASAP7_75t_L g18997 ( 
.A(n_18843),
.B(n_18045),
.Y(n_18997)
);

INVx1_ASAP7_75t_L g18998 ( 
.A(n_18629),
.Y(n_18998)
);

INVx1_ASAP7_75t_L g18999 ( 
.A(n_18475),
.Y(n_18999)
);

INVx1_ASAP7_75t_L g19000 ( 
.A(n_18661),
.Y(n_19000)
);

AND2x2_ASAP7_75t_L g19001 ( 
.A(n_18560),
.B(n_18329),
.Y(n_19001)
);

OAI21xp33_ASAP7_75t_L g19002 ( 
.A1(n_18677),
.A2(n_18030),
.B(n_18323),
.Y(n_19002)
);

AND2x2_ASAP7_75t_L g19003 ( 
.A(n_18836),
.B(n_18896),
.Y(n_19003)
);

AOI21xp5_ASAP7_75t_L g19004 ( 
.A1(n_18482),
.A2(n_18032),
.B(n_18005),
.Y(n_19004)
);

INVx1_ASAP7_75t_L g19005 ( 
.A(n_18495),
.Y(n_19005)
);

INVxp67_ASAP7_75t_SL g19006 ( 
.A(n_18457),
.Y(n_19006)
);

AOI211xp5_ASAP7_75t_L g19007 ( 
.A1(n_18483),
.A2(n_18335),
.B(n_18400),
.C(n_18443),
.Y(n_19007)
);

NOR2xp33_ASAP7_75t_L g19008 ( 
.A(n_18730),
.B(n_18341),
.Y(n_19008)
);

INVx1_ASAP7_75t_L g19009 ( 
.A(n_18513),
.Y(n_19009)
);

OR2x2_ASAP7_75t_L g19010 ( 
.A(n_18702),
.B(n_18410),
.Y(n_19010)
);

NAND2xp5_ASAP7_75t_L g19011 ( 
.A(n_18567),
.B(n_18250),
.Y(n_19011)
);

INVxp67_ASAP7_75t_L g19012 ( 
.A(n_18815),
.Y(n_19012)
);

AND2x2_ASAP7_75t_L g19013 ( 
.A(n_18708),
.B(n_18217),
.Y(n_19013)
);

AOI22xp5_ASAP7_75t_L g19014 ( 
.A1(n_18596),
.A2(n_10110),
.B1(n_10181),
.B2(n_11341),
.Y(n_19014)
);

NAND2xp5_ASAP7_75t_L g19015 ( 
.A(n_18711),
.B(n_10963),
.Y(n_19015)
);

NOR2xp33_ASAP7_75t_L g19016 ( 
.A(n_18741),
.B(n_7996),
.Y(n_19016)
);

INVxp67_ASAP7_75t_SL g19017 ( 
.A(n_18736),
.Y(n_19017)
);

INVx1_ASAP7_75t_L g19018 ( 
.A(n_18514),
.Y(n_19018)
);

NAND2xp5_ASAP7_75t_L g19019 ( 
.A(n_18714),
.B(n_10963),
.Y(n_19019)
);

NAND2xp5_ASAP7_75t_L g19020 ( 
.A(n_18757),
.B(n_10963),
.Y(n_19020)
);

AOI22xp5_ASAP7_75t_L g19021 ( 
.A1(n_18614),
.A2(n_10110),
.B1(n_10181),
.B2(n_11341),
.Y(n_19021)
);

HB1xp67_ASAP7_75t_L g19022 ( 
.A(n_18568),
.Y(n_19022)
);

INVx1_ASAP7_75t_L g19023 ( 
.A(n_18474),
.Y(n_19023)
);

NAND2x1p5_ASAP7_75t_L g19024 ( 
.A(n_18690),
.B(n_9636),
.Y(n_19024)
);

NAND2xp5_ASAP7_75t_L g19025 ( 
.A(n_18744),
.B(n_10963),
.Y(n_19025)
);

NAND2xp5_ASAP7_75t_L g19026 ( 
.A(n_18616),
.B(n_10963),
.Y(n_19026)
);

NAND2xp5_ASAP7_75t_L g19027 ( 
.A(n_18618),
.B(n_10963),
.Y(n_19027)
);

AND2x2_ASAP7_75t_L g19028 ( 
.A(n_18797),
.B(n_8638),
.Y(n_19028)
);

AOI22xp5_ASAP7_75t_L g19029 ( 
.A1(n_18601),
.A2(n_10110),
.B1(n_10181),
.B2(n_11341),
.Y(n_19029)
);

AOI22xp5_ASAP7_75t_L g19030 ( 
.A1(n_18615),
.A2(n_10110),
.B1(n_10181),
.B2(n_11341),
.Y(n_19030)
);

INVx2_ASAP7_75t_SL g19031 ( 
.A(n_18736),
.Y(n_19031)
);

INVx1_ASAP7_75t_L g19032 ( 
.A(n_18458),
.Y(n_19032)
);

INVx2_ASAP7_75t_L g19033 ( 
.A(n_18564),
.Y(n_19033)
);

INVx1_ASAP7_75t_L g19034 ( 
.A(n_18604),
.Y(n_19034)
);

INVx1_ASAP7_75t_L g19035 ( 
.A(n_18539),
.Y(n_19035)
);

NOR2xp33_ASAP7_75t_L g19036 ( 
.A(n_18620),
.B(n_18621),
.Y(n_19036)
);

AND2x4_ASAP7_75t_SL g19037 ( 
.A(n_18841),
.B(n_7782),
.Y(n_19037)
);

AND2x2_ASAP7_75t_L g19038 ( 
.A(n_18801),
.B(n_8638),
.Y(n_19038)
);

INVx1_ASAP7_75t_L g19039 ( 
.A(n_18519),
.Y(n_19039)
);

INVx2_ASAP7_75t_L g19040 ( 
.A(n_18575),
.Y(n_19040)
);

INVx2_ASAP7_75t_SL g19041 ( 
.A(n_18718),
.Y(n_19041)
);

INVx2_ASAP7_75t_L g19042 ( 
.A(n_18585),
.Y(n_19042)
);

INVx1_ASAP7_75t_L g19043 ( 
.A(n_18471),
.Y(n_19043)
);

INVx1_ASAP7_75t_L g19044 ( 
.A(n_18630),
.Y(n_19044)
);

INVx1_ASAP7_75t_L g19045 ( 
.A(n_18693),
.Y(n_19045)
);

INVx1_ASAP7_75t_L g19046 ( 
.A(n_18587),
.Y(n_19046)
);

INVxp67_ASAP7_75t_SL g19047 ( 
.A(n_18840),
.Y(n_19047)
);

A2O1A1Ixp33_ASAP7_75t_L g19048 ( 
.A1(n_18463),
.A2(n_10868),
.B(n_10871),
.C(n_10842),
.Y(n_19048)
);

OR2x2_ASAP7_75t_L g19049 ( 
.A(n_18852),
.B(n_11617),
.Y(n_19049)
);

NOR2x1_ASAP7_75t_L g19050 ( 
.A(n_18484),
.B(n_11904),
.Y(n_19050)
);

INVx1_ASAP7_75t_L g19051 ( 
.A(n_18595),
.Y(n_19051)
);

NAND2xp5_ASAP7_75t_L g19052 ( 
.A(n_18864),
.B(n_18867),
.Y(n_19052)
);

NAND2xp5_ASAP7_75t_L g19053 ( 
.A(n_18496),
.B(n_10966),
.Y(n_19053)
);

AND2x2_ASAP7_75t_L g19054 ( 
.A(n_18709),
.B(n_8638),
.Y(n_19054)
);

OR2x2_ASAP7_75t_L g19055 ( 
.A(n_18881),
.B(n_11617),
.Y(n_19055)
);

INVx1_ASAP7_75t_L g19056 ( 
.A(n_18612),
.Y(n_19056)
);

INVx1_ASAP7_75t_L g19057 ( 
.A(n_18527),
.Y(n_19057)
);

OR2x2_ASAP7_75t_L g19058 ( 
.A(n_18862),
.B(n_11617),
.Y(n_19058)
);

INVx1_ASAP7_75t_L g19059 ( 
.A(n_18529),
.Y(n_19059)
);

AND2x4_ASAP7_75t_SL g19060 ( 
.A(n_18787),
.B(n_18823),
.Y(n_19060)
);

OAI21xp33_ASAP7_75t_L g19061 ( 
.A1(n_18740),
.A2(n_10112),
.B(n_10081),
.Y(n_19061)
);

NAND2xp5_ASAP7_75t_L g19062 ( 
.A(n_18878),
.B(n_10966),
.Y(n_19062)
);

OAI32xp33_ASAP7_75t_L g19063 ( 
.A1(n_18473),
.A2(n_9843),
.A3(n_9859),
.B1(n_9809),
.B2(n_9796),
.Y(n_19063)
);

AND2x2_ASAP7_75t_L g19064 ( 
.A(n_18608),
.B(n_8638),
.Y(n_19064)
);

OR2x6_ASAP7_75t_L g19065 ( 
.A(n_18691),
.B(n_9005),
.Y(n_19065)
);

OR2x2_ASAP7_75t_L g19066 ( 
.A(n_18530),
.B(n_11617),
.Y(n_19066)
);

INVx1_ASAP7_75t_SL g19067 ( 
.A(n_18491),
.Y(n_19067)
);

AND2x2_ASAP7_75t_L g19068 ( 
.A(n_18742),
.B(n_8681),
.Y(n_19068)
);

NAND2xp5_ASAP7_75t_L g19069 ( 
.A(n_18627),
.B(n_10966),
.Y(n_19069)
);

OR2x2_ASAP7_75t_L g19070 ( 
.A(n_18583),
.B(n_11617),
.Y(n_19070)
);

OR2x2_ASAP7_75t_L g19071 ( 
.A(n_18597),
.B(n_11617),
.Y(n_19071)
);

INVx2_ASAP7_75t_L g19072 ( 
.A(n_18658),
.Y(n_19072)
);

AND2x2_ASAP7_75t_L g19073 ( 
.A(n_18745),
.B(n_8681),
.Y(n_19073)
);

INVx1_ASAP7_75t_L g19074 ( 
.A(n_18869),
.Y(n_19074)
);

INVx1_ASAP7_75t_L g19075 ( 
.A(n_18901),
.Y(n_19075)
);

INVx2_ASAP7_75t_L g19076 ( 
.A(n_18652),
.Y(n_19076)
);

AND2x2_ASAP7_75t_L g19077 ( 
.A(n_18761),
.B(n_8681),
.Y(n_19077)
);

NAND2xp5_ASAP7_75t_L g19078 ( 
.A(n_18649),
.B(n_10966),
.Y(n_19078)
);

NAND2xp5_ASAP7_75t_L g19079 ( 
.A(n_18760),
.B(n_10966),
.Y(n_19079)
);

INVx1_ASAP7_75t_L g19080 ( 
.A(n_18553),
.Y(n_19080)
);

NOR2xp33_ASAP7_75t_L g19081 ( 
.A(n_18559),
.B(n_7996),
.Y(n_19081)
);

INVx1_ASAP7_75t_L g19082 ( 
.A(n_18569),
.Y(n_19082)
);

INVxp67_ASAP7_75t_L g19083 ( 
.A(n_18549),
.Y(n_19083)
);

NAND2xp5_ASAP7_75t_SL g19084 ( 
.A(n_18540),
.B(n_10181),
.Y(n_19084)
);

OR2x2_ASAP7_75t_L g19085 ( 
.A(n_18571),
.B(n_10531),
.Y(n_19085)
);

AND2x2_ASAP7_75t_L g19086 ( 
.A(n_18771),
.B(n_8681),
.Y(n_19086)
);

AND2x2_ASAP7_75t_L g19087 ( 
.A(n_18494),
.B(n_8687),
.Y(n_19087)
);

INVx1_ASAP7_75t_L g19088 ( 
.A(n_18573),
.Y(n_19088)
);

INVxp67_ASAP7_75t_SL g19089 ( 
.A(n_18814),
.Y(n_19089)
);

NAND2xp5_ASAP7_75t_L g19090 ( 
.A(n_18734),
.B(n_10966),
.Y(n_19090)
);

NAND2xp5_ASAP7_75t_L g19091 ( 
.A(n_18609),
.B(n_11423),
.Y(n_19091)
);

NAND2xp5_ASAP7_75t_L g19092 ( 
.A(n_18579),
.B(n_11423),
.Y(n_19092)
);

INVx1_ASAP7_75t_L g19093 ( 
.A(n_18858),
.Y(n_19093)
);

AND2x2_ASAP7_75t_L g19094 ( 
.A(n_18521),
.B(n_8687),
.Y(n_19094)
);

INVx1_ASAP7_75t_L g19095 ( 
.A(n_18455),
.Y(n_19095)
);

INVx1_ASAP7_75t_L g19096 ( 
.A(n_18525),
.Y(n_19096)
);

OAI21xp33_ASAP7_75t_L g19097 ( 
.A1(n_18754),
.A2(n_10112),
.B(n_10081),
.Y(n_19097)
);

AND2x2_ASAP7_75t_L g19098 ( 
.A(n_18717),
.B(n_8687),
.Y(n_19098)
);

INVx1_ASAP7_75t_L g19099 ( 
.A(n_18593),
.Y(n_19099)
);

INVx1_ASAP7_75t_L g19100 ( 
.A(n_18576),
.Y(n_19100)
);

OAI211xp5_ASAP7_75t_L g19101 ( 
.A1(n_18493),
.A2(n_11904),
.B(n_9675),
.C(n_9848),
.Y(n_19101)
);

OR2x2_ASAP7_75t_L g19102 ( 
.A(n_18642),
.B(n_10531),
.Y(n_19102)
);

INVx2_ASAP7_75t_L g19103 ( 
.A(n_18647),
.Y(n_19103)
);

BUFx2_ASAP7_75t_L g19104 ( 
.A(n_18735),
.Y(n_19104)
);

OR2x2_ASAP7_75t_L g19105 ( 
.A(n_18657),
.B(n_10531),
.Y(n_19105)
);

AND2x2_ASAP7_75t_L g19106 ( 
.A(n_18592),
.B(n_8687),
.Y(n_19106)
);

AND2x2_ASAP7_75t_L g19107 ( 
.A(n_18726),
.B(n_9785),
.Y(n_19107)
);

NAND2xp5_ASAP7_75t_L g19108 ( 
.A(n_18581),
.B(n_11429),
.Y(n_19108)
);

OR2x2_ASAP7_75t_L g19109 ( 
.A(n_18631),
.B(n_10531),
.Y(n_19109)
);

OAI21xp33_ASAP7_75t_L g19110 ( 
.A1(n_18664),
.A2(n_10112),
.B(n_10081),
.Y(n_19110)
);

INVx1_ASAP7_75t_L g19111 ( 
.A(n_18507),
.Y(n_19111)
);

INVx2_ASAP7_75t_L g19112 ( 
.A(n_18759),
.Y(n_19112)
);

INVx1_ASAP7_75t_L g19113 ( 
.A(n_18546),
.Y(n_19113)
);

INVxp67_ASAP7_75t_SL g19114 ( 
.A(n_18544),
.Y(n_19114)
);

AND2x2_ASAP7_75t_L g19115 ( 
.A(n_18598),
.B(n_9785),
.Y(n_19115)
);

OAI22xp5_ASAP7_75t_L g19116 ( 
.A1(n_18622),
.A2(n_10181),
.B1(n_9809),
.B2(n_9843),
.Y(n_19116)
);

INVx1_ASAP7_75t_L g19117 ( 
.A(n_18547),
.Y(n_19117)
);

AND2x2_ASAP7_75t_L g19118 ( 
.A(n_18611),
.B(n_9785),
.Y(n_19118)
);

INVx2_ASAP7_75t_L g19119 ( 
.A(n_18668),
.Y(n_19119)
);

OAI32xp33_ASAP7_75t_L g19120 ( 
.A1(n_18503),
.A2(n_9862),
.A3(n_9864),
.B1(n_9859),
.B2(n_9796),
.Y(n_19120)
);

AND2x2_ASAP7_75t_L g19121 ( 
.A(n_18863),
.B(n_9827),
.Y(n_19121)
);

INVx1_ASAP7_75t_SL g19122 ( 
.A(n_18793),
.Y(n_19122)
);

AND2x4_ASAP7_75t_L g19123 ( 
.A(n_18551),
.B(n_11293),
.Y(n_19123)
);

OAI21xp5_ASAP7_75t_SL g19124 ( 
.A1(n_18537),
.A2(n_18586),
.B(n_18703),
.Y(n_19124)
);

INVx2_ASAP7_75t_L g19125 ( 
.A(n_18656),
.Y(n_19125)
);

NAND2xp5_ASAP7_75t_L g19126 ( 
.A(n_18449),
.B(n_11429),
.Y(n_19126)
);

AND2x2_ASAP7_75t_L g19127 ( 
.A(n_18650),
.B(n_9827),
.Y(n_19127)
);

INVx2_ASAP7_75t_L g19128 ( 
.A(n_18743),
.Y(n_19128)
);

NAND2xp5_ASAP7_75t_L g19129 ( 
.A(n_18669),
.B(n_11441),
.Y(n_19129)
);

NAND3xp33_ASAP7_75t_L g19130 ( 
.A(n_18641),
.B(n_10026),
.C(n_10007),
.Y(n_19130)
);

INVx1_ASAP7_75t_L g19131 ( 
.A(n_18550),
.Y(n_19131)
);

INVx1_ASAP7_75t_L g19132 ( 
.A(n_18554),
.Y(n_19132)
);

HB1xp67_ASAP7_75t_L g19133 ( 
.A(n_18696),
.Y(n_19133)
);

OAI21xp33_ASAP7_75t_SL g19134 ( 
.A1(n_18518),
.A2(n_10868),
.B(n_10871),
.Y(n_19134)
);

INVx1_ASAP7_75t_L g19135 ( 
.A(n_18555),
.Y(n_19135)
);

INVx2_ASAP7_75t_SL g19136 ( 
.A(n_18638),
.Y(n_19136)
);

NAND2xp5_ASAP7_75t_L g19137 ( 
.A(n_18748),
.B(n_11441),
.Y(n_19137)
);

INVxp67_ASAP7_75t_L g19138 ( 
.A(n_18541),
.Y(n_19138)
);

HB1xp67_ASAP7_75t_L g19139 ( 
.A(n_18535),
.Y(n_19139)
);

NAND2xp5_ASAP7_75t_L g19140 ( 
.A(n_18750),
.B(n_11445),
.Y(n_19140)
);

NAND2xp5_ASAP7_75t_L g19141 ( 
.A(n_18753),
.B(n_11445),
.Y(n_19141)
);

NOR2x1_ASAP7_75t_L g19142 ( 
.A(n_18645),
.B(n_12887),
.Y(n_19142)
);

INVx1_ASAP7_75t_L g19143 ( 
.A(n_18557),
.Y(n_19143)
);

AND2x4_ASAP7_75t_L g19144 ( 
.A(n_18763),
.B(n_10081),
.Y(n_19144)
);

AND2x2_ASAP7_75t_L g19145 ( 
.A(n_18650),
.B(n_9827),
.Y(n_19145)
);

INVx1_ASAP7_75t_L g19146 ( 
.A(n_18561),
.Y(n_19146)
);

AND2x2_ASAP7_75t_L g19147 ( 
.A(n_18670),
.B(n_9827),
.Y(n_19147)
);

NAND2xp5_ASAP7_75t_L g19148 ( 
.A(n_18674),
.B(n_11450),
.Y(n_19148)
);

AND2x2_ASAP7_75t_L g19149 ( 
.A(n_18686),
.B(n_9827),
.Y(n_19149)
);

AND2x4_ASAP7_75t_L g19150 ( 
.A(n_18662),
.B(n_11293),
.Y(n_19150)
);

AND2x2_ASAP7_75t_L g19151 ( 
.A(n_18692),
.B(n_9827),
.Y(n_19151)
);

INVx2_ASAP7_75t_L g19152 ( 
.A(n_18574),
.Y(n_19152)
);

INVx1_ASAP7_75t_L g19153 ( 
.A(n_18578),
.Y(n_19153)
);

AND2x2_ASAP7_75t_L g19154 ( 
.A(n_18700),
.B(n_9827),
.Y(n_19154)
);

AND2x2_ASAP7_75t_L g19155 ( 
.A(n_18710),
.B(n_9827),
.Y(n_19155)
);

INVx1_ASAP7_75t_L g19156 ( 
.A(n_18589),
.Y(n_19156)
);

NAND2xp5_ASAP7_75t_L g19157 ( 
.A(n_18778),
.B(n_11450),
.Y(n_19157)
);

AOI22xp5_ASAP7_75t_L g19158 ( 
.A1(n_18719),
.A2(n_10181),
.B1(n_11358),
.B2(n_11341),
.Y(n_19158)
);

AND2x2_ASAP7_75t_L g19159 ( 
.A(n_18707),
.B(n_9827),
.Y(n_19159)
);

NAND2xp5_ASAP7_75t_L g19160 ( 
.A(n_18666),
.B(n_11451),
.Y(n_19160)
);

INVxp67_ASAP7_75t_L g19161 ( 
.A(n_18506),
.Y(n_19161)
);

INVx1_ASAP7_75t_L g19162 ( 
.A(n_18552),
.Y(n_19162)
);

INVxp33_ASAP7_75t_L g19163 ( 
.A(n_18790),
.Y(n_19163)
);

INVx1_ASAP7_75t_L g19164 ( 
.A(n_18524),
.Y(n_19164)
);

NAND2xp5_ASAP7_75t_L g19165 ( 
.A(n_18722),
.B(n_11451),
.Y(n_19165)
);

NAND2xp5_ASAP7_75t_L g19166 ( 
.A(n_18725),
.B(n_11454),
.Y(n_19166)
);

AND2x2_ASAP7_75t_L g19167 ( 
.A(n_18818),
.B(n_18536),
.Y(n_19167)
);

AND2x2_ASAP7_75t_L g19168 ( 
.A(n_18538),
.B(n_9829),
.Y(n_19168)
);

INVx1_ASAP7_75t_SL g19169 ( 
.A(n_18599),
.Y(n_19169)
);

OR2x2_ASAP7_75t_L g19170 ( 
.A(n_18485),
.B(n_10531),
.Y(n_19170)
);

INVx1_ASAP7_75t_SL g19171 ( 
.A(n_18628),
.Y(n_19171)
);

AND2x2_ASAP7_75t_L g19172 ( 
.A(n_18756),
.B(n_9829),
.Y(n_19172)
);

A2O1A1Ixp33_ASAP7_75t_L g19173 ( 
.A1(n_18847),
.A2(n_10842),
.B(n_10856),
.C(n_10852),
.Y(n_19173)
);

INVx1_ASAP7_75t_L g19174 ( 
.A(n_18570),
.Y(n_19174)
);

INVx1_ASAP7_75t_L g19175 ( 
.A(n_18523),
.Y(n_19175)
);

AOI21xp33_ASAP7_75t_SL g19176 ( 
.A1(n_18772),
.A2(n_10047),
.B(n_10011),
.Y(n_19176)
);

AND2x2_ASAP7_75t_L g19177 ( 
.A(n_18526),
.B(n_9829),
.Y(n_19177)
);

AND2x2_ASAP7_75t_L g19178 ( 
.A(n_18735),
.B(n_9829),
.Y(n_19178)
);

AND2x2_ASAP7_75t_L g19179 ( 
.A(n_18533),
.B(n_9829),
.Y(n_19179)
);

INVx1_ASAP7_75t_SL g19180 ( 
.A(n_18625),
.Y(n_19180)
);

OAI21xp5_ASAP7_75t_L g19181 ( 
.A1(n_18904),
.A2(n_10668),
.B(n_10679),
.Y(n_19181)
);

INVx1_ASAP7_75t_L g19182 ( 
.A(n_18792),
.Y(n_19182)
);

NOR2xp67_ASAP7_75t_L g19183 ( 
.A(n_18635),
.B(n_11293),
.Y(n_19183)
);

BUFx2_ASAP7_75t_L g19184 ( 
.A(n_18900),
.Y(n_19184)
);

AND2x2_ASAP7_75t_L g19185 ( 
.A(n_18520),
.B(n_9829),
.Y(n_19185)
);

NAND2xp5_ASAP7_75t_L g19186 ( 
.A(n_18728),
.B(n_11454),
.Y(n_19186)
);

INVx1_ASAP7_75t_L g19187 ( 
.A(n_18563),
.Y(n_19187)
);

INVx1_ASAP7_75t_L g19188 ( 
.A(n_18633),
.Y(n_19188)
);

NOR2x1_ASAP7_75t_L g19189 ( 
.A(n_18729),
.B(n_12887),
.Y(n_19189)
);

AOI22xp5_ASAP7_75t_L g19190 ( 
.A1(n_18887),
.A2(n_10181),
.B1(n_11502),
.B2(n_11358),
.Y(n_19190)
);

AND2x2_ASAP7_75t_L g19191 ( 
.A(n_18679),
.B(n_9829),
.Y(n_19191)
);

INVx1_ASAP7_75t_L g19192 ( 
.A(n_18636),
.Y(n_19192)
);

NAND2xp5_ASAP7_75t_L g19193 ( 
.A(n_18731),
.B(n_11456),
.Y(n_19193)
);

AND2x2_ASAP7_75t_L g19194 ( 
.A(n_18688),
.B(n_9829),
.Y(n_19194)
);

INVx1_ASAP7_75t_L g19195 ( 
.A(n_18637),
.Y(n_19195)
);

INVx1_ASAP7_75t_L g19196 ( 
.A(n_18676),
.Y(n_19196)
);

INVx1_ASAP7_75t_L g19197 ( 
.A(n_18678),
.Y(n_19197)
);

INVx2_ASAP7_75t_L g19198 ( 
.A(n_18781),
.Y(n_19198)
);

INVx1_ASAP7_75t_L g19199 ( 
.A(n_18681),
.Y(n_19199)
);

INVx1_ASAP7_75t_L g19200 ( 
.A(n_18687),
.Y(n_19200)
);

AND2x2_ASAP7_75t_L g19201 ( 
.A(n_18517),
.B(n_9829),
.Y(n_19201)
);

AND2x2_ASAP7_75t_L g19202 ( 
.A(n_18883),
.B(n_9858),
.Y(n_19202)
);

INVx1_ASAP7_75t_L g19203 ( 
.A(n_18746),
.Y(n_19203)
);

AND2x2_ASAP7_75t_L g19204 ( 
.A(n_18602),
.B(n_9858),
.Y(n_19204)
);

INVx1_ASAP7_75t_L g19205 ( 
.A(n_18766),
.Y(n_19205)
);

NOR2x1_ASAP7_75t_L g19206 ( 
.A(n_18768),
.B(n_18769),
.Y(n_19206)
);

INVx1_ASAP7_75t_L g19207 ( 
.A(n_18773),
.Y(n_19207)
);

INVx2_ASAP7_75t_SL g19208 ( 
.A(n_18580),
.Y(n_19208)
);

NOR2x1p5_ASAP7_75t_SL g19209 ( 
.A(n_18644),
.B(n_11305),
.Y(n_19209)
);

INVx1_ASAP7_75t_L g19210 ( 
.A(n_18780),
.Y(n_19210)
);

INVx2_ASAP7_75t_L g19211 ( 
.A(n_18783),
.Y(n_19211)
);

INVx1_ASAP7_75t_SL g19212 ( 
.A(n_18640),
.Y(n_19212)
);

AND2x2_ASAP7_75t_L g19213 ( 
.A(n_18602),
.B(n_9858),
.Y(n_19213)
);

NAND2xp5_ASAP7_75t_L g19214 ( 
.A(n_18789),
.B(n_11456),
.Y(n_19214)
);

NOR2xp33_ASAP7_75t_L g19215 ( 
.A(n_18791),
.B(n_8037),
.Y(n_19215)
);

OR2x2_ASAP7_75t_L g19216 ( 
.A(n_18865),
.B(n_10531),
.Y(n_19216)
);

INVx1_ASAP7_75t_L g19217 ( 
.A(n_18794),
.Y(n_19217)
);

INVx1_ASAP7_75t_L g19218 ( 
.A(n_18798),
.Y(n_19218)
);

INVx2_ASAP7_75t_L g19219 ( 
.A(n_18824),
.Y(n_19219)
);

INVxp67_ASAP7_75t_L g19220 ( 
.A(n_18804),
.Y(n_19220)
);

INVx2_ASAP7_75t_L g19221 ( 
.A(n_18882),
.Y(n_19221)
);

INVxp67_ASAP7_75t_L g19222 ( 
.A(n_18805),
.Y(n_19222)
);

AND2x2_ASAP7_75t_L g19223 ( 
.A(n_18653),
.B(n_18807),
.Y(n_19223)
);

NAND2xp5_ASAP7_75t_L g19224 ( 
.A(n_18809),
.B(n_11459),
.Y(n_19224)
);

NAND2xp5_ASAP7_75t_L g19225 ( 
.A(n_18817),
.B(n_11459),
.Y(n_19225)
);

INVx1_ASAP7_75t_L g19226 ( 
.A(n_18819),
.Y(n_19226)
);

NAND2xp5_ASAP7_75t_L g19227 ( 
.A(n_18826),
.B(n_11462),
.Y(n_19227)
);

INVx1_ASAP7_75t_L g19228 ( 
.A(n_18827),
.Y(n_19228)
);

NAND2xp5_ASAP7_75t_L g19229 ( 
.A(n_18884),
.B(n_11462),
.Y(n_19229)
);

INVxp67_ASAP7_75t_SL g19230 ( 
.A(n_18682),
.Y(n_19230)
);

INVx2_ASAP7_75t_L g19231 ( 
.A(n_18831),
.Y(n_19231)
);

AOI221xp5_ASAP7_75t_L g19232 ( 
.A1(n_18870),
.A2(n_9294),
.B1(n_9329),
.B2(n_9108),
.C(n_9001),
.Y(n_19232)
);

INVx2_ASAP7_75t_L g19233 ( 
.A(n_18839),
.Y(n_19233)
);

INVx1_ASAP7_75t_L g19234 ( 
.A(n_18845),
.Y(n_19234)
);

INVx1_ASAP7_75t_L g19235 ( 
.A(n_18857),
.Y(n_19235)
);

AND2x2_ASAP7_75t_L g19236 ( 
.A(n_18685),
.B(n_9858),
.Y(n_19236)
);

AND2x2_ASAP7_75t_L g19237 ( 
.A(n_18727),
.B(n_9858),
.Y(n_19237)
);

AOI22xp33_ASAP7_75t_L g19238 ( 
.A1(n_18888),
.A2(n_11169),
.B1(n_11172),
.B2(n_11157),
.Y(n_19238)
);

INVx1_ASAP7_75t_L g19239 ( 
.A(n_18868),
.Y(n_19239)
);

INVx2_ASAP7_75t_SL g19240 ( 
.A(n_18800),
.Y(n_19240)
);

OR2x2_ASAP7_75t_L g19241 ( 
.A(n_18830),
.B(n_10531),
.Y(n_19241)
);

AND2x2_ASAP7_75t_L g19242 ( 
.A(n_18738),
.B(n_9858),
.Y(n_19242)
);

NAND2xp5_ASAP7_75t_L g19243 ( 
.A(n_18829),
.B(n_11468),
.Y(n_19243)
);

AND2x2_ASAP7_75t_L g19244 ( 
.A(n_18764),
.B(n_9858),
.Y(n_19244)
);

NOR2x1_ASAP7_75t_L g19245 ( 
.A(n_18872),
.B(n_12887),
.Y(n_19245)
);

INVxp67_ASAP7_75t_L g19246 ( 
.A(n_18481),
.Y(n_19246)
);

INVx1_ASAP7_75t_L g19247 ( 
.A(n_18873),
.Y(n_19247)
);

AOI22xp5_ASAP7_75t_L g19248 ( 
.A1(n_18825),
.A2(n_11358),
.B1(n_11502),
.B2(n_10112),
.Y(n_19248)
);

AND2x2_ASAP7_75t_L g19249 ( 
.A(n_18765),
.B(n_18774),
.Y(n_19249)
);

OAI21xp33_ASAP7_75t_L g19250 ( 
.A1(n_18892),
.A2(n_10112),
.B(n_9779),
.Y(n_19250)
);

INVx1_ASAP7_75t_L g19251 ( 
.A(n_18874),
.Y(n_19251)
);

AOI22xp5_ASAP7_75t_L g19252 ( 
.A1(n_18808),
.A2(n_11502),
.B1(n_11358),
.B2(n_9077),
.Y(n_19252)
);

AND2x2_ASAP7_75t_L g19253 ( 
.A(n_18543),
.B(n_9858),
.Y(n_19253)
);

OR2x2_ASAP7_75t_L g19254 ( 
.A(n_18663),
.B(n_10238),
.Y(n_19254)
);

INVx1_ASAP7_75t_L g19255 ( 
.A(n_18877),
.Y(n_19255)
);

NAND2x1p5_ASAP7_75t_L g19256 ( 
.A(n_18834),
.B(n_9636),
.Y(n_19256)
);

INVx1_ASAP7_75t_L g19257 ( 
.A(n_18879),
.Y(n_19257)
);

AND2x2_ASAP7_75t_L g19258 ( 
.A(n_18895),
.B(n_18835),
.Y(n_19258)
);

AND2x2_ASAP7_75t_L g19259 ( 
.A(n_18837),
.B(n_9858),
.Y(n_19259)
);

NAND2xp5_ASAP7_75t_SL g19260 ( 
.A(n_18660),
.B(n_9060),
.Y(n_19260)
);

NAND2xp5_ASAP7_75t_L g19261 ( 
.A(n_18838),
.B(n_18844),
.Y(n_19261)
);

HB1xp67_ASAP7_75t_L g19262 ( 
.A(n_18900),
.Y(n_19262)
);

NAND2xp5_ASAP7_75t_L g19263 ( 
.A(n_18902),
.B(n_11468),
.Y(n_19263)
);

NOR2xp33_ASAP7_75t_L g19264 ( 
.A(n_18849),
.B(n_8037),
.Y(n_19264)
);

INVx1_ASAP7_75t_L g19265 ( 
.A(n_18889),
.Y(n_19265)
);

AND2x2_ASAP7_75t_L g19266 ( 
.A(n_18891),
.B(n_9186),
.Y(n_19266)
);

OR2x2_ASAP7_75t_L g19267 ( 
.A(n_18672),
.B(n_10238),
.Y(n_19267)
);

INVxp67_ASAP7_75t_L g19268 ( 
.A(n_18784),
.Y(n_19268)
);

INVx2_ASAP7_75t_L g19269 ( 
.A(n_18786),
.Y(n_19269)
);

INVx2_ASAP7_75t_L g19270 ( 
.A(n_18795),
.Y(n_19270)
);

AND2x2_ASAP7_75t_L g19271 ( 
.A(n_18903),
.B(n_9214),
.Y(n_19271)
);

INVx1_ASAP7_75t_L g19272 ( 
.A(n_18675),
.Y(n_19272)
);

AND2x2_ASAP7_75t_L g19273 ( 
.A(n_18859),
.B(n_9214),
.Y(n_19273)
);

NAND2xp5_ASAP7_75t_L g19274 ( 
.A(n_18866),
.B(n_11474),
.Y(n_19274)
);

AND2x4_ASAP7_75t_L g19275 ( 
.A(n_18810),
.B(n_9214),
.Y(n_19275)
);

INVx2_ASAP7_75t_L g19276 ( 
.A(n_18812),
.Y(n_19276)
);

NAND2xp5_ASAP7_75t_L g19277 ( 
.A(n_18886),
.B(n_11474),
.Y(n_19277)
);

AND2x2_ASAP7_75t_L g19278 ( 
.A(n_18813),
.B(n_9214),
.Y(n_19278)
);

NAND2xp5_ASAP7_75t_L g19279 ( 
.A(n_18854),
.B(n_11488),
.Y(n_19279)
);

AND2x2_ASAP7_75t_L g19280 ( 
.A(n_18820),
.B(n_9214),
.Y(n_19280)
);

NAND2xp5_ASAP7_75t_L g19281 ( 
.A(n_18785),
.B(n_11488),
.Y(n_19281)
);

AND2x2_ASAP7_75t_L g19282 ( 
.A(n_18822),
.B(n_9214),
.Y(n_19282)
);

INVx1_ASAP7_75t_L g19283 ( 
.A(n_18695),
.Y(n_19283)
);

OR2x2_ASAP7_75t_L g19284 ( 
.A(n_18799),
.B(n_18806),
.Y(n_19284)
);

INVx1_ASAP7_75t_SL g19285 ( 
.A(n_18720),
.Y(n_19285)
);

INVx2_ASAP7_75t_L g19286 ( 
.A(n_18846),
.Y(n_19286)
);

OR2x2_ASAP7_75t_L g19287 ( 
.A(n_18811),
.B(n_10238),
.Y(n_19287)
);

AND2x2_ASAP7_75t_L g19288 ( 
.A(n_18848),
.B(n_9214),
.Y(n_19288)
);

OR2x2_ASAP7_75t_L g19289 ( 
.A(n_18885),
.B(n_10238),
.Y(n_19289)
);

INVx1_ASAP7_75t_L g19290 ( 
.A(n_18721),
.Y(n_19290)
);

INVx1_ASAP7_75t_L g19291 ( 
.A(n_18732),
.Y(n_19291)
);

INVx1_ASAP7_75t_L g19292 ( 
.A(n_18755),
.Y(n_19292)
);

OAI21xp33_ASAP7_75t_L g19293 ( 
.A1(n_18716),
.A2(n_9779),
.B(n_9778),
.Y(n_19293)
);

AND2x2_ASAP7_75t_L g19294 ( 
.A(n_18706),
.B(n_9214),
.Y(n_19294)
);

INVx1_ASAP7_75t_SL g19295 ( 
.A(n_18683),
.Y(n_19295)
);

NAND2xp5_ASAP7_75t_L g19296 ( 
.A(n_18853),
.B(n_11501),
.Y(n_19296)
);

INVx2_ASAP7_75t_L g19297 ( 
.A(n_18788),
.Y(n_19297)
);

AND2x2_ASAP7_75t_L g19298 ( 
.A(n_18816),
.B(n_9245),
.Y(n_19298)
);

INVx2_ASAP7_75t_SL g19299 ( 
.A(n_18698),
.Y(n_19299)
);

AND2x4_ASAP7_75t_L g19300 ( 
.A(n_18832),
.B(n_11305),
.Y(n_19300)
);

INVx2_ASAP7_75t_L g19301 ( 
.A(n_18779),
.Y(n_19301)
);

INVx2_ASAP7_75t_L g19302 ( 
.A(n_18802),
.Y(n_19302)
);

NOR2xp33_ASAP7_75t_L g19303 ( 
.A(n_18899),
.B(n_8037),
.Y(n_19303)
);

OR2x2_ASAP7_75t_L g19304 ( 
.A(n_18851),
.B(n_10238),
.Y(n_19304)
);

NAND2xp5_ASAP7_75t_L g19305 ( 
.A(n_18646),
.B(n_18648),
.Y(n_19305)
);

NOR2x1_ASAP7_75t_SL g19306 ( 
.A(n_18775),
.B(n_9763),
.Y(n_19306)
);

AND2x2_ASAP7_75t_L g19307 ( 
.A(n_18861),
.B(n_9245),
.Y(n_19307)
);

NAND2x1p5_ASAP7_75t_L g19308 ( 
.A(n_18803),
.B(n_9636),
.Y(n_19308)
);

NAND2xp5_ASAP7_75t_L g19309 ( 
.A(n_18767),
.B(n_11501),
.Y(n_19309)
);

INVx2_ASAP7_75t_L g19310 ( 
.A(n_18875),
.Y(n_19310)
);

AND2x2_ASAP7_75t_L g19311 ( 
.A(n_18876),
.B(n_18880),
.Y(n_19311)
);

OR2x2_ASAP7_75t_L g19312 ( 
.A(n_18890),
.B(n_10238),
.Y(n_19312)
);

NAND2xp5_ASAP7_75t_L g19313 ( 
.A(n_18777),
.B(n_11517),
.Y(n_19313)
);

INVx1_ASAP7_75t_L g19314 ( 
.A(n_18673),
.Y(n_19314)
);

OR2x2_ASAP7_75t_L g19315 ( 
.A(n_18893),
.B(n_10238),
.Y(n_19315)
);

AND2x2_ASAP7_75t_L g19316 ( 
.A(n_18751),
.B(n_9245),
.Y(n_19316)
);

INVx1_ASAP7_75t_SL g19317 ( 
.A(n_18897),
.Y(n_19317)
);

INVx1_ASAP7_75t_L g19318 ( 
.A(n_18860),
.Y(n_19318)
);

OR2x2_ASAP7_75t_L g19319 ( 
.A(n_18833),
.B(n_10238),
.Y(n_19319)
);

NOR2xp33_ASAP7_75t_L g19320 ( 
.A(n_18733),
.B(n_8037),
.Y(n_19320)
);

INVx1_ASAP7_75t_L g19321 ( 
.A(n_18850),
.Y(n_19321)
);

OR2x2_ASAP7_75t_L g19322 ( 
.A(n_18739),
.B(n_11358),
.Y(n_19322)
);

INVx1_ASAP7_75t_L g19323 ( 
.A(n_18821),
.Y(n_19323)
);

NAND2xp5_ASAP7_75t_L g19324 ( 
.A(n_18758),
.B(n_18667),
.Y(n_19324)
);

OR2x2_ASAP7_75t_L g19325 ( 
.A(n_18762),
.B(n_11502),
.Y(n_19325)
);

OAI22xp5_ASAP7_75t_L g19326 ( 
.A1(n_18694),
.A2(n_18699),
.B1(n_18871),
.B2(n_18654),
.Y(n_19326)
);

AND2x2_ASAP7_75t_L g19327 ( 
.A(n_18689),
.B(n_9245),
.Y(n_19327)
);

INVx1_ASAP7_75t_L g19328 ( 
.A(n_18723),
.Y(n_19328)
);

AND2x2_ASAP7_75t_L g19329 ( 
.A(n_18701),
.B(n_9245),
.Y(n_19329)
);

INVx1_ASAP7_75t_L g19330 ( 
.A(n_18724),
.Y(n_19330)
);

INVx1_ASAP7_75t_L g19331 ( 
.A(n_18737),
.Y(n_19331)
);

INVx1_ASAP7_75t_L g19332 ( 
.A(n_18752),
.Y(n_19332)
);

OR2x2_ASAP7_75t_L g19333 ( 
.A(n_18715),
.B(n_11502),
.Y(n_19333)
);

INVx1_ASAP7_75t_L g19334 ( 
.A(n_18680),
.Y(n_19334)
);

INVx1_ASAP7_75t_L g19335 ( 
.A(n_18776),
.Y(n_19335)
);

INVxp67_ASAP7_75t_L g19336 ( 
.A(n_18796),
.Y(n_19336)
);

INVx1_ASAP7_75t_L g19337 ( 
.A(n_18566),
.Y(n_19337)
);

NOR2xp33_ASAP7_75t_SL g19338 ( 
.A(n_18936),
.B(n_18894),
.Y(n_19338)
);

AOI22xp5_ASAP7_75t_L g19339 ( 
.A1(n_19122),
.A2(n_18558),
.B1(n_18747),
.B2(n_18516),
.Y(n_19339)
);

INVx1_ASAP7_75t_L g19340 ( 
.A(n_19139),
.Y(n_19340)
);

A2O1A1Ixp33_ASAP7_75t_L g19341 ( 
.A1(n_18949),
.A2(n_18610),
.B(n_18480),
.C(n_18855),
.Y(n_19341)
);

INVx1_ASAP7_75t_L g19342 ( 
.A(n_18925),
.Y(n_19342)
);

AND2x2_ASAP7_75t_L g19343 ( 
.A(n_18923),
.B(n_9245),
.Y(n_19343)
);

NAND2xp5_ASAP7_75t_L g19344 ( 
.A(n_18929),
.B(n_10897),
.Y(n_19344)
);

AND2x2_ASAP7_75t_L g19345 ( 
.A(n_18919),
.B(n_9245),
.Y(n_19345)
);

INVx1_ASAP7_75t_L g19346 ( 
.A(n_18935),
.Y(n_19346)
);

INVx1_ASAP7_75t_L g19347 ( 
.A(n_18924),
.Y(n_19347)
);

OR2x2_ASAP7_75t_L g19348 ( 
.A(n_18965),
.B(n_11305),
.Y(n_19348)
);

AOI22xp5_ASAP7_75t_L g19349 ( 
.A1(n_18930),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19349)
);

AOI21xp33_ASAP7_75t_L g19350 ( 
.A1(n_18950),
.A2(n_12771),
.B(n_12772),
.Y(n_19350)
);

AND2x2_ASAP7_75t_L g19351 ( 
.A(n_19003),
.B(n_9245),
.Y(n_19351)
);

OR2x2_ASAP7_75t_L g19352 ( 
.A(n_18912),
.B(n_11325),
.Y(n_19352)
);

INVx1_ASAP7_75t_L g19353 ( 
.A(n_18938),
.Y(n_19353)
);

INVx1_ASAP7_75t_L g19354 ( 
.A(n_18931),
.Y(n_19354)
);

INVx2_ASAP7_75t_L g19355 ( 
.A(n_18948),
.Y(n_19355)
);

INVx1_ASAP7_75t_L g19356 ( 
.A(n_18933),
.Y(n_19356)
);

OAI22xp5_ASAP7_75t_L g19357 ( 
.A1(n_18951),
.A2(n_9859),
.B1(n_9862),
.B2(n_9796),
.Y(n_19357)
);

INVx1_ASAP7_75t_L g19358 ( 
.A(n_18956),
.Y(n_19358)
);

OAI222xp33_ASAP7_75t_L g19359 ( 
.A1(n_19067),
.A2(n_9329),
.B1(n_9001),
.B2(n_9387),
.C1(n_9332),
.C2(n_9108),
.Y(n_19359)
);

INVx1_ASAP7_75t_L g19360 ( 
.A(n_19060),
.Y(n_19360)
);

OAI21xp5_ASAP7_75t_L g19361 ( 
.A1(n_18960),
.A2(n_11572),
.B(n_11571),
.Y(n_19361)
);

INVx1_ASAP7_75t_L g19362 ( 
.A(n_18915),
.Y(n_19362)
);

INVx2_ASAP7_75t_L g19363 ( 
.A(n_18988),
.Y(n_19363)
);

NAND2xp5_ASAP7_75t_L g19364 ( 
.A(n_18916),
.B(n_18917),
.Y(n_19364)
);

INVx1_ASAP7_75t_SL g19365 ( 
.A(n_18988),
.Y(n_19365)
);

OAI22xp5_ASAP7_75t_L g19366 ( 
.A1(n_19089),
.A2(n_9862),
.B1(n_9864),
.B2(n_9859),
.Y(n_19366)
);

OR2x2_ASAP7_75t_L g19367 ( 
.A(n_19052),
.B(n_18953),
.Y(n_19367)
);

AND2x4_ASAP7_75t_L g19368 ( 
.A(n_18945),
.B(n_9271),
.Y(n_19368)
);

AOI22xp5_ASAP7_75t_L g19369 ( 
.A1(n_19107),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19369)
);

AND2x2_ASAP7_75t_L g19370 ( 
.A(n_18911),
.B(n_9271),
.Y(n_19370)
);

A2O1A1Ixp33_ASAP7_75t_L g19371 ( 
.A1(n_19008),
.A2(n_10842),
.B(n_10856),
.C(n_10852),
.Y(n_19371)
);

NAND2xp5_ASAP7_75t_L g19372 ( 
.A(n_18914),
.B(n_10897),
.Y(n_19372)
);

AOI21xp5_ASAP7_75t_L g19373 ( 
.A1(n_18927),
.A2(n_12771),
.B(n_12363),
.Y(n_19373)
);

INVx1_ASAP7_75t_SL g19374 ( 
.A(n_18989),
.Y(n_19374)
);

INVx1_ASAP7_75t_L g19375 ( 
.A(n_18905),
.Y(n_19375)
);

NOR2xp33_ASAP7_75t_L g19376 ( 
.A(n_19169),
.B(n_8037),
.Y(n_19376)
);

OAI22xp33_ASAP7_75t_L g19377 ( 
.A1(n_18979),
.A2(n_9862),
.B1(n_9864),
.B2(n_9859),
.Y(n_19377)
);

AND2x2_ASAP7_75t_SL g19378 ( 
.A(n_18928),
.B(n_9077),
.Y(n_19378)
);

NAND2xp5_ASAP7_75t_L g19379 ( 
.A(n_18974),
.B(n_11517),
.Y(n_19379)
);

INVx1_ASAP7_75t_L g19380 ( 
.A(n_19022),
.Y(n_19380)
);

AOI322xp5_ASAP7_75t_L g19381 ( 
.A1(n_18941),
.A2(n_9914),
.A3(n_9862),
.B1(n_9920),
.B2(n_9983),
.C1(n_9864),
.C2(n_9859),
.Y(n_19381)
);

INVx1_ASAP7_75t_L g19382 ( 
.A(n_18913),
.Y(n_19382)
);

AOI22xp5_ASAP7_75t_L g19383 ( 
.A1(n_19095),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19383)
);

NAND2xp5_ASAP7_75t_L g19384 ( 
.A(n_18969),
.B(n_11524),
.Y(n_19384)
);

INVx2_ASAP7_75t_SL g19385 ( 
.A(n_19037),
.Y(n_19385)
);

INVx1_ASAP7_75t_L g19386 ( 
.A(n_18957),
.Y(n_19386)
);

INVxp67_ASAP7_75t_L g19387 ( 
.A(n_18997),
.Y(n_19387)
);

INVx1_ASAP7_75t_L g19388 ( 
.A(n_18993),
.Y(n_19388)
);

AOI22xp5_ASAP7_75t_L g19389 ( 
.A1(n_19121),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19389)
);

AOI22xp5_ASAP7_75t_L g19390 ( 
.A1(n_19016),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19390)
);

NAND2xp5_ASAP7_75t_L g19391 ( 
.A(n_19114),
.B(n_18940),
.Y(n_19391)
);

AOI31xp33_ASAP7_75t_SL g19392 ( 
.A1(n_19246),
.A2(n_9864),
.A3(n_9914),
.B(n_9862),
.Y(n_19392)
);

NAND3x2_ASAP7_75t_L g19393 ( 
.A(n_19184),
.B(n_9008),
.C(n_8977),
.Y(n_19393)
);

AO22x2_ASAP7_75t_L g19394 ( 
.A1(n_18952),
.A2(n_10198),
.B1(n_10221),
.B2(n_10195),
.Y(n_19394)
);

AND2x2_ASAP7_75t_L g19395 ( 
.A(n_19249),
.B(n_9271),
.Y(n_19395)
);

AND2x2_ASAP7_75t_L g19396 ( 
.A(n_18986),
.B(n_9271),
.Y(n_19396)
);

OAI222xp33_ASAP7_75t_L g19397 ( 
.A1(n_19065),
.A2(n_19171),
.B1(n_19075),
.B2(n_19212),
.C1(n_19074),
.C2(n_18964),
.Y(n_19397)
);

OAI322xp33_ASAP7_75t_L g19398 ( 
.A1(n_18958),
.A2(n_9329),
.A3(n_9001),
.B1(n_9332),
.B2(n_9404),
.C1(n_9387),
.C2(n_10195),
.Y(n_19398)
);

AOI22xp5_ASAP7_75t_L g19399 ( 
.A1(n_19031),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19399)
);

INVx2_ASAP7_75t_L g19400 ( 
.A(n_18954),
.Y(n_19400)
);

AND2x2_ASAP7_75t_L g19401 ( 
.A(n_19033),
.B(n_9271),
.Y(n_19401)
);

INVx2_ASAP7_75t_SL g19402 ( 
.A(n_18954),
.Y(n_19402)
);

AOI211xp5_ASAP7_75t_L g19403 ( 
.A1(n_18959),
.A2(n_18966),
.B(n_18970),
.C(n_18972),
.Y(n_19403)
);

NAND2xp5_ASAP7_75t_L g19404 ( 
.A(n_19017),
.B(n_11524),
.Y(n_19404)
);

INVx2_ASAP7_75t_L g19405 ( 
.A(n_19028),
.Y(n_19405)
);

NAND2xp5_ASAP7_75t_L g19406 ( 
.A(n_18998),
.B(n_11530),
.Y(n_19406)
);

INVx1_ASAP7_75t_L g19407 ( 
.A(n_18963),
.Y(n_19407)
);

AND2x4_ASAP7_75t_L g19408 ( 
.A(n_19206),
.B(n_11325),
.Y(n_19408)
);

INVx1_ASAP7_75t_L g19409 ( 
.A(n_18991),
.Y(n_19409)
);

NAND2xp33_ASAP7_75t_SL g19410 ( 
.A(n_19240),
.B(n_9077),
.Y(n_19410)
);

OR2x2_ASAP7_75t_L g19411 ( 
.A(n_18907),
.B(n_19040),
.Y(n_19411)
);

AND2x2_ASAP7_75t_L g19412 ( 
.A(n_19042),
.B(n_9271),
.Y(n_19412)
);

INVx1_ASAP7_75t_L g19413 ( 
.A(n_18985),
.Y(n_19413)
);

INVx2_ASAP7_75t_L g19414 ( 
.A(n_19038),
.Y(n_19414)
);

INVx1_ASAP7_75t_L g19415 ( 
.A(n_18921),
.Y(n_19415)
);

INVx1_ASAP7_75t_L g19416 ( 
.A(n_18962),
.Y(n_19416)
);

OAI322xp33_ASAP7_75t_L g19417 ( 
.A1(n_19012),
.A2(n_9387),
.A3(n_9404),
.B1(n_9332),
.B2(n_10221),
.C1(n_10198),
.C2(n_10195),
.Y(n_19417)
);

INVx1_ASAP7_75t_SL g19418 ( 
.A(n_19104),
.Y(n_19418)
);

INVx3_ASAP7_75t_L g19419 ( 
.A(n_18920),
.Y(n_19419)
);

NAND2xp5_ASAP7_75t_L g19420 ( 
.A(n_18994),
.B(n_11530),
.Y(n_19420)
);

OAI22xp5_ASAP7_75t_L g19421 ( 
.A1(n_19045),
.A2(n_9914),
.B1(n_9920),
.B2(n_9864),
.Y(n_19421)
);

AND2x4_ASAP7_75t_L g19422 ( 
.A(n_19198),
.B(n_9271),
.Y(n_19422)
);

AND2x2_ASAP7_75t_L g19423 ( 
.A(n_19211),
.B(n_9271),
.Y(n_19423)
);

O2A1O1Ixp33_ASAP7_75t_L g19424 ( 
.A1(n_19262),
.A2(n_9652),
.B(n_9621),
.C(n_9083),
.Y(n_19424)
);

NAND2xp5_ASAP7_75t_L g19425 ( 
.A(n_19100),
.B(n_11537),
.Y(n_19425)
);

NAND2xp5_ASAP7_75t_L g19426 ( 
.A(n_18920),
.B(n_19006),
.Y(n_19426)
);

AOI22xp5_ASAP7_75t_L g19427 ( 
.A1(n_19046),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19427)
);

AOI22xp5_ASAP7_75t_L g19428 ( 
.A1(n_19221),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19428)
);

AOI22xp5_ASAP7_75t_L g19429 ( 
.A1(n_19231),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19429)
);

INVx1_ASAP7_75t_L g19430 ( 
.A(n_18922),
.Y(n_19430)
);

INVx1_ASAP7_75t_L g19431 ( 
.A(n_18908),
.Y(n_19431)
);

INVx1_ASAP7_75t_L g19432 ( 
.A(n_18909),
.Y(n_19432)
);

O2A1O1Ixp33_ASAP7_75t_L g19433 ( 
.A1(n_18978),
.A2(n_18968),
.B(n_19011),
.C(n_19043),
.Y(n_19433)
);

INVx1_ASAP7_75t_L g19434 ( 
.A(n_19219),
.Y(n_19434)
);

AOI31xp33_ASAP7_75t_L g19435 ( 
.A1(n_19047),
.A2(n_10104),
.A3(n_10131),
.B(n_10047),
.Y(n_19435)
);

INVx1_ASAP7_75t_L g19436 ( 
.A(n_19010),
.Y(n_19436)
);

NAND2xp5_ASAP7_75t_L g19437 ( 
.A(n_19233),
.B(n_11537),
.Y(n_19437)
);

OAI221xp5_ASAP7_75t_SL g19438 ( 
.A1(n_19124),
.A2(n_9404),
.B1(n_9387),
.B2(n_9332),
.C(n_9333),
.Y(n_19438)
);

INVx1_ASAP7_75t_L g19439 ( 
.A(n_18942),
.Y(n_19439)
);

NAND2xp5_ASAP7_75t_L g19440 ( 
.A(n_19119),
.B(n_11538),
.Y(n_19440)
);

INVx1_ASAP7_75t_L g19441 ( 
.A(n_18961),
.Y(n_19441)
);

INVx1_ASAP7_75t_L g19442 ( 
.A(n_18996),
.Y(n_19442)
);

A2O1A1Ixp33_ASAP7_75t_L g19443 ( 
.A1(n_19002),
.A2(n_10852),
.B(n_10856),
.C(n_11607),
.Y(n_19443)
);

AND2x2_ASAP7_75t_L g19444 ( 
.A(n_19269),
.B(n_9282),
.Y(n_19444)
);

NAND2xp5_ASAP7_75t_L g19445 ( 
.A(n_19270),
.B(n_11538),
.Y(n_19445)
);

AOI22xp33_ASAP7_75t_L g19446 ( 
.A1(n_18946),
.A2(n_11169),
.B1(n_11172),
.B2(n_11157),
.Y(n_19446)
);

INVx1_ASAP7_75t_L g19447 ( 
.A(n_19223),
.Y(n_19447)
);

INVxp67_ASAP7_75t_L g19448 ( 
.A(n_19036),
.Y(n_19448)
);

INVx1_ASAP7_75t_L g19449 ( 
.A(n_18955),
.Y(n_19449)
);

O2A1O1Ixp33_ASAP7_75t_L g19450 ( 
.A1(n_19230),
.A2(n_9652),
.B(n_9621),
.C(n_9083),
.Y(n_19450)
);

XOR2x2_ASAP7_75t_L g19451 ( 
.A(n_18947),
.B(n_10047),
.Y(n_19451)
);

NAND2xp5_ASAP7_75t_L g19452 ( 
.A(n_19276),
.B(n_11545),
.Y(n_19452)
);

INVx1_ASAP7_75t_L g19453 ( 
.A(n_19286),
.Y(n_19453)
);

OAI22xp5_ASAP7_75t_L g19454 ( 
.A1(n_18918),
.A2(n_9920),
.B1(n_9983),
.B2(n_9914),
.Y(n_19454)
);

INVxp67_ASAP7_75t_L g19455 ( 
.A(n_18937),
.Y(n_19455)
);

AOI21xp33_ASAP7_75t_L g19456 ( 
.A1(n_19163),
.A2(n_12771),
.B(n_12772),
.Y(n_19456)
);

AOI21xp33_ASAP7_75t_L g19457 ( 
.A1(n_18990),
.A2(n_12816),
.B(n_12772),
.Y(n_19457)
);

AND2x4_ASAP7_75t_L g19458 ( 
.A(n_19136),
.B(n_11325),
.Y(n_19458)
);

INVx1_ASAP7_75t_SL g19459 ( 
.A(n_19258),
.Y(n_19459)
);

INVx1_ASAP7_75t_L g19460 ( 
.A(n_18987),
.Y(n_19460)
);

INVx1_ASAP7_75t_L g19461 ( 
.A(n_19125),
.Y(n_19461)
);

AOI21xp5_ASAP7_75t_L g19462 ( 
.A1(n_19133),
.A2(n_12363),
.B(n_12816),
.Y(n_19462)
);

INVx1_ASAP7_75t_L g19463 ( 
.A(n_19000),
.Y(n_19463)
);

AOI21xp33_ASAP7_75t_SL g19464 ( 
.A1(n_19314),
.A2(n_10104),
.B(n_10047),
.Y(n_19464)
);

OAI21xp33_ASAP7_75t_L g19465 ( 
.A1(n_19087),
.A2(n_9779),
.B(n_9778),
.Y(n_19465)
);

OAI211xp5_ASAP7_75t_L g19466 ( 
.A1(n_18906),
.A2(n_9563),
.B(n_9848),
.C(n_9675),
.Y(n_19466)
);

AOI32xp33_ASAP7_75t_L g19467 ( 
.A1(n_19001),
.A2(n_9920),
.A3(n_9999),
.B1(n_9983),
.B2(n_9914),
.Y(n_19467)
);

NAND2xp5_ASAP7_75t_L g19468 ( 
.A(n_19112),
.B(n_11545),
.Y(n_19468)
);

NAND2xp5_ASAP7_75t_L g19469 ( 
.A(n_19128),
.B(n_11547),
.Y(n_19469)
);

NOR2xp33_ASAP7_75t_L g19470 ( 
.A(n_19103),
.B(n_8037),
.Y(n_19470)
);

INVx1_ASAP7_75t_L g19471 ( 
.A(n_19072),
.Y(n_19471)
);

NAND2xp5_ASAP7_75t_L g19472 ( 
.A(n_19096),
.B(n_11547),
.Y(n_19472)
);

INVx1_ASAP7_75t_L g19473 ( 
.A(n_18939),
.Y(n_19473)
);

NAND3xp33_ASAP7_75t_SL g19474 ( 
.A(n_19007),
.B(n_10104),
.C(n_10047),
.Y(n_19474)
);

NOR2xp33_ASAP7_75t_L g19475 ( 
.A(n_19034),
.B(n_8037),
.Y(n_19475)
);

NAND2xp5_ASAP7_75t_L g19476 ( 
.A(n_19098),
.B(n_11548),
.Y(n_19476)
);

INVx1_ASAP7_75t_L g19477 ( 
.A(n_18980),
.Y(n_19477)
);

AOI211x1_ASAP7_75t_SL g19478 ( 
.A1(n_19326),
.A2(n_11369),
.B(n_11364),
.C(n_9920),
.Y(n_19478)
);

NAND2xp5_ASAP7_75t_L g19479 ( 
.A(n_19041),
.B(n_11548),
.Y(n_19479)
);

INVx1_ASAP7_75t_L g19480 ( 
.A(n_18934),
.Y(n_19480)
);

OAI21xp33_ASAP7_75t_L g19481 ( 
.A1(n_19054),
.A2(n_9789),
.B(n_9784),
.Y(n_19481)
);

INVx1_ASAP7_75t_L g19482 ( 
.A(n_18932),
.Y(n_19482)
);

AOI32xp33_ASAP7_75t_L g19483 ( 
.A1(n_19202),
.A2(n_9920),
.A3(n_9999),
.B1(n_9983),
.B2(n_9914),
.Y(n_19483)
);

AOI22xp5_ASAP7_75t_L g19484 ( 
.A1(n_19093),
.A2(n_9141),
.B1(n_9361),
.B2(n_9077),
.Y(n_19484)
);

INVx1_ASAP7_75t_L g19485 ( 
.A(n_18982),
.Y(n_19485)
);

OAI22xp5_ASAP7_75t_L g19486 ( 
.A1(n_19065),
.A2(n_9999),
.B1(n_10022),
.B2(n_9983),
.Y(n_19486)
);

INVx1_ASAP7_75t_L g19487 ( 
.A(n_18943),
.Y(n_19487)
);

INVx2_ASAP7_75t_L g19488 ( 
.A(n_19068),
.Y(n_19488)
);

AND2x4_ASAP7_75t_SL g19489 ( 
.A(n_19167),
.B(n_9141),
.Y(n_19489)
);

AOI211xp5_ASAP7_75t_L g19490 ( 
.A1(n_19081),
.A2(n_9159),
.B(n_9386),
.C(n_9211),
.Y(n_19490)
);

INVx2_ASAP7_75t_SL g19491 ( 
.A(n_19144),
.Y(n_19491)
);

INVx1_ASAP7_75t_L g19492 ( 
.A(n_18973),
.Y(n_19492)
);

OR2x2_ASAP7_75t_L g19493 ( 
.A(n_19035),
.B(n_11364),
.Y(n_19493)
);

INVx3_ASAP7_75t_L g19494 ( 
.A(n_19178),
.Y(n_19494)
);

INVx1_ASAP7_75t_L g19495 ( 
.A(n_18967),
.Y(n_19495)
);

AOI22xp33_ASAP7_75t_SL g19496 ( 
.A1(n_19208),
.A2(n_9141),
.B1(n_9391),
.B2(n_9361),
.Y(n_19496)
);

AND2x2_ASAP7_75t_L g19497 ( 
.A(n_19118),
.B(n_9282),
.Y(n_19497)
);

INVx2_ASAP7_75t_L g19498 ( 
.A(n_19073),
.Y(n_19498)
);

OAI22xp5_ASAP7_75t_L g19499 ( 
.A1(n_19138),
.A2(n_9999),
.B1(n_10022),
.B2(n_9983),
.Y(n_19499)
);

NOR2xp67_ASAP7_75t_L g19500 ( 
.A(n_19162),
.B(n_11364),
.Y(n_19500)
);

NAND2xp5_ASAP7_75t_L g19501 ( 
.A(n_18975),
.B(n_11574),
.Y(n_19501)
);

INVx1_ASAP7_75t_L g19502 ( 
.A(n_18976),
.Y(n_19502)
);

AOI21xp5_ASAP7_75t_L g19503 ( 
.A1(n_19324),
.A2(n_12363),
.B(n_12816),
.Y(n_19503)
);

OAI22xp5_ASAP7_75t_L g19504 ( 
.A1(n_19220),
.A2(n_10022),
.B1(n_10029),
.B2(n_9999),
.Y(n_19504)
);

NAND3x2_ASAP7_75t_L g19505 ( 
.A(n_18910),
.B(n_9008),
.C(n_8977),
.Y(n_19505)
);

AND2x4_ASAP7_75t_L g19506 ( 
.A(n_19152),
.B(n_9282),
.Y(n_19506)
);

INVx2_ASAP7_75t_L g19507 ( 
.A(n_19077),
.Y(n_19507)
);

AND2x4_ASAP7_75t_L g19508 ( 
.A(n_19044),
.B(n_9282),
.Y(n_19508)
);

OAI22xp5_ASAP7_75t_L g19509 ( 
.A1(n_19222),
.A2(n_10022),
.B1(n_10029),
.B2(n_9999),
.Y(n_19509)
);

INVx2_ASAP7_75t_L g19510 ( 
.A(n_19086),
.Y(n_19510)
);

OR2x6_ASAP7_75t_L g19511 ( 
.A(n_18926),
.B(n_9005),
.Y(n_19511)
);

INVx1_ASAP7_75t_L g19512 ( 
.A(n_18977),
.Y(n_19512)
);

CKINVDCx5p33_ASAP7_75t_R g19513 ( 
.A(n_19023),
.Y(n_19513)
);

NAND2xp5_ASAP7_75t_L g19514 ( 
.A(n_18981),
.B(n_11574),
.Y(n_19514)
);

OAI21xp5_ASAP7_75t_L g19515 ( 
.A1(n_19083),
.A2(n_11572),
.B(n_11571),
.Y(n_19515)
);

AND2x2_ASAP7_75t_L g19516 ( 
.A(n_19191),
.B(n_9282),
.Y(n_19516)
);

INVx1_ASAP7_75t_SL g19517 ( 
.A(n_18995),
.Y(n_19517)
);

OAI21xp33_ASAP7_75t_L g19518 ( 
.A1(n_19215),
.A2(n_9789),
.B(n_9784),
.Y(n_19518)
);

AND2x2_ASAP7_75t_L g19519 ( 
.A(n_19194),
.B(n_9282),
.Y(n_19519)
);

INVx2_ASAP7_75t_L g19520 ( 
.A(n_19094),
.Y(n_19520)
);

INVx2_ASAP7_75t_L g19521 ( 
.A(n_19168),
.Y(n_19521)
);

OAI21xp33_ASAP7_75t_L g19522 ( 
.A1(n_19264),
.A2(n_9789),
.B(n_9784),
.Y(n_19522)
);

INVx1_ASAP7_75t_L g19523 ( 
.A(n_18983),
.Y(n_19523)
);

NAND2xp5_ASAP7_75t_SL g19524 ( 
.A(n_19099),
.B(n_9141),
.Y(n_19524)
);

INVx1_ASAP7_75t_SL g19525 ( 
.A(n_19013),
.Y(n_19525)
);

INVx1_ASAP7_75t_L g19526 ( 
.A(n_18992),
.Y(n_19526)
);

NAND2xp5_ASAP7_75t_L g19527 ( 
.A(n_18999),
.B(n_19174),
.Y(n_19527)
);

INVx1_ASAP7_75t_L g19528 ( 
.A(n_19039),
.Y(n_19528)
);

OAI21xp33_ASAP7_75t_SL g19529 ( 
.A1(n_19142),
.A2(n_10924),
.B(n_10672),
.Y(n_19529)
);

AND2x4_ASAP7_75t_L g19530 ( 
.A(n_19051),
.B(n_19056),
.Y(n_19530)
);

INVxp67_ASAP7_75t_L g19531 ( 
.A(n_18971),
.Y(n_19531)
);

INVx1_ASAP7_75t_L g19532 ( 
.A(n_19057),
.Y(n_19532)
);

INVx1_ASAP7_75t_L g19533 ( 
.A(n_19059),
.Y(n_19533)
);

OAI211xp5_ASAP7_75t_L g19534 ( 
.A1(n_18984),
.A2(n_9563),
.B(n_9848),
.C(n_9675),
.Y(n_19534)
);

OR2x6_ASAP7_75t_L g19535 ( 
.A(n_19080),
.B(n_9005),
.Y(n_19535)
);

INVx2_ASAP7_75t_SL g19536 ( 
.A(n_19266),
.Y(n_19536)
);

INVx1_ASAP7_75t_L g19537 ( 
.A(n_19082),
.Y(n_19537)
);

INVx1_ASAP7_75t_L g19538 ( 
.A(n_19088),
.Y(n_19538)
);

OAI22xp5_ASAP7_75t_L g19539 ( 
.A1(n_19048),
.A2(n_19234),
.B1(n_19239),
.B2(n_19235),
.Y(n_19539)
);

BUFx2_ASAP7_75t_L g19540 ( 
.A(n_19175),
.Y(n_19540)
);

NAND2x2_ASAP7_75t_L g19541 ( 
.A(n_18944),
.B(n_8442),
.Y(n_19541)
);

INVx1_ASAP7_75t_L g19542 ( 
.A(n_19005),
.Y(n_19542)
);

INVx1_ASAP7_75t_L g19543 ( 
.A(n_19009),
.Y(n_19543)
);

INVx1_ASAP7_75t_L g19544 ( 
.A(n_19018),
.Y(n_19544)
);

INVx1_ASAP7_75t_L g19545 ( 
.A(n_19032),
.Y(n_19545)
);

NAND2xp5_ASAP7_75t_L g19546 ( 
.A(n_19247),
.B(n_11582),
.Y(n_19546)
);

OAI33xp33_ASAP7_75t_L g19547 ( 
.A1(n_19251),
.A2(n_11589),
.A3(n_11592),
.B1(n_11618),
.B2(n_11582),
.B3(n_9789),
.Y(n_19547)
);

INVx2_ASAP7_75t_L g19548 ( 
.A(n_19177),
.Y(n_19548)
);

INVx1_ASAP7_75t_L g19549 ( 
.A(n_19255),
.Y(n_19549)
);

INVx1_ASAP7_75t_L g19550 ( 
.A(n_19257),
.Y(n_19550)
);

OAI21xp33_ASAP7_75t_L g19551 ( 
.A1(n_19303),
.A2(n_9784),
.B(n_9482),
.Y(n_19551)
);

OR2x2_ASAP7_75t_L g19552 ( 
.A(n_19265),
.B(n_11369),
.Y(n_19552)
);

NOR2xp33_ASAP7_75t_L g19553 ( 
.A(n_19161),
.B(n_8449),
.Y(n_19553)
);

HB1xp67_ASAP7_75t_L g19554 ( 
.A(n_19189),
.Y(n_19554)
);

NAND2xp5_ASAP7_75t_L g19555 ( 
.A(n_19196),
.B(n_11589),
.Y(n_19555)
);

OAI22xp5_ASAP7_75t_L g19556 ( 
.A1(n_19182),
.A2(n_10029),
.B1(n_10040),
.B2(n_10022),
.Y(n_19556)
);

OAI22xp33_ASAP7_75t_L g19557 ( 
.A1(n_19055),
.A2(n_10022),
.B1(n_10040),
.B2(n_10029),
.Y(n_19557)
);

INVx1_ASAP7_75t_L g19558 ( 
.A(n_19076),
.Y(n_19558)
);

NAND2xp5_ASAP7_75t_L g19559 ( 
.A(n_19197),
.B(n_11592),
.Y(n_19559)
);

INVx1_ASAP7_75t_L g19560 ( 
.A(n_19199),
.Y(n_19560)
);

INVx1_ASAP7_75t_L g19561 ( 
.A(n_19200),
.Y(n_19561)
);

INVx1_ASAP7_75t_L g19562 ( 
.A(n_19203),
.Y(n_19562)
);

AND2x2_ASAP7_75t_L g19563 ( 
.A(n_19259),
.B(n_9282),
.Y(n_19563)
);

INVx2_ASAP7_75t_SL g19564 ( 
.A(n_19271),
.Y(n_19564)
);

OR2x2_ASAP7_75t_L g19565 ( 
.A(n_19170),
.B(n_19205),
.Y(n_19565)
);

AND2x2_ASAP7_75t_L g19566 ( 
.A(n_19311),
.B(n_9282),
.Y(n_19566)
);

AOI32xp33_ASAP7_75t_L g19567 ( 
.A1(n_19320),
.A2(n_10040),
.A3(n_10067),
.B1(n_10061),
.B2(n_10029),
.Y(n_19567)
);

INVx1_ASAP7_75t_L g19568 ( 
.A(n_19207),
.Y(n_19568)
);

NAND2xp5_ASAP7_75t_L g19569 ( 
.A(n_19210),
.B(n_11618),
.Y(n_19569)
);

NAND2xp5_ASAP7_75t_L g19570 ( 
.A(n_19217),
.B(n_11169),
.Y(n_19570)
);

INVx2_ASAP7_75t_L g19571 ( 
.A(n_19300),
.Y(n_19571)
);

INVx1_ASAP7_75t_L g19572 ( 
.A(n_19218),
.Y(n_19572)
);

INVx1_ASAP7_75t_L g19573 ( 
.A(n_19226),
.Y(n_19573)
);

AND2x2_ASAP7_75t_L g19574 ( 
.A(n_19253),
.B(n_19179),
.Y(n_19574)
);

NAND2x1p5_ASAP7_75t_L g19575 ( 
.A(n_19187),
.B(n_9174),
.Y(n_19575)
);

NAND3xp33_ASAP7_75t_SL g19576 ( 
.A(n_19180),
.B(n_10131),
.C(n_10104),
.Y(n_19576)
);

OR2x2_ASAP7_75t_L g19577 ( 
.A(n_19228),
.B(n_11369),
.Y(n_19577)
);

OR2x2_ASAP7_75t_L g19578 ( 
.A(n_19058),
.B(n_11317),
.Y(n_19578)
);

NAND2xp5_ASAP7_75t_L g19579 ( 
.A(n_19164),
.B(n_11169),
.Y(n_19579)
);

INVx1_ASAP7_75t_L g19580 ( 
.A(n_19297),
.Y(n_19580)
);

NAND2xp5_ASAP7_75t_L g19581 ( 
.A(n_19111),
.B(n_11172),
.Y(n_19581)
);

A2O1A1Ixp33_ASAP7_75t_L g19582 ( 
.A1(n_19209),
.A2(n_11607),
.B(n_10863),
.C(n_10679),
.Y(n_19582)
);

INVx1_ASAP7_75t_L g19583 ( 
.A(n_19301),
.Y(n_19583)
);

INVx1_ASAP7_75t_L g19584 ( 
.A(n_19302),
.Y(n_19584)
);

OAI22xp5_ASAP7_75t_L g19585 ( 
.A1(n_19049),
.A2(n_10040),
.B1(n_10061),
.B2(n_10029),
.Y(n_19585)
);

INVxp67_ASAP7_75t_L g19586 ( 
.A(n_19113),
.Y(n_19586)
);

AND2x2_ASAP7_75t_L g19587 ( 
.A(n_19185),
.B(n_9301),
.Y(n_19587)
);

NOR2xp33_ASAP7_75t_L g19588 ( 
.A(n_19317),
.B(n_19117),
.Y(n_19588)
);

INVx1_ASAP7_75t_L g19589 ( 
.A(n_19310),
.Y(n_19589)
);

OAI22xp5_ASAP7_75t_SL g19590 ( 
.A1(n_19131),
.A2(n_10180),
.B1(n_10061),
.B2(n_10067),
.Y(n_19590)
);

INVxp67_ASAP7_75t_L g19591 ( 
.A(n_19132),
.Y(n_19591)
);

INVx1_ASAP7_75t_L g19592 ( 
.A(n_19318),
.Y(n_19592)
);

INVx1_ASAP7_75t_L g19593 ( 
.A(n_19321),
.Y(n_19593)
);

INVx1_ASAP7_75t_SL g19594 ( 
.A(n_19085),
.Y(n_19594)
);

NAND2xp5_ASAP7_75t_L g19595 ( 
.A(n_19135),
.B(n_11172),
.Y(n_19595)
);

OAI21xp33_ASAP7_75t_L g19596 ( 
.A1(n_19159),
.A2(n_19201),
.B(n_19172),
.Y(n_19596)
);

OAI21xp33_ASAP7_75t_L g19597 ( 
.A1(n_19127),
.A2(n_9482),
.B(n_9411),
.Y(n_19597)
);

NAND2xp5_ASAP7_75t_L g19598 ( 
.A(n_19143),
.B(n_11157),
.Y(n_19598)
);

INVxp67_ASAP7_75t_L g19599 ( 
.A(n_19146),
.Y(n_19599)
);

OAI322xp33_ASAP7_75t_L g19600 ( 
.A1(n_19025),
.A2(n_9404),
.A3(n_10221),
.B1(n_10347),
.B2(n_10350),
.C1(n_10198),
.C2(n_10195),
.Y(n_19600)
);

NAND2xp5_ASAP7_75t_L g19601 ( 
.A(n_19153),
.B(n_11157),
.Y(n_19601)
);

INVx1_ASAP7_75t_L g19602 ( 
.A(n_19323),
.Y(n_19602)
);

AND2x2_ASAP7_75t_L g19603 ( 
.A(n_19145),
.B(n_9301),
.Y(n_19603)
);

NAND2xp5_ASAP7_75t_L g19604 ( 
.A(n_19156),
.B(n_11157),
.Y(n_19604)
);

INVxp67_ASAP7_75t_L g19605 ( 
.A(n_19188),
.Y(n_19605)
);

NAND2xp5_ASAP7_75t_L g19606 ( 
.A(n_19285),
.B(n_11330),
.Y(n_19606)
);

INVx1_ASAP7_75t_L g19607 ( 
.A(n_19272),
.Y(n_19607)
);

INVx1_ASAP7_75t_L g19608 ( 
.A(n_19283),
.Y(n_19608)
);

AND2x2_ASAP7_75t_L g19609 ( 
.A(n_19204),
.B(n_9301),
.Y(n_19609)
);

NAND2xp5_ASAP7_75t_L g19610 ( 
.A(n_19337),
.B(n_11330),
.Y(n_19610)
);

INVx1_ASAP7_75t_L g19611 ( 
.A(n_19290),
.Y(n_19611)
);

INVxp67_ASAP7_75t_SL g19612 ( 
.A(n_19050),
.Y(n_19612)
);

OAI21xp5_ASAP7_75t_L g19613 ( 
.A1(n_19053),
.A2(n_11572),
.B(n_11571),
.Y(n_19613)
);

NAND2xp5_ASAP7_75t_L g19614 ( 
.A(n_19192),
.B(n_11330),
.Y(n_19614)
);

OR2x2_ASAP7_75t_L g19615 ( 
.A(n_19216),
.B(n_11317),
.Y(n_19615)
);

AOI22xp5_ASAP7_75t_L g19616 ( 
.A1(n_19147),
.A2(n_9391),
.B1(n_9455),
.B2(n_9361),
.Y(n_19616)
);

NAND2xp5_ASAP7_75t_L g19617 ( 
.A(n_19195),
.B(n_11330),
.Y(n_19617)
);

OR2x2_ASAP7_75t_L g19618 ( 
.A(n_19090),
.B(n_11317),
.Y(n_19618)
);

INVxp67_ASAP7_75t_L g19619 ( 
.A(n_19261),
.Y(n_19619)
);

OAI21xp5_ASAP7_75t_L g19620 ( 
.A1(n_19004),
.A2(n_11580),
.B(n_11573),
.Y(n_19620)
);

NAND2xp5_ASAP7_75t_L g19621 ( 
.A(n_19273),
.B(n_11330),
.Y(n_19621)
);

NAND2xp5_ASAP7_75t_L g19622 ( 
.A(n_19291),
.B(n_7696),
.Y(n_19622)
);

INVx2_ASAP7_75t_SL g19623 ( 
.A(n_19307),
.Y(n_19623)
);

AOI322xp5_ASAP7_75t_L g19624 ( 
.A1(n_19295),
.A2(n_10080),
.A3(n_10061),
.B1(n_10127),
.B2(n_10067),
.C1(n_10040),
.C2(n_9091),
.Y(n_19624)
);

AND2x2_ASAP7_75t_L g19625 ( 
.A(n_19213),
.B(n_9301),
.Y(n_19625)
);

INVx1_ASAP7_75t_L g19626 ( 
.A(n_19126),
.Y(n_19626)
);

OR2x2_ASAP7_75t_L g19627 ( 
.A(n_19229),
.B(n_11317),
.Y(n_19627)
);

INVx1_ASAP7_75t_L g19628 ( 
.A(n_19091),
.Y(n_19628)
);

OR2x2_ASAP7_75t_L g19629 ( 
.A(n_19105),
.B(n_19109),
.Y(n_19629)
);

AND2x2_ASAP7_75t_SL g19630 ( 
.A(n_19284),
.B(n_9361),
.Y(n_19630)
);

INVx1_ASAP7_75t_L g19631 ( 
.A(n_19092),
.Y(n_19631)
);

INVxp67_ASAP7_75t_L g19632 ( 
.A(n_19263),
.Y(n_19632)
);

OAI211xp5_ASAP7_75t_L g19633 ( 
.A1(n_19336),
.A2(n_9563),
.B(n_8992),
.C(n_10815),
.Y(n_19633)
);

INVx1_ASAP7_75t_L g19634 ( 
.A(n_19108),
.Y(n_19634)
);

INVx1_ASAP7_75t_L g19635 ( 
.A(n_19129),
.Y(n_19635)
);

INVx1_ASAP7_75t_L g19636 ( 
.A(n_19137),
.Y(n_19636)
);

AO21x1_ASAP7_75t_L g19637 ( 
.A1(n_19150),
.A2(n_10221),
.B(n_10198),
.Y(n_19637)
);

OAI22xp5_ASAP7_75t_L g19638 ( 
.A1(n_19275),
.A2(n_10061),
.B1(n_10067),
.B2(n_10040),
.Y(n_19638)
);

INVxp67_ASAP7_75t_L g19639 ( 
.A(n_19150),
.Y(n_19639)
);

NAND3xp33_ASAP7_75t_L g19640 ( 
.A(n_19268),
.B(n_10026),
.C(n_10007),
.Y(n_19640)
);

INVx1_ASAP7_75t_L g19641 ( 
.A(n_19140),
.Y(n_19641)
);

INVx1_ASAP7_75t_L g19642 ( 
.A(n_19141),
.Y(n_19642)
);

INVx1_ASAP7_75t_L g19643 ( 
.A(n_19148),
.Y(n_19643)
);

AOI21xp33_ASAP7_75t_L g19644 ( 
.A1(n_19334),
.A2(n_12110),
.B(n_12093),
.Y(n_19644)
);

INVx1_ASAP7_75t_L g19645 ( 
.A(n_19160),
.Y(n_19645)
);

OR2x2_ASAP7_75t_L g19646 ( 
.A(n_19066),
.B(n_11317),
.Y(n_19646)
);

BUFx2_ASAP7_75t_L g19647 ( 
.A(n_19024),
.Y(n_19647)
);

HB1xp67_ASAP7_75t_L g19648 ( 
.A(n_19245),
.Y(n_19648)
);

INVx1_ASAP7_75t_L g19649 ( 
.A(n_19165),
.Y(n_19649)
);

INVx2_ASAP7_75t_L g19650 ( 
.A(n_19300),
.Y(n_19650)
);

INVx2_ASAP7_75t_L g19651 ( 
.A(n_19244),
.Y(n_19651)
);

OAI21xp33_ASAP7_75t_L g19652 ( 
.A1(n_19149),
.A2(n_9482),
.B(n_9411),
.Y(n_19652)
);

INVx1_ASAP7_75t_SL g19653 ( 
.A(n_19070),
.Y(n_19653)
);

INVxp67_ASAP7_75t_L g19654 ( 
.A(n_19287),
.Y(n_19654)
);

AND2x2_ASAP7_75t_L g19655 ( 
.A(n_19064),
.B(n_9301),
.Y(n_19655)
);

AOI21xp5_ASAP7_75t_SL g19656 ( 
.A1(n_19299),
.A2(n_19306),
.B(n_19123),
.Y(n_19656)
);

AND2x2_ASAP7_75t_L g19657 ( 
.A(n_19151),
.B(n_9301),
.Y(n_19657)
);

INVx1_ASAP7_75t_L g19658 ( 
.A(n_19166),
.Y(n_19658)
);

NAND2x1p5_ASAP7_75t_L g19659 ( 
.A(n_19123),
.B(n_9636),
.Y(n_19659)
);

INVx1_ASAP7_75t_L g19660 ( 
.A(n_19186),
.Y(n_19660)
);

INVx1_ASAP7_75t_L g19661 ( 
.A(n_19193),
.Y(n_19661)
);

OR2x2_ASAP7_75t_L g19662 ( 
.A(n_19020),
.B(n_11317),
.Y(n_19662)
);

AOI22xp5_ASAP7_75t_L g19663 ( 
.A1(n_19154),
.A2(n_9455),
.B1(n_9456),
.B2(n_9391),
.Y(n_19663)
);

NAND2xp5_ASAP7_75t_L g19664 ( 
.A(n_19335),
.B(n_7696),
.Y(n_19664)
);

INVx1_ASAP7_75t_L g19665 ( 
.A(n_19214),
.Y(n_19665)
);

NAND2xp5_ASAP7_75t_L g19666 ( 
.A(n_19328),
.B(n_19330),
.Y(n_19666)
);

INVxp67_ASAP7_75t_SL g19667 ( 
.A(n_19256),
.Y(n_19667)
);

INVxp67_ASAP7_75t_SL g19668 ( 
.A(n_19308),
.Y(n_19668)
);

INVx1_ASAP7_75t_L g19669 ( 
.A(n_19224),
.Y(n_19669)
);

OAI21xp5_ASAP7_75t_L g19670 ( 
.A1(n_19260),
.A2(n_11580),
.B(n_11573),
.Y(n_19670)
);

INVx2_ASAP7_75t_L g19671 ( 
.A(n_19236),
.Y(n_19671)
);

NAND2xp5_ASAP7_75t_L g19672 ( 
.A(n_19331),
.B(n_7869),
.Y(n_19672)
);

NAND3xp33_ASAP7_75t_L g19673 ( 
.A(n_19069),
.B(n_10026),
.C(n_10007),
.Y(n_19673)
);

INVx1_ASAP7_75t_L g19674 ( 
.A(n_19225),
.Y(n_19674)
);

OAI211xp5_ASAP7_75t_SL g19675 ( 
.A1(n_19332),
.A2(n_9766),
.B(n_9717),
.C(n_9659),
.Y(n_19675)
);

INVx1_ASAP7_75t_L g19676 ( 
.A(n_19227),
.Y(n_19676)
);

AOI21xp33_ASAP7_75t_L g19677 ( 
.A1(n_19305),
.A2(n_12110),
.B(n_12093),
.Y(n_19677)
);

NOR2x1_ASAP7_75t_L g19678 ( 
.A(n_19292),
.B(n_19304),
.Y(n_19678)
);

INVx1_ASAP7_75t_L g19679 ( 
.A(n_19243),
.Y(n_19679)
);

INVxp67_ASAP7_75t_SL g19680 ( 
.A(n_19078),
.Y(n_19680)
);

A2O1A1Ixp33_ASAP7_75t_L g19681 ( 
.A1(n_19062),
.A2(n_10863),
.B(n_10679),
.C(n_11368),
.Y(n_19681)
);

INVx1_ASAP7_75t_L g19682 ( 
.A(n_19274),
.Y(n_19682)
);

OAI32xp33_ASAP7_75t_L g19683 ( 
.A1(n_19241),
.A2(n_10080),
.A3(n_10127),
.B1(n_10067),
.B2(n_10061),
.Y(n_19683)
);

OAI22xp33_ASAP7_75t_L g19684 ( 
.A1(n_19102),
.A2(n_10080),
.B1(n_10127),
.B2(n_10067),
.Y(n_19684)
);

OAI22xp33_ASAP7_75t_SL g19685 ( 
.A1(n_19071),
.A2(n_19254),
.B1(n_19267),
.B2(n_19079),
.Y(n_19685)
);

INVx1_ASAP7_75t_L g19686 ( 
.A(n_19279),
.Y(n_19686)
);

AND2x2_ASAP7_75t_L g19687 ( 
.A(n_19155),
.B(n_9301),
.Y(n_19687)
);

AOI21xp5_ASAP7_75t_L g19688 ( 
.A1(n_19015),
.A2(n_12760),
.B(n_12461),
.Y(n_19688)
);

AND2x2_ASAP7_75t_L g19689 ( 
.A(n_19237),
.B(n_9301),
.Y(n_19689)
);

INVx1_ASAP7_75t_L g19690 ( 
.A(n_19277),
.Y(n_19690)
);

AOI221xp5_ASAP7_75t_L g19691 ( 
.A1(n_19019),
.A2(n_9652),
.B1(n_9621),
.B2(n_9595),
.C(n_9578),
.Y(n_19691)
);

OAI22xp5_ASAP7_75t_L g19692 ( 
.A1(n_19021),
.A2(n_10127),
.B1(n_10080),
.B2(n_8977),
.Y(n_19692)
);

INVx1_ASAP7_75t_SL g19693 ( 
.A(n_19289),
.Y(n_19693)
);

INVx1_ASAP7_75t_L g19694 ( 
.A(n_19296),
.Y(n_19694)
);

OAI22xp5_ASAP7_75t_L g19695 ( 
.A1(n_19029),
.A2(n_10127),
.B1(n_10080),
.B2(n_9075),
.Y(n_19695)
);

NAND3xp33_ASAP7_75t_L g19696 ( 
.A(n_19026),
.B(n_10026),
.C(n_10007),
.Y(n_19696)
);

INVx2_ASAP7_75t_L g19697 ( 
.A(n_19242),
.Y(n_19697)
);

AND2x2_ASAP7_75t_L g19698 ( 
.A(n_19106),
.B(n_19115),
.Y(n_19698)
);

INVx1_ASAP7_75t_SL g19699 ( 
.A(n_19312),
.Y(n_19699)
);

INVx2_ASAP7_75t_L g19700 ( 
.A(n_19278),
.Y(n_19700)
);

INVx1_ASAP7_75t_L g19701 ( 
.A(n_19281),
.Y(n_19701)
);

OAI21xp5_ASAP7_75t_L g19702 ( 
.A1(n_19027),
.A2(n_11580),
.B(n_11573),
.Y(n_19702)
);

INVx1_ASAP7_75t_L g19703 ( 
.A(n_19315),
.Y(n_19703)
);

OR2x6_ASAP7_75t_L g19704 ( 
.A(n_19363),
.B(n_19402),
.Y(n_19704)
);

INVx2_ASAP7_75t_L g19705 ( 
.A(n_19419),
.Y(n_19705)
);

INVx2_ASAP7_75t_L g19706 ( 
.A(n_19400),
.Y(n_19706)
);

INVx2_ASAP7_75t_L g19707 ( 
.A(n_19365),
.Y(n_19707)
);

OAI221xp5_ASAP7_75t_L g19708 ( 
.A1(n_19338),
.A2(n_19319),
.B1(n_19097),
.B2(n_19061),
.C(n_19110),
.Y(n_19708)
);

OR2x2_ASAP7_75t_L g19709 ( 
.A(n_19459),
.B(n_19316),
.Y(n_19709)
);

AOI22xp5_ASAP7_75t_L g19710 ( 
.A1(n_19418),
.A2(n_19327),
.B1(n_19298),
.B2(n_19294),
.Y(n_19710)
);

INVx1_ASAP7_75t_L g19711 ( 
.A(n_19648),
.Y(n_19711)
);

INVx1_ASAP7_75t_L g19712 ( 
.A(n_19554),
.Y(n_19712)
);

INVx1_ASAP7_75t_L g19713 ( 
.A(n_19360),
.Y(n_19713)
);

NOR2x1_ASAP7_75t_L g19714 ( 
.A(n_19388),
.B(n_19183),
.Y(n_19714)
);

INVx1_ASAP7_75t_L g19715 ( 
.A(n_19571),
.Y(n_19715)
);

INVx1_ASAP7_75t_L g19716 ( 
.A(n_19650),
.Y(n_19716)
);

OAI32xp33_ASAP7_75t_L g19717 ( 
.A1(n_19541),
.A2(n_19309),
.A3(n_19313),
.B1(n_19325),
.B2(n_19322),
.Y(n_19717)
);

INVx1_ASAP7_75t_L g19718 ( 
.A(n_19380),
.Y(n_19718)
);

OAI221xp5_ASAP7_75t_L g19719 ( 
.A1(n_19403),
.A2(n_19293),
.B1(n_19250),
.B2(n_19134),
.C(n_19333),
.Y(n_19719)
);

AOI21xp33_ASAP7_75t_SL g19720 ( 
.A1(n_19441),
.A2(n_19084),
.B(n_19116),
.Y(n_19720)
);

NAND2xp5_ASAP7_75t_L g19721 ( 
.A(n_19416),
.B(n_19280),
.Y(n_19721)
);

INVx1_ASAP7_75t_L g19722 ( 
.A(n_19342),
.Y(n_19722)
);

INVxp67_ASAP7_75t_L g19723 ( 
.A(n_19540),
.Y(n_19723)
);

INVx1_ASAP7_75t_SL g19724 ( 
.A(n_19378),
.Y(n_19724)
);

NAND2xp5_ASAP7_75t_L g19725 ( 
.A(n_19447),
.B(n_19282),
.Y(n_19725)
);

INVx1_ASAP7_75t_L g19726 ( 
.A(n_19612),
.Y(n_19726)
);

INVx2_ASAP7_75t_L g19727 ( 
.A(n_19408),
.Y(n_19727)
);

OAI22xp5_ASAP7_75t_L g19728 ( 
.A1(n_19387),
.A2(n_19130),
.B1(n_19030),
.B2(n_19014),
.Y(n_19728)
);

AOI322xp5_ASAP7_75t_L g19729 ( 
.A1(n_19525),
.A2(n_19288),
.A3(n_19329),
.B1(n_19157),
.B2(n_19238),
.C1(n_19232),
.C2(n_19158),
.Y(n_19729)
);

INVx1_ASAP7_75t_L g19730 ( 
.A(n_19460),
.Y(n_19730)
);

AOI221xp5_ASAP7_75t_L g19731 ( 
.A1(n_19397),
.A2(n_19176),
.B1(n_19120),
.B2(n_19063),
.C(n_19181),
.Y(n_19731)
);

O2A1O1Ixp33_ASAP7_75t_L g19732 ( 
.A1(n_19415),
.A2(n_19173),
.B(n_19101),
.C(n_9083),
.Y(n_19732)
);

AOI22xp5_ASAP7_75t_L g19733 ( 
.A1(n_19374),
.A2(n_19248),
.B1(n_19190),
.B2(n_19252),
.Y(n_19733)
);

INVxp67_ASAP7_75t_L g19734 ( 
.A(n_19502),
.Y(n_19734)
);

OAI32xp33_ASAP7_75t_L g19735 ( 
.A1(n_19347),
.A2(n_19354),
.A3(n_19358),
.B1(n_19356),
.B2(n_19434),
.Y(n_19735)
);

AOI21xp5_ASAP7_75t_L g19736 ( 
.A1(n_19656),
.A2(n_12760),
.B(n_12461),
.Y(n_19736)
);

AOI21xp33_ASAP7_75t_L g19737 ( 
.A1(n_19433),
.A2(n_12274),
.B(n_12367),
.Y(n_19737)
);

AOI21xp5_ASAP7_75t_L g19738 ( 
.A1(n_19391),
.A2(n_12760),
.B(n_12461),
.Y(n_19738)
);

INVx1_ASAP7_75t_L g19739 ( 
.A(n_19411),
.Y(n_19739)
);

OR2x2_ASAP7_75t_L g19740 ( 
.A(n_19517),
.B(n_12343),
.Y(n_19740)
);

AOI22xp33_ASAP7_75t_L g19741 ( 
.A1(n_19386),
.A2(n_10039),
.B1(n_10055),
.B2(n_10026),
.Y(n_19741)
);

INVx1_ASAP7_75t_L g19742 ( 
.A(n_19340),
.Y(n_19742)
);

INVx1_ASAP7_75t_L g19743 ( 
.A(n_19492),
.Y(n_19743)
);

INVx2_ASAP7_75t_L g19744 ( 
.A(n_19408),
.Y(n_19744)
);

OAI21xp5_ASAP7_75t_L g19745 ( 
.A1(n_19341),
.A2(n_11595),
.B(n_11583),
.Y(n_19745)
);

OAI221xp5_ASAP7_75t_SL g19746 ( 
.A1(n_19339),
.A2(n_9377),
.B1(n_9333),
.B2(n_10127),
.C(n_10080),
.Y(n_19746)
);

NAND2xp5_ASAP7_75t_L g19747 ( 
.A(n_19494),
.B(n_10039),
.Y(n_19747)
);

INVxp33_ASAP7_75t_L g19748 ( 
.A(n_19376),
.Y(n_19748)
);

OAI322xp33_ASAP7_75t_L g19749 ( 
.A1(n_19353),
.A2(n_10359),
.A3(n_10350),
.B1(n_10372),
.B2(n_10389),
.C1(n_10353),
.C2(n_10347),
.Y(n_19749)
);

AOI221xp5_ASAP7_75t_L g19750 ( 
.A1(n_19539),
.A2(n_10353),
.B1(n_10359),
.B2(n_10350),
.C(n_10347),
.Y(n_19750)
);

AOI322xp5_ASAP7_75t_L g19751 ( 
.A1(n_19453),
.A2(n_9091),
.A3(n_9013),
.B1(n_9093),
.B2(n_9189),
.C1(n_9078),
.C2(n_9075),
.Y(n_19751)
);

NAND4xp25_ASAP7_75t_L g19752 ( 
.A(n_19553),
.B(n_8020),
.C(n_8460),
.D(n_8088),
.Y(n_19752)
);

OAI21xp33_ASAP7_75t_L g19753 ( 
.A1(n_19596),
.A2(n_9562),
.B(n_9559),
.Y(n_19753)
);

INVx1_ASAP7_75t_L g19754 ( 
.A(n_19439),
.Y(n_19754)
);

INVx2_ASAP7_75t_SL g19755 ( 
.A(n_19489),
.Y(n_19755)
);

NAND2xp5_ASAP7_75t_L g19756 ( 
.A(n_19482),
.B(n_19449),
.Y(n_19756)
);

AOI21xp33_ASAP7_75t_L g19757 ( 
.A1(n_19461),
.A2(n_12274),
.B(n_12367),
.Y(n_19757)
);

NOR2xp67_ASAP7_75t_SL g19758 ( 
.A(n_19485),
.B(n_19367),
.Y(n_19758)
);

AOI21xp5_ASAP7_75t_L g19759 ( 
.A1(n_19426),
.A2(n_12471),
.B(n_12451),
.Y(n_19759)
);

INVx1_ASAP7_75t_L g19760 ( 
.A(n_19364),
.Y(n_19760)
);

INVx1_ASAP7_75t_L g19761 ( 
.A(n_19574),
.Y(n_19761)
);

INVx1_ASAP7_75t_L g19762 ( 
.A(n_19698),
.Y(n_19762)
);

NOR2x1_ASAP7_75t_L g19763 ( 
.A(n_19436),
.B(n_10180),
.Y(n_19763)
);

NOR2xp67_ASAP7_75t_L g19764 ( 
.A(n_19639),
.B(n_10815),
.Y(n_19764)
);

INVx1_ASAP7_75t_L g19765 ( 
.A(n_19405),
.Y(n_19765)
);

AOI21xp33_ASAP7_75t_L g19766 ( 
.A1(n_19413),
.A2(n_12274),
.B(n_12367),
.Y(n_19766)
);

OAI22xp5_ASAP7_75t_L g19767 ( 
.A1(n_19531),
.A2(n_19455),
.B1(n_19448),
.B2(n_19393),
.Y(n_19767)
);

A2O1A1Ixp33_ASAP7_75t_L g19768 ( 
.A1(n_19470),
.A2(n_10863),
.B(n_11379),
.C(n_11368),
.Y(n_19768)
);

OAI21xp5_ASAP7_75t_L g19769 ( 
.A1(n_19619),
.A2(n_11595),
.B(n_11583),
.Y(n_19769)
);

OR2x2_ASAP7_75t_L g19770 ( 
.A(n_19651),
.B(n_12343),
.Y(n_19770)
);

INVx1_ASAP7_75t_L g19771 ( 
.A(n_19671),
.Y(n_19771)
);

HB1xp67_ASAP7_75t_L g19772 ( 
.A(n_19500),
.Y(n_19772)
);

INVx1_ASAP7_75t_L g19773 ( 
.A(n_19697),
.Y(n_19773)
);

AND2x2_ASAP7_75t_L g19774 ( 
.A(n_19521),
.B(n_9345),
.Y(n_19774)
);

INVx1_ASAP7_75t_L g19775 ( 
.A(n_19548),
.Y(n_19775)
);

INVx1_ASAP7_75t_L g19776 ( 
.A(n_19362),
.Y(n_19776)
);

AOI22xp33_ASAP7_75t_SL g19777 ( 
.A1(n_19375),
.A2(n_9455),
.B1(n_9456),
.B2(n_9391),
.Y(n_19777)
);

AND2x2_ASAP7_75t_L g19778 ( 
.A(n_19520),
.B(n_9345),
.Y(n_19778)
);

NAND2xp5_ASAP7_75t_L g19779 ( 
.A(n_19368),
.B(n_10039),
.Y(n_19779)
);

NAND2xp5_ASAP7_75t_L g19780 ( 
.A(n_19370),
.B(n_10039),
.Y(n_19780)
);

NAND2xp5_ASAP7_75t_L g19781 ( 
.A(n_19491),
.B(n_10039),
.Y(n_19781)
);

INVx1_ASAP7_75t_L g19782 ( 
.A(n_19471),
.Y(n_19782)
);

INVx3_ASAP7_75t_L g19783 ( 
.A(n_19458),
.Y(n_19783)
);

NAND2xp5_ASAP7_75t_L g19784 ( 
.A(n_19536),
.B(n_10039),
.Y(n_19784)
);

INVx2_ASAP7_75t_L g19785 ( 
.A(n_19345),
.Y(n_19785)
);

NAND2xp5_ASAP7_75t_L g19786 ( 
.A(n_19564),
.B(n_10039),
.Y(n_19786)
);

INVx1_ASAP7_75t_L g19787 ( 
.A(n_19512),
.Y(n_19787)
);

INVx1_ASAP7_75t_L g19788 ( 
.A(n_19558),
.Y(n_19788)
);

AOI22xp33_ASAP7_75t_SL g19789 ( 
.A1(n_19580),
.A2(n_9455),
.B1(n_9456),
.B2(n_9391),
.Y(n_19789)
);

INVx1_ASAP7_75t_L g19790 ( 
.A(n_19527),
.Y(n_19790)
);

INVx1_ASAP7_75t_L g19791 ( 
.A(n_19583),
.Y(n_19791)
);

OAI22xp33_ASAP7_75t_L g19792 ( 
.A1(n_19349),
.A2(n_12471),
.B1(n_12496),
.B2(n_12451),
.Y(n_19792)
);

NAND3x2_ASAP7_75t_L g19793 ( 
.A(n_19647),
.B(n_9075),
.C(n_9013),
.Y(n_19793)
);

AOI32xp33_ASAP7_75t_L g19794 ( 
.A1(n_19430),
.A2(n_9013),
.A3(n_9093),
.B1(n_9091),
.B2(n_9078),
.Y(n_19794)
);

CKINVDCx14_ASAP7_75t_R g19795 ( 
.A(n_19513),
.Y(n_19795)
);

OAI21xp5_ASAP7_75t_L g19796 ( 
.A1(n_19584),
.A2(n_11595),
.B(n_11583),
.Y(n_19796)
);

HB1xp67_ASAP7_75t_L g19797 ( 
.A(n_19535),
.Y(n_19797)
);

INVx2_ASAP7_75t_SL g19798 ( 
.A(n_19535),
.Y(n_19798)
);

INVx2_ASAP7_75t_SL g19799 ( 
.A(n_19422),
.Y(n_19799)
);

INVx1_ASAP7_75t_L g19800 ( 
.A(n_19589),
.Y(n_19800)
);

OR2x2_ASAP7_75t_L g19801 ( 
.A(n_19414),
.B(n_12343),
.Y(n_19801)
);

AND2x2_ASAP7_75t_L g19802 ( 
.A(n_19488),
.B(n_9345),
.Y(n_19802)
);

AND2x2_ASAP7_75t_L g19803 ( 
.A(n_19498),
.B(n_9345),
.Y(n_19803)
);

INVx1_ASAP7_75t_L g19804 ( 
.A(n_19463),
.Y(n_19804)
);

NOR2x1_ASAP7_75t_L g19805 ( 
.A(n_19565),
.B(n_10180),
.Y(n_19805)
);

INVx1_ASAP7_75t_L g19806 ( 
.A(n_19495),
.Y(n_19806)
);

INVx1_ASAP7_75t_L g19807 ( 
.A(n_19507),
.Y(n_19807)
);

INVx1_ASAP7_75t_L g19808 ( 
.A(n_19510),
.Y(n_19808)
);

OAI22xp5_ASAP7_75t_L g19809 ( 
.A1(n_19383),
.A2(n_9091),
.B1(n_9093),
.B2(n_9078),
.Y(n_19809)
);

OAI221xp5_ASAP7_75t_L g19810 ( 
.A1(n_19346),
.A2(n_10131),
.B1(n_10104),
.B2(n_9156),
.C(n_9266),
.Y(n_19810)
);

AO22x1_ASAP7_75t_L g19811 ( 
.A1(n_19680),
.A2(n_9078),
.B1(n_9189),
.B2(n_9093),
.Y(n_19811)
);

INVx1_ASAP7_75t_L g19812 ( 
.A(n_19549),
.Y(n_19812)
);

OAI21xp33_ASAP7_75t_L g19813 ( 
.A1(n_19382),
.A2(n_9562),
.B(n_9559),
.Y(n_19813)
);

NOR2xp33_ASAP7_75t_L g19814 ( 
.A(n_19487),
.B(n_8449),
.Y(n_19814)
);

AOI22xp5_ASAP7_75t_L g19815 ( 
.A1(n_19395),
.A2(n_9455),
.B1(n_9456),
.B2(n_9391),
.Y(n_19815)
);

OAI22xp5_ASAP7_75t_L g19816 ( 
.A1(n_19505),
.A2(n_9295),
.B1(n_9189),
.B2(n_8981),
.Y(n_19816)
);

OAI22xp5_ASAP7_75t_L g19817 ( 
.A1(n_19473),
.A2(n_19399),
.B1(n_19480),
.B2(n_19432),
.Y(n_19817)
);

INVxp33_ASAP7_75t_L g19818 ( 
.A(n_19475),
.Y(n_19818)
);

INVx2_ASAP7_75t_L g19819 ( 
.A(n_19343),
.Y(n_19819)
);

INVx2_ASAP7_75t_L g19820 ( 
.A(n_19351),
.Y(n_19820)
);

AOI22xp5_ASAP7_75t_L g19821 ( 
.A1(n_19431),
.A2(n_9455),
.B1(n_9456),
.B2(n_9391),
.Y(n_19821)
);

INVx1_ASAP7_75t_L g19822 ( 
.A(n_19550),
.Y(n_19822)
);

INVx1_ASAP7_75t_L g19823 ( 
.A(n_19592),
.Y(n_19823)
);

INVx1_ASAP7_75t_L g19824 ( 
.A(n_19593),
.Y(n_19824)
);

INVx1_ASAP7_75t_L g19825 ( 
.A(n_19602),
.Y(n_19825)
);

NAND2xp5_ASAP7_75t_L g19826 ( 
.A(n_19508),
.B(n_10039),
.Y(n_19826)
);

INVx1_ASAP7_75t_L g19827 ( 
.A(n_19530),
.Y(n_19827)
);

OR2x2_ASAP7_75t_L g19828 ( 
.A(n_19355),
.B(n_12421),
.Y(n_19828)
);

AOI32xp33_ASAP7_75t_L g19829 ( 
.A1(n_19423),
.A2(n_9189),
.A3(n_9295),
.B1(n_10350),
.B2(n_10347),
.Y(n_19829)
);

AND2x2_ASAP7_75t_L g19830 ( 
.A(n_19511),
.B(n_9345),
.Y(n_19830)
);

O2A1O1Ixp33_ASAP7_75t_L g19831 ( 
.A1(n_19685),
.A2(n_10359),
.B(n_10372),
.C(n_10353),
.Y(n_19831)
);

OAI21xp33_ASAP7_75t_SL g19832 ( 
.A1(n_19381),
.A2(n_10924),
.B(n_10672),
.Y(n_19832)
);

INVx1_ASAP7_75t_L g19833 ( 
.A(n_19607),
.Y(n_19833)
);

NOR2xp33_ASAP7_75t_L g19834 ( 
.A(n_19700),
.B(n_8449),
.Y(n_19834)
);

INVx1_ASAP7_75t_L g19835 ( 
.A(n_19608),
.Y(n_19835)
);

INVxp67_ASAP7_75t_SL g19836 ( 
.A(n_19678),
.Y(n_19836)
);

NAND2xp5_ASAP7_75t_L g19837 ( 
.A(n_19385),
.B(n_10039),
.Y(n_19837)
);

INVx1_ASAP7_75t_L g19838 ( 
.A(n_19611),
.Y(n_19838)
);

NAND2xp5_ASAP7_75t_L g19839 ( 
.A(n_19523),
.B(n_10055),
.Y(n_19839)
);

A2O1A1Ixp33_ASAP7_75t_L g19840 ( 
.A1(n_19588),
.A2(n_11379),
.B(n_11368),
.C(n_11251),
.Y(n_19840)
);

INVx1_ASAP7_75t_L g19841 ( 
.A(n_19407),
.Y(n_19841)
);

NAND2xp5_ASAP7_75t_L g19842 ( 
.A(n_19526),
.B(n_10055),
.Y(n_19842)
);

NAND2xp5_ASAP7_75t_L g19843 ( 
.A(n_19401),
.B(n_19412),
.Y(n_19843)
);

OAI22xp5_ASAP7_75t_L g19844 ( 
.A1(n_19477),
.A2(n_9295),
.B1(n_8981),
.B2(n_9084),
.Y(n_19844)
);

NOR2x1_ASAP7_75t_L g19845 ( 
.A(n_19629),
.B(n_10180),
.Y(n_19845)
);

OAI21xp33_ASAP7_75t_L g19846 ( 
.A1(n_19444),
.A2(n_9562),
.B(n_9559),
.Y(n_19846)
);

NAND2xp5_ASAP7_75t_L g19847 ( 
.A(n_19528),
.B(n_10055),
.Y(n_19847)
);

AOI22xp33_ASAP7_75t_SL g19848 ( 
.A1(n_19396),
.A2(n_9455),
.B1(n_9456),
.B2(n_9391),
.Y(n_19848)
);

INVx1_ASAP7_75t_L g19849 ( 
.A(n_19409),
.Y(n_19849)
);

INVx1_ASAP7_75t_L g19850 ( 
.A(n_19552),
.Y(n_19850)
);

INVx1_ASAP7_75t_L g19851 ( 
.A(n_19532),
.Y(n_19851)
);

OAI22xp33_ASAP7_75t_L g19852 ( 
.A1(n_19484),
.A2(n_12471),
.B1(n_12496),
.B2(n_12451),
.Y(n_19852)
);

AOI22xp5_ASAP7_75t_L g19853 ( 
.A1(n_19506),
.A2(n_9391),
.B1(n_9456),
.B2(n_9455),
.Y(n_19853)
);

AOI22xp33_ASAP7_75t_L g19854 ( 
.A1(n_19474),
.A2(n_10078),
.B1(n_10094),
.B2(n_10055),
.Y(n_19854)
);

INVx1_ASAP7_75t_L g19855 ( 
.A(n_19533),
.Y(n_19855)
);

AOI21xp5_ASAP7_75t_L g19856 ( 
.A1(n_19667),
.A2(n_12556),
.B(n_12496),
.Y(n_19856)
);

INVx2_ASAP7_75t_SL g19857 ( 
.A(n_19511),
.Y(n_19857)
);

AOI21x1_ASAP7_75t_L g19858 ( 
.A1(n_19442),
.A2(n_10931),
.B(n_10876),
.Y(n_19858)
);

NAND2xp5_ASAP7_75t_L g19859 ( 
.A(n_19537),
.B(n_10055),
.Y(n_19859)
);

INVxp67_ASAP7_75t_L g19860 ( 
.A(n_19538),
.Y(n_19860)
);

AOI32xp33_ASAP7_75t_L g19861 ( 
.A1(n_19410),
.A2(n_19542),
.A3(n_19545),
.B1(n_19544),
.B2(n_19543),
.Y(n_19861)
);

AOI22xp5_ASAP7_75t_SL g19862 ( 
.A1(n_19560),
.A2(n_9763),
.B1(n_10006),
.B2(n_9828),
.Y(n_19862)
);

INVx1_ASAP7_75t_L g19863 ( 
.A(n_19561),
.Y(n_19863)
);

NAND2x1p5_ASAP7_75t_L g19864 ( 
.A(n_19562),
.B(n_9636),
.Y(n_19864)
);

NAND2xp5_ASAP7_75t_L g19865 ( 
.A(n_19568),
.B(n_19572),
.Y(n_19865)
);

INVx1_ASAP7_75t_L g19866 ( 
.A(n_19573),
.Y(n_19866)
);

AOI21xp5_ASAP7_75t_L g19867 ( 
.A1(n_19668),
.A2(n_12585),
.B(n_12556),
.Y(n_19867)
);

OAI21xp5_ASAP7_75t_L g19868 ( 
.A1(n_19605),
.A2(n_19591),
.B(n_19586),
.Y(n_19868)
);

OAI22xp33_ASAP7_75t_L g19869 ( 
.A1(n_19427),
.A2(n_12585),
.B1(n_12556),
.B2(n_10353),
.Y(n_19869)
);

NAND2xp5_ASAP7_75t_L g19870 ( 
.A(n_19623),
.B(n_10055),
.Y(n_19870)
);

OAI22xp5_ASAP7_75t_L g19871 ( 
.A1(n_19428),
.A2(n_9295),
.B1(n_8981),
.B2(n_9084),
.Y(n_19871)
);

INVx1_ASAP7_75t_L g19872 ( 
.A(n_19479),
.Y(n_19872)
);

NAND2x1_ASAP7_75t_L g19873 ( 
.A(n_19458),
.B(n_9662),
.Y(n_19873)
);

INVxp33_ASAP7_75t_L g19874 ( 
.A(n_19622),
.Y(n_19874)
);

OAI21xp5_ASAP7_75t_L g19875 ( 
.A1(n_19599),
.A2(n_11604),
.B(n_11596),
.Y(n_19875)
);

AOI22xp5_ASAP7_75t_L g19876 ( 
.A1(n_19566),
.A2(n_9455),
.B1(n_9456),
.B2(n_9391),
.Y(n_19876)
);

OR2x2_ASAP7_75t_L g19877 ( 
.A(n_19352),
.B(n_12421),
.Y(n_19877)
);

OAI21xp5_ASAP7_75t_L g19878 ( 
.A1(n_19451),
.A2(n_11604),
.B(n_11596),
.Y(n_19878)
);

INVxp67_ASAP7_75t_L g19879 ( 
.A(n_19626),
.Y(n_19879)
);

INVx1_ASAP7_75t_L g19880 ( 
.A(n_19493),
.Y(n_19880)
);

NAND2xp5_ASAP7_75t_L g19881 ( 
.A(n_19594),
.B(n_10055),
.Y(n_19881)
);

NOR2xp33_ASAP7_75t_L g19882 ( 
.A(n_19693),
.B(n_8449),
.Y(n_19882)
);

OAI22xp33_ASAP7_75t_L g19883 ( 
.A1(n_19429),
.A2(n_12585),
.B1(n_10372),
.B2(n_10389),
.Y(n_19883)
);

BUFx2_ASAP7_75t_L g19884 ( 
.A(n_19348),
.Y(n_19884)
);

OR2x2_ASAP7_75t_L g19885 ( 
.A(n_19420),
.B(n_12421),
.Y(n_19885)
);

NAND2xp5_ASAP7_75t_L g19886 ( 
.A(n_19653),
.B(n_10055),
.Y(n_19886)
);

OAI32xp33_ASAP7_75t_L g19887 ( 
.A1(n_19478),
.A2(n_19699),
.A3(n_19437),
.B1(n_19452),
.B2(n_19445),
.Y(n_19887)
);

INVxp33_ASAP7_75t_L g19888 ( 
.A(n_19404),
.Y(n_19888)
);

OR2x2_ASAP7_75t_L g19889 ( 
.A(n_19440),
.B(n_12093),
.Y(n_19889)
);

NAND3xp33_ASAP7_75t_SL g19890 ( 
.A(n_19666),
.B(n_10131),
.C(n_10104),
.Y(n_19890)
);

NAND2xp5_ASAP7_75t_L g19891 ( 
.A(n_19628),
.B(n_10078),
.Y(n_19891)
);

AND2x2_ASAP7_75t_L g19892 ( 
.A(n_19603),
.B(n_9345),
.Y(n_19892)
);

INVx2_ASAP7_75t_L g19893 ( 
.A(n_19689),
.Y(n_19893)
);

AND2x2_ASAP7_75t_L g19894 ( 
.A(n_19609),
.B(n_9345),
.Y(n_19894)
);

NAND2xp5_ASAP7_75t_L g19895 ( 
.A(n_19631),
.B(n_10078),
.Y(n_19895)
);

INVx2_ASAP7_75t_SL g19896 ( 
.A(n_19630),
.Y(n_19896)
);

INVxp67_ASAP7_75t_SL g19897 ( 
.A(n_19577),
.Y(n_19897)
);

AOI221xp5_ASAP7_75t_L g19898 ( 
.A1(n_19524),
.A2(n_10389),
.B1(n_10486),
.B2(n_10372),
.C(n_10359),
.Y(n_19898)
);

NAND2xp5_ASAP7_75t_L g19899 ( 
.A(n_19634),
.B(n_10078),
.Y(n_19899)
);

HB1xp67_ASAP7_75t_L g19900 ( 
.A(n_19659),
.Y(n_19900)
);

AND2x2_ASAP7_75t_L g19901 ( 
.A(n_19625),
.B(n_9345),
.Y(n_19901)
);

OAI22xp5_ASAP7_75t_L g19902 ( 
.A1(n_19496),
.A2(n_9084),
.B1(n_9744),
.B2(n_9636),
.Y(n_19902)
);

INVx2_ASAP7_75t_L g19903 ( 
.A(n_19657),
.Y(n_19903)
);

INVx1_ASAP7_75t_L g19904 ( 
.A(n_19379),
.Y(n_19904)
);

BUFx2_ASAP7_75t_SL g19905 ( 
.A(n_19703),
.Y(n_19905)
);

AND2x2_ASAP7_75t_L g19906 ( 
.A(n_19516),
.B(n_9445),
.Y(n_19906)
);

INVx1_ASAP7_75t_L g19907 ( 
.A(n_19384),
.Y(n_19907)
);

INVx1_ASAP7_75t_L g19908 ( 
.A(n_19546),
.Y(n_19908)
);

OAI211xp5_ASAP7_75t_SL g19909 ( 
.A1(n_19632),
.A2(n_9766),
.B(n_9717),
.C(n_9659),
.Y(n_19909)
);

INVx2_ASAP7_75t_SL g19910 ( 
.A(n_19468),
.Y(n_19910)
);

NAND2xp5_ASAP7_75t_L g19911 ( 
.A(n_19635),
.B(n_10078),
.Y(n_19911)
);

OAI22xp33_ASAP7_75t_SL g19912 ( 
.A1(n_19615),
.A2(n_10131),
.B1(n_10486),
.B2(n_10389),
.Y(n_19912)
);

OR2x2_ASAP7_75t_L g19913 ( 
.A(n_19469),
.B(n_19425),
.Y(n_19913)
);

OAI21xp33_ASAP7_75t_L g19914 ( 
.A1(n_19519),
.A2(n_9562),
.B(n_9559),
.Y(n_19914)
);

NAND2xp5_ASAP7_75t_SL g19915 ( 
.A(n_19529),
.B(n_9391),
.Y(n_19915)
);

INVx1_ASAP7_75t_L g19916 ( 
.A(n_19472),
.Y(n_19916)
);

NOR2xp33_ASAP7_75t_L g19917 ( 
.A(n_19654),
.B(n_8449),
.Y(n_19917)
);

INVx1_ASAP7_75t_L g19918 ( 
.A(n_19501),
.Y(n_19918)
);

INVx1_ASAP7_75t_L g19919 ( 
.A(n_19514),
.Y(n_19919)
);

INVxp67_ASAP7_75t_L g19920 ( 
.A(n_19664),
.Y(n_19920)
);

INVxp67_ASAP7_75t_L g19921 ( 
.A(n_19672),
.Y(n_19921)
);

INVx1_ASAP7_75t_L g19922 ( 
.A(n_19555),
.Y(n_19922)
);

AND2x2_ASAP7_75t_L g19923 ( 
.A(n_19497),
.B(n_9445),
.Y(n_19923)
);

INVx1_ASAP7_75t_SL g19924 ( 
.A(n_19344),
.Y(n_19924)
);

INVx1_ASAP7_75t_SL g19925 ( 
.A(n_19686),
.Y(n_19925)
);

NAND2x1p5_ASAP7_75t_L g19926 ( 
.A(n_19690),
.B(n_9636),
.Y(n_19926)
);

INVxp67_ASAP7_75t_L g19927 ( 
.A(n_19636),
.Y(n_19927)
);

AND2x2_ASAP7_75t_L g19928 ( 
.A(n_19563),
.B(n_9445),
.Y(n_19928)
);

INVx1_ASAP7_75t_L g19929 ( 
.A(n_19559),
.Y(n_19929)
);

OAI221xp5_ASAP7_75t_SL g19930 ( 
.A1(n_19551),
.A2(n_9377),
.B1(n_9333),
.B2(n_9725),
.C(n_9704),
.Y(n_19930)
);

INVx1_ASAP7_75t_L g19931 ( 
.A(n_19569),
.Y(n_19931)
);

AOI21xp5_ASAP7_75t_L g19932 ( 
.A1(n_19372),
.A2(n_12683),
.B(n_12626),
.Y(n_19932)
);

INVx1_ASAP7_75t_L g19933 ( 
.A(n_19406),
.Y(n_19933)
);

INVx1_ASAP7_75t_L g19934 ( 
.A(n_19641),
.Y(n_19934)
);

NOR3xp33_ASAP7_75t_L g19935 ( 
.A(n_19679),
.B(n_8088),
.C(n_8020),
.Y(n_19935)
);

INVx1_ASAP7_75t_L g19936 ( 
.A(n_19642),
.Y(n_19936)
);

AND2x2_ASAP7_75t_L g19937 ( 
.A(n_19687),
.B(n_9445),
.Y(n_19937)
);

NOR2x1_ASAP7_75t_L g19938 ( 
.A(n_19643),
.B(n_10180),
.Y(n_19938)
);

NAND2xp5_ASAP7_75t_L g19939 ( 
.A(n_19645),
.B(n_10078),
.Y(n_19939)
);

AOI21xp5_ASAP7_75t_L g19940 ( 
.A1(n_19606),
.A2(n_12683),
.B(n_12626),
.Y(n_19940)
);

INVx1_ASAP7_75t_L g19941 ( 
.A(n_19649),
.Y(n_19941)
);

INVx1_ASAP7_75t_L g19942 ( 
.A(n_19658),
.Y(n_19942)
);

INVx1_ASAP7_75t_L g19943 ( 
.A(n_19660),
.Y(n_19943)
);

AOI22xp33_ASAP7_75t_SL g19944 ( 
.A1(n_19587),
.A2(n_9391),
.B1(n_9456),
.B2(n_9455),
.Y(n_19944)
);

AND2x4_ASAP7_75t_L g19945 ( 
.A(n_19661),
.B(n_10931),
.Y(n_19945)
);

INVx1_ASAP7_75t_L g19946 ( 
.A(n_19665),
.Y(n_19946)
);

OR2x2_ASAP7_75t_L g19947 ( 
.A(n_19476),
.B(n_12110),
.Y(n_19947)
);

INVx1_ASAP7_75t_L g19948 ( 
.A(n_19669),
.Y(n_19948)
);

NOR2xp33_ASAP7_75t_L g19949 ( 
.A(n_19674),
.B(n_8449),
.Y(n_19949)
);

OAI22xp33_ASAP7_75t_L g19950 ( 
.A1(n_19390),
.A2(n_10506),
.B1(n_10511),
.B2(n_10486),
.Y(n_19950)
);

AND2x2_ASAP7_75t_L g19951 ( 
.A(n_19676),
.B(n_9445),
.Y(n_19951)
);

INVx3_ASAP7_75t_L g19952 ( 
.A(n_19646),
.Y(n_19952)
);

INVx1_ASAP7_75t_L g19953 ( 
.A(n_19682),
.Y(n_19953)
);

NAND2xp5_ASAP7_75t_L g19954 ( 
.A(n_19694),
.B(n_19701),
.Y(n_19954)
);

NOR2xp67_ASAP7_75t_SL g19955 ( 
.A(n_19618),
.B(n_19610),
.Y(n_19955)
);

INVxp67_ASAP7_75t_L g19956 ( 
.A(n_19614),
.Y(n_19956)
);

INVx1_ASAP7_75t_L g19957 ( 
.A(n_19617),
.Y(n_19957)
);

BUFx4f_ASAP7_75t_SL g19958 ( 
.A(n_19578),
.Y(n_19958)
);

INVx1_ASAP7_75t_L g19959 ( 
.A(n_19570),
.Y(n_19959)
);

NAND4xp25_ASAP7_75t_SL g19960 ( 
.A(n_19503),
.B(n_19579),
.C(n_19601),
.D(n_19598),
.Y(n_19960)
);

OAI21xp5_ASAP7_75t_L g19961 ( 
.A1(n_19581),
.A2(n_11604),
.B(n_11596),
.Y(n_19961)
);

NAND2xp5_ASAP7_75t_L g19962 ( 
.A(n_19655),
.B(n_10078),
.Y(n_19962)
);

INVxp67_ASAP7_75t_SL g19963 ( 
.A(n_19604),
.Y(n_19963)
);

OR2x2_ASAP7_75t_L g19964 ( 
.A(n_19576),
.B(n_12176),
.Y(n_19964)
);

OAI21xp33_ASAP7_75t_SL g19965 ( 
.A1(n_19350),
.A2(n_10924),
.B(n_10672),
.Y(n_19965)
);

INVx1_ASAP7_75t_L g19966 ( 
.A(n_19595),
.Y(n_19966)
);

INVx1_ASAP7_75t_L g19967 ( 
.A(n_19627),
.Y(n_19967)
);

OR2x2_ASAP7_75t_L g19968 ( 
.A(n_19575),
.B(n_12176),
.Y(n_19968)
);

INVx2_ASAP7_75t_L g19969 ( 
.A(n_19662),
.Y(n_19969)
);

INVx1_ASAP7_75t_L g19970 ( 
.A(n_19637),
.Y(n_19970)
);

AOI22xp5_ASAP7_75t_L g19971 ( 
.A1(n_19597),
.A2(n_19652),
.B1(n_19522),
.B2(n_19684),
.Y(n_19971)
);

AND2x2_ASAP7_75t_L g19972 ( 
.A(n_19464),
.B(n_9445),
.Y(n_19972)
);

AOI21xp33_ASAP7_75t_SL g19973 ( 
.A1(n_19457),
.A2(n_10131),
.B(n_9156),
.Y(n_19973)
);

OA21x2_ASAP7_75t_L g19974 ( 
.A1(n_19373),
.A2(n_11252),
.B(n_11251),
.Y(n_19974)
);

OAI21xp33_ASAP7_75t_L g19975 ( 
.A1(n_19438),
.A2(n_9586),
.B(n_9576),
.Y(n_19975)
);

NOR2x1_ASAP7_75t_L g19976 ( 
.A(n_19696),
.B(n_10180),
.Y(n_19976)
);

OR2x2_ASAP7_75t_L g19977 ( 
.A(n_19621),
.B(n_12176),
.Y(n_19977)
);

NAND2xp5_ASAP7_75t_L g19978 ( 
.A(n_19557),
.B(n_10078),
.Y(n_19978)
);

A2O1A1Ixp33_ASAP7_75t_L g19979 ( 
.A1(n_19462),
.A2(n_11379),
.B(n_11251),
.C(n_11252),
.Y(n_19979)
);

OAI21xp5_ASAP7_75t_SL g19980 ( 
.A1(n_19435),
.A2(n_10131),
.B(n_9156),
.Y(n_19980)
);

AOI222xp33_ASAP7_75t_L g19981 ( 
.A1(n_19518),
.A2(n_10486),
.B1(n_10511),
.B2(n_10542),
.C1(n_10522),
.C2(n_10506),
.Y(n_19981)
);

AOI21xp33_ASAP7_75t_L g19982 ( 
.A1(n_19670),
.A2(n_19673),
.B(n_19640),
.Y(n_19982)
);

OAI21xp5_ASAP7_75t_L g19983 ( 
.A1(n_19443),
.A2(n_10802),
.B(n_10205),
.Y(n_19983)
);

AOI21xp33_ASAP7_75t_SL g19984 ( 
.A1(n_19456),
.A2(n_9156),
.B(n_9065),
.Y(n_19984)
);

OR2x2_ASAP7_75t_L g19985 ( 
.A(n_19695),
.B(n_12248),
.Y(n_19985)
);

NAND2xp5_ASAP7_75t_L g19986 ( 
.A(n_19369),
.B(n_10078),
.Y(n_19986)
);

AND2x2_ASAP7_75t_L g19987 ( 
.A(n_19389),
.B(n_9445),
.Y(n_19987)
);

OAI211xp5_ASAP7_75t_L g19988 ( 
.A1(n_19644),
.A2(n_8992),
.B(n_9199),
.C(n_9145),
.Y(n_19988)
);

AND2x2_ASAP7_75t_L g19989 ( 
.A(n_19616),
.B(n_9445),
.Y(n_19989)
);

OAI322xp33_ASAP7_75t_L g19990 ( 
.A1(n_19590),
.A2(n_10542),
.A3(n_10511),
.B1(n_10549),
.B2(n_10563),
.C1(n_10522),
.C2(n_10506),
.Y(n_19990)
);

AOI22xp5_ASAP7_75t_L g19991 ( 
.A1(n_19585),
.A2(n_9391),
.B1(n_9456),
.B2(n_9455),
.Y(n_19991)
);

INVx1_ASAP7_75t_L g19992 ( 
.A(n_19394),
.Y(n_19992)
);

INVx1_ASAP7_75t_L g19993 ( 
.A(n_19394),
.Y(n_19993)
);

INVx2_ASAP7_75t_L g19994 ( 
.A(n_19692),
.Y(n_19994)
);

OAI21xp5_ASAP7_75t_L g19995 ( 
.A1(n_19663),
.A2(n_10802),
.B(n_10205),
.Y(n_19995)
);

NAND2xp5_ASAP7_75t_L g19996 ( 
.A(n_19567),
.B(n_10094),
.Y(n_19996)
);

AOI22xp33_ASAP7_75t_SL g19997 ( 
.A1(n_19466),
.A2(n_9455),
.B1(n_9468),
.B2(n_9456),
.Y(n_19997)
);

AOI21xp33_ASAP7_75t_SL g19998 ( 
.A1(n_19677),
.A2(n_9156),
.B(n_9065),
.Y(n_19998)
);

OAI32xp33_ASAP7_75t_L g19999 ( 
.A1(n_19675),
.A2(n_10522),
.A3(n_10542),
.B1(n_10511),
.B2(n_10506),
.Y(n_19999)
);

OAI22x1_ASAP7_75t_L g20000 ( 
.A1(n_19392),
.A2(n_9199),
.B1(n_8992),
.B2(n_9145),
.Y(n_20000)
);

INVx2_ASAP7_75t_L g20001 ( 
.A(n_19366),
.Y(n_20001)
);

NAND2xp5_ASAP7_75t_SL g20002 ( 
.A(n_19424),
.B(n_9455),
.Y(n_20002)
);

NAND2xp5_ASAP7_75t_L g20003 ( 
.A(n_19483),
.B(n_10094),
.Y(n_20003)
);

INVx2_ASAP7_75t_L g20004 ( 
.A(n_19454),
.Y(n_20004)
);

INVx1_ASAP7_75t_L g20005 ( 
.A(n_19481),
.Y(n_20005)
);

AOI22xp33_ASAP7_75t_L g20006 ( 
.A1(n_19547),
.A2(n_10118),
.B1(n_10139),
.B2(n_10094),
.Y(n_20006)
);

AOI21xp33_ASAP7_75t_L g20007 ( 
.A1(n_19450),
.A2(n_12257),
.B(n_12248),
.Y(n_20007)
);

AOI221xp5_ASAP7_75t_L g20008 ( 
.A1(n_19683),
.A2(n_10549),
.B1(n_10563),
.B2(n_10542),
.C(n_10522),
.Y(n_20008)
);

NAND2xp5_ASAP7_75t_L g20009 ( 
.A(n_19465),
.B(n_10094),
.Y(n_20009)
);

INVx1_ASAP7_75t_L g20010 ( 
.A(n_19600),
.Y(n_20010)
);

INVx2_ASAP7_75t_SL g20011 ( 
.A(n_19486),
.Y(n_20011)
);

INVx1_ASAP7_75t_L g20012 ( 
.A(n_19398),
.Y(n_20012)
);

OAI21xp33_ASAP7_75t_L g20013 ( 
.A1(n_19446),
.A2(n_9586),
.B(n_9576),
.Y(n_20013)
);

INVx1_ASAP7_75t_L g20014 ( 
.A(n_19688),
.Y(n_20014)
);

INVx1_ASAP7_75t_L g20015 ( 
.A(n_19783),
.Y(n_20015)
);

AND2x2_ASAP7_75t_L g20016 ( 
.A(n_19704),
.B(n_19490),
.Y(n_20016)
);

NAND2xp5_ASAP7_75t_L g20017 ( 
.A(n_19705),
.B(n_19371),
.Y(n_20017)
);

AO21x1_ASAP7_75t_L g20018 ( 
.A1(n_19992),
.A2(n_19359),
.B(n_19377),
.Y(n_20018)
);

NAND2xp5_ASAP7_75t_L g20019 ( 
.A(n_19713),
.B(n_19633),
.Y(n_20019)
);

OAI32xp33_ASAP7_75t_L g20020 ( 
.A1(n_20010),
.A2(n_19620),
.A3(n_19357),
.B1(n_19556),
.B2(n_19421),
.Y(n_20020)
);

NAND2xp5_ASAP7_75t_L g20021 ( 
.A(n_19762),
.B(n_19467),
.Y(n_20021)
);

INVx1_ASAP7_75t_L g20022 ( 
.A(n_19783),
.Y(n_20022)
);

AOI322xp5_ASAP7_75t_L g20023 ( 
.A1(n_19836),
.A2(n_19761),
.A3(n_19765),
.B1(n_19773),
.B2(n_19775),
.C1(n_19771),
.C2(n_19707),
.Y(n_20023)
);

XNOR2x1_ASAP7_75t_L g20024 ( 
.A(n_19704),
.B(n_19361),
.Y(n_20024)
);

AOI21xp5_ASAP7_75t_L g20025 ( 
.A1(n_19756),
.A2(n_19723),
.B(n_19896),
.Y(n_20025)
);

NAND2xp5_ASAP7_75t_L g20026 ( 
.A(n_19706),
.B(n_19691),
.Y(n_20026)
);

AND2x2_ASAP7_75t_L g20027 ( 
.A(n_19827),
.B(n_19624),
.Y(n_20027)
);

INVx1_ASAP7_75t_L g20028 ( 
.A(n_19772),
.Y(n_20028)
);

INVx1_ASAP7_75t_L g20029 ( 
.A(n_19993),
.Y(n_20029)
);

INVx2_ASAP7_75t_SL g20030 ( 
.A(n_19714),
.Y(n_20030)
);

AOI22xp33_ASAP7_75t_SL g20031 ( 
.A1(n_19795),
.A2(n_19534),
.B1(n_19638),
.B2(n_19499),
.Y(n_20031)
);

INVx1_ASAP7_75t_L g20032 ( 
.A(n_19758),
.Y(n_20032)
);

OAI222xp33_ASAP7_75t_L g20033 ( 
.A1(n_19734),
.A2(n_19504),
.B1(n_19509),
.B2(n_19417),
.C1(n_19681),
.C2(n_19582),
.Y(n_20033)
);

AOI222xp33_ASAP7_75t_L g20034 ( 
.A1(n_19958),
.A2(n_19702),
.B1(n_19613),
.B2(n_19515),
.C1(n_10549),
.C2(n_10575),
.Y(n_20034)
);

OAI21xp5_ASAP7_75t_L g20035 ( 
.A1(n_19860),
.A2(n_10802),
.B(n_10205),
.Y(n_20035)
);

AND2x2_ASAP7_75t_L g20036 ( 
.A(n_19807),
.B(n_9452),
.Y(n_20036)
);

OR2x2_ASAP7_75t_L g20037 ( 
.A(n_19715),
.B(n_12248),
.Y(n_20037)
);

AOI21xp33_ASAP7_75t_L g20038 ( 
.A1(n_19735),
.A2(n_12257),
.B(n_12626),
.Y(n_20038)
);

NOR2xp33_ASAP7_75t_SL g20039 ( 
.A(n_19739),
.B(n_9411),
.Y(n_20039)
);

NAND2xp5_ASAP7_75t_L g20040 ( 
.A(n_19716),
.B(n_10094),
.Y(n_20040)
);

NAND3xp33_ASAP7_75t_L g20041 ( 
.A(n_19861),
.B(n_9468),
.C(n_9456),
.Y(n_20041)
);

AOI221xp5_ASAP7_75t_L g20042 ( 
.A1(n_19720),
.A2(n_10575),
.B1(n_10578),
.B2(n_10563),
.C(n_10549),
.Y(n_20042)
);

NAND2xp5_ASAP7_75t_SL g20043 ( 
.A(n_19731),
.B(n_9456),
.Y(n_20043)
);

INVx1_ASAP7_75t_L g20044 ( 
.A(n_19730),
.Y(n_20044)
);

OAI31xp33_ASAP7_75t_L g20045 ( 
.A1(n_19719),
.A2(n_9578),
.A3(n_9595),
.B(n_9493),
.Y(n_20045)
);

OAI22xp5_ASAP7_75t_L g20046 ( 
.A1(n_19742),
.A2(n_9744),
.B1(n_9636),
.B2(n_9586),
.Y(n_20046)
);

AOI22xp5_ASAP7_75t_L g20047 ( 
.A1(n_19808),
.A2(n_9476),
.B1(n_9566),
.B2(n_9468),
.Y(n_20047)
);

INVx1_ASAP7_75t_L g20048 ( 
.A(n_19884),
.Y(n_20048)
);

INVx1_ASAP7_75t_L g20049 ( 
.A(n_19727),
.Y(n_20049)
);

INVx1_ASAP7_75t_L g20050 ( 
.A(n_19744),
.Y(n_20050)
);

NAND2xp5_ASAP7_75t_L g20051 ( 
.A(n_19787),
.B(n_10094),
.Y(n_20051)
);

OAI21xp33_ASAP7_75t_L g20052 ( 
.A1(n_19814),
.A2(n_19834),
.B(n_19748),
.Y(n_20052)
);

INVx1_ASAP7_75t_L g20053 ( 
.A(n_19722),
.Y(n_20053)
);

NAND2xp5_ASAP7_75t_L g20054 ( 
.A(n_20011),
.B(n_10094),
.Y(n_20054)
);

INVxp67_ASAP7_75t_L g20055 ( 
.A(n_19905),
.Y(n_20055)
);

INVx1_ASAP7_75t_L g20056 ( 
.A(n_19797),
.Y(n_20056)
);

NAND2xp5_ASAP7_75t_SL g20057 ( 
.A(n_19789),
.B(n_9468),
.Y(n_20057)
);

NOR3xp33_ASAP7_75t_L g20058 ( 
.A(n_19868),
.B(n_8088),
.C(n_8020),
.Y(n_20058)
);

INVxp33_ASAP7_75t_L g20059 ( 
.A(n_19882),
.Y(n_20059)
);

NOR2xp33_ASAP7_75t_SL g20060 ( 
.A(n_19743),
.B(n_9411),
.Y(n_20060)
);

INVx1_ASAP7_75t_L g20061 ( 
.A(n_19721),
.Y(n_20061)
);

AOI32xp33_ASAP7_75t_L g20062 ( 
.A1(n_20012),
.A2(n_10578),
.A3(n_10589),
.B1(n_10575),
.B2(n_10563),
.Y(n_20062)
);

NAND3x2_ASAP7_75t_L g20063 ( 
.A(n_19740),
.B(n_9066),
.C(n_9576),
.Y(n_20063)
);

OR2x2_ASAP7_75t_L g20064 ( 
.A(n_19709),
.B(n_12257),
.Y(n_20064)
);

OR2x2_ASAP7_75t_L g20065 ( 
.A(n_19754),
.B(n_12683),
.Y(n_20065)
);

AND2x2_ASAP7_75t_L g20066 ( 
.A(n_19774),
.B(n_9452),
.Y(n_20066)
);

OAI22xp33_ASAP7_75t_SL g20067 ( 
.A1(n_19915),
.A2(n_10578),
.B1(n_10589),
.B2(n_10575),
.Y(n_20067)
);

INVx1_ASAP7_75t_L g20068 ( 
.A(n_19718),
.Y(n_20068)
);

INVx3_ASAP7_75t_L g20069 ( 
.A(n_19778),
.Y(n_20069)
);

AO22x1_ASAP7_75t_L g20070 ( 
.A1(n_19897),
.A2(n_10589),
.B1(n_10590),
.B2(n_10578),
.Y(n_20070)
);

INVx1_ASAP7_75t_L g20071 ( 
.A(n_19725),
.Y(n_20071)
);

NAND3xp33_ASAP7_75t_L g20072 ( 
.A(n_19711),
.B(n_9476),
.C(n_9468),
.Y(n_20072)
);

NAND2xp5_ASAP7_75t_L g20073 ( 
.A(n_19712),
.B(n_10094),
.Y(n_20073)
);

INVx1_ASAP7_75t_L g20074 ( 
.A(n_19782),
.Y(n_20074)
);

AO22x1_ASAP7_75t_L g20075 ( 
.A1(n_19888),
.A2(n_10590),
.B1(n_10596),
.B2(n_10589),
.Y(n_20075)
);

INVx2_ASAP7_75t_L g20076 ( 
.A(n_19802),
.Y(n_20076)
);

OAI22xp33_ASAP7_75t_SL g20077 ( 
.A1(n_19970),
.A2(n_10596),
.B1(n_10599),
.B2(n_10590),
.Y(n_20077)
);

AOI22xp33_ASAP7_75t_L g20078 ( 
.A1(n_19806),
.A2(n_11265),
.B1(n_11264),
.B2(n_10139),
.Y(n_20078)
);

OAI22xp5_ASAP7_75t_L g20079 ( 
.A1(n_19710),
.A2(n_9744),
.B1(n_9636),
.B2(n_9586),
.Y(n_20079)
);

AOI21xp5_ASAP7_75t_L g20080 ( 
.A1(n_19724),
.A2(n_12725),
.B(n_12707),
.Y(n_20080)
);

NOR2xp33_ASAP7_75t_L g20081 ( 
.A(n_19788),
.B(n_8449),
.Y(n_20081)
);

OR2x2_ASAP7_75t_L g20082 ( 
.A(n_19791),
.B(n_12707),
.Y(n_20082)
);

AOI221x1_ASAP7_75t_SL g20083 ( 
.A1(n_19767),
.A2(n_9576),
.B1(n_9602),
.B2(n_9594),
.C(n_9588),
.Y(n_20083)
);

INVx2_ASAP7_75t_L g20084 ( 
.A(n_19803),
.Y(n_20084)
);

AOI222xp33_ASAP7_75t_L g20085 ( 
.A1(n_19726),
.A2(n_10590),
.B1(n_10599),
.B2(n_10675),
.C1(n_10606),
.C2(n_10596),
.Y(n_20085)
);

OAI21xp33_ASAP7_75t_SL g20086 ( 
.A1(n_19805),
.A2(n_10659),
.B(n_10639),
.Y(n_20086)
);

AOI21xp5_ASAP7_75t_L g20087 ( 
.A1(n_19865),
.A2(n_12725),
.B(n_12707),
.Y(n_20087)
);

AOI21xp5_ASAP7_75t_SL g20088 ( 
.A1(n_19857),
.A2(n_10180),
.B(n_9377),
.Y(n_20088)
);

AOI22xp5_ASAP7_75t_L g20089 ( 
.A1(n_19917),
.A2(n_9476),
.B1(n_9566),
.B2(n_9468),
.Y(n_20089)
);

NOR2xp67_ASAP7_75t_SL g20090 ( 
.A(n_19800),
.B(n_9005),
.Y(n_20090)
);

INVxp67_ASAP7_75t_L g20091 ( 
.A(n_19776),
.Y(n_20091)
);

INVx2_ASAP7_75t_L g20092 ( 
.A(n_19830),
.Y(n_20092)
);

AOI22xp5_ASAP7_75t_L g20093 ( 
.A1(n_19949),
.A2(n_9476),
.B1(n_9566),
.B2(n_9468),
.Y(n_20093)
);

OAI221xp5_ASAP7_75t_L g20094 ( 
.A1(n_19971),
.A2(n_9156),
.B1(n_9266),
.B2(n_9261),
.C(n_9065),
.Y(n_20094)
);

NAND2xp5_ASAP7_75t_L g20095 ( 
.A(n_20004),
.B(n_10118),
.Y(n_20095)
);

NAND2xp5_ASAP7_75t_L g20096 ( 
.A(n_19799),
.B(n_10118),
.Y(n_20096)
);

AOI22xp5_ASAP7_75t_L g20097 ( 
.A1(n_19760),
.A2(n_9476),
.B1(n_9566),
.B2(n_9468),
.Y(n_20097)
);

INVx2_ASAP7_75t_L g20098 ( 
.A(n_19937),
.Y(n_20098)
);

AOI22xp5_ASAP7_75t_L g20099 ( 
.A1(n_19925),
.A2(n_19790),
.B1(n_19824),
.B2(n_19823),
.Y(n_20099)
);

OAI31xp33_ASAP7_75t_L g20100 ( 
.A1(n_19708),
.A2(n_19728),
.A3(n_19817),
.B(n_19825),
.Y(n_20100)
);

AOI31xp33_ASAP7_75t_L g20101 ( 
.A1(n_19818),
.A2(n_9156),
.A3(n_9261),
.B(n_9065),
.Y(n_20101)
);

AOI221xp5_ASAP7_75t_L g20102 ( 
.A1(n_19982),
.A2(n_10606),
.B1(n_10675),
.B2(n_10599),
.C(n_10596),
.Y(n_20102)
);

AND2x4_ASAP7_75t_L g20103 ( 
.A(n_19820),
.B(n_19819),
.Y(n_20103)
);

INVx1_ASAP7_75t_L g20104 ( 
.A(n_19833),
.Y(n_20104)
);

INVx1_ASAP7_75t_L g20105 ( 
.A(n_19835),
.Y(n_20105)
);

OAI21xp33_ASAP7_75t_SL g20106 ( 
.A1(n_19763),
.A2(n_10659),
.B(n_10639),
.Y(n_20106)
);

INVx2_ASAP7_75t_SL g20107 ( 
.A(n_19951),
.Y(n_20107)
);

OAI32xp33_ASAP7_75t_L g20108 ( 
.A1(n_19838),
.A2(n_10675),
.A3(n_10743),
.B1(n_10606),
.B2(n_10599),
.Y(n_20108)
);

NOR2xp33_ASAP7_75t_L g20109 ( 
.A(n_19785),
.B(n_19893),
.Y(n_20109)
);

INVx1_ASAP7_75t_L g20110 ( 
.A(n_19952),
.Y(n_20110)
);

OAI21xp5_ASAP7_75t_L g20111 ( 
.A1(n_19879),
.A2(n_10210),
.B(n_10204),
.Y(n_20111)
);

AND2x2_ASAP7_75t_L g20112 ( 
.A(n_19903),
.B(n_9452),
.Y(n_20112)
);

AND2x2_ASAP7_75t_L g20113 ( 
.A(n_19994),
.B(n_9452),
.Y(n_20113)
);

INVx1_ASAP7_75t_L g20114 ( 
.A(n_19952),
.Y(n_20114)
);

INVx1_ASAP7_75t_L g20115 ( 
.A(n_19804),
.Y(n_20115)
);

NOR2xp33_ASAP7_75t_SL g20116 ( 
.A(n_19798),
.B(n_9411),
.Y(n_20116)
);

O2A1O1Ixp33_ASAP7_75t_L g20117 ( 
.A1(n_19900),
.A2(n_10675),
.B(n_10743),
.C(n_10606),
.Y(n_20117)
);

OR2x2_ASAP7_75t_L g20118 ( 
.A(n_19841),
.B(n_12725),
.Y(n_20118)
);

OR2x2_ASAP7_75t_L g20119 ( 
.A(n_19849),
.B(n_12730),
.Y(n_20119)
);

BUFx2_ASAP7_75t_SL g20120 ( 
.A(n_19755),
.Y(n_20120)
);

NAND2xp5_ASAP7_75t_L g20121 ( 
.A(n_20001),
.B(n_10118),
.Y(n_20121)
);

NAND2xp5_ASAP7_75t_L g20122 ( 
.A(n_19812),
.B(n_10118),
.Y(n_20122)
);

INVx1_ASAP7_75t_L g20123 ( 
.A(n_19822),
.Y(n_20123)
);

INVx2_ASAP7_75t_L g20124 ( 
.A(n_19892),
.Y(n_20124)
);

NAND2xp5_ASAP7_75t_L g20125 ( 
.A(n_19851),
.B(n_10118),
.Y(n_20125)
);

AND2x2_ASAP7_75t_L g20126 ( 
.A(n_19855),
.B(n_9452),
.Y(n_20126)
);

NAND2xp5_ASAP7_75t_L g20127 ( 
.A(n_19863),
.B(n_10118),
.Y(n_20127)
);

OAI22xp5_ASAP7_75t_L g20128 ( 
.A1(n_19793),
.A2(n_9744),
.B1(n_9636),
.B2(n_9594),
.Y(n_20128)
);

AOI22xp5_ASAP7_75t_L g20129 ( 
.A1(n_19935),
.A2(n_9468),
.B1(n_9566),
.B2(n_9476),
.Y(n_20129)
);

NAND4xp25_ASAP7_75t_SL g20130 ( 
.A(n_19732),
.B(n_8779),
.C(n_8783),
.D(n_9704),
.Y(n_20130)
);

O2A1O1Ixp33_ASAP7_75t_L g20131 ( 
.A1(n_19887),
.A2(n_10745),
.B(n_10775),
.C(n_10743),
.Y(n_20131)
);

OAI211xp5_ASAP7_75t_L g20132 ( 
.A1(n_19733),
.A2(n_8992),
.B(n_9199),
.C(n_12730),
.Y(n_20132)
);

AOI222xp33_ASAP7_75t_L g20133 ( 
.A1(n_19832),
.A2(n_19965),
.B1(n_19975),
.B2(n_19753),
.C1(n_20002),
.C2(n_20014),
.Y(n_20133)
);

NOR2xp33_ASAP7_75t_L g20134 ( 
.A(n_19874),
.B(n_8497),
.Y(n_20134)
);

NAND2x1p5_ASAP7_75t_L g20135 ( 
.A(n_19866),
.B(n_8504),
.Y(n_20135)
);

INVx1_ASAP7_75t_L g20136 ( 
.A(n_19850),
.Y(n_20136)
);

INVxp67_ASAP7_75t_L g20137 ( 
.A(n_19843),
.Y(n_20137)
);

AOI22xp5_ASAP7_75t_L g20138 ( 
.A1(n_19752),
.A2(n_9468),
.B1(n_9566),
.B2(n_9476),
.Y(n_20138)
);

OAI22xp33_ASAP7_75t_L g20139 ( 
.A1(n_19821),
.A2(n_10745),
.B1(n_10775),
.B2(n_10743),
.Y(n_20139)
);

INVx2_ASAP7_75t_L g20140 ( 
.A(n_19894),
.Y(n_20140)
);

AND2x2_ASAP7_75t_L g20141 ( 
.A(n_19927),
.B(n_9452),
.Y(n_20141)
);

NOR2x1p5_ASAP7_75t_L g20142 ( 
.A(n_19954),
.B(n_19934),
.Y(n_20142)
);

INVx1_ASAP7_75t_L g20143 ( 
.A(n_19880),
.Y(n_20143)
);

INVx2_ASAP7_75t_L g20144 ( 
.A(n_19901),
.Y(n_20144)
);

INVx1_ASAP7_75t_L g20145 ( 
.A(n_19913),
.Y(n_20145)
);

OAI21xp5_ASAP7_75t_SL g20146 ( 
.A1(n_19920),
.A2(n_19921),
.B(n_19936),
.Y(n_20146)
);

AOI21xp5_ASAP7_75t_L g20147 ( 
.A1(n_19717),
.A2(n_12730),
.B(n_11265),
.Y(n_20147)
);

NAND2xp5_ASAP7_75t_L g20148 ( 
.A(n_19729),
.B(n_10118),
.Y(n_20148)
);

INVx1_ASAP7_75t_L g20149 ( 
.A(n_19955),
.Y(n_20149)
);

INVx1_ASAP7_75t_L g20150 ( 
.A(n_19941),
.Y(n_20150)
);

NAND2xp5_ASAP7_75t_L g20151 ( 
.A(n_19910),
.B(n_10118),
.Y(n_20151)
);

OAI222xp33_ASAP7_75t_L g20152 ( 
.A1(n_19747),
.A2(n_9578),
.B1(n_9595),
.B2(n_9694),
.C1(n_9622),
.C2(n_9493),
.Y(n_20152)
);

INVx1_ASAP7_75t_L g20153 ( 
.A(n_19942),
.Y(n_20153)
);

INVx1_ASAP7_75t_L g20154 ( 
.A(n_19943),
.Y(n_20154)
);

AOI221xp5_ASAP7_75t_L g20155 ( 
.A1(n_19737),
.A2(n_20005),
.B1(n_19946),
.B2(n_19953),
.C(n_19948),
.Y(n_20155)
);

INVxp67_ASAP7_75t_L g20156 ( 
.A(n_19872),
.Y(n_20156)
);

INVx1_ASAP7_75t_L g20157 ( 
.A(n_19969),
.Y(n_20157)
);

NAND2xp5_ASAP7_75t_L g20158 ( 
.A(n_19907),
.B(n_10139),
.Y(n_20158)
);

OAI221xp5_ASAP7_75t_L g20159 ( 
.A1(n_19745),
.A2(n_9065),
.B1(n_9924),
.B2(n_9266),
.C(n_9261),
.Y(n_20159)
);

AND2x2_ASAP7_75t_L g20160 ( 
.A(n_19904),
.B(n_9452),
.Y(n_20160)
);

BUFx2_ASAP7_75t_L g20161 ( 
.A(n_19864),
.Y(n_20161)
);

INVx2_ASAP7_75t_L g20162 ( 
.A(n_19770),
.Y(n_20162)
);

AOI21xp5_ASAP7_75t_L g20163 ( 
.A1(n_19967),
.A2(n_11265),
.B(n_11264),
.Y(n_20163)
);

NAND2xp5_ASAP7_75t_L g20164 ( 
.A(n_19916),
.B(n_10139),
.Y(n_20164)
);

NAND2xp5_ASAP7_75t_SL g20165 ( 
.A(n_19777),
.B(n_9468),
.Y(n_20165)
);

INVx3_ASAP7_75t_L g20166 ( 
.A(n_19926),
.Y(n_20166)
);

INVx1_ASAP7_75t_L g20167 ( 
.A(n_19908),
.Y(n_20167)
);

INVx1_ASAP7_75t_SL g20168 ( 
.A(n_19828),
.Y(n_20168)
);

O2A1O1Ixp33_ASAP7_75t_SL g20169 ( 
.A1(n_19918),
.A2(n_9549),
.B(n_9568),
.C(n_9482),
.Y(n_20169)
);

AOI22xp5_ASAP7_75t_L g20170 ( 
.A1(n_19837),
.A2(n_9468),
.B1(n_9566),
.B2(n_9476),
.Y(n_20170)
);

NOR2xp33_ASAP7_75t_L g20171 ( 
.A(n_19919),
.B(n_8497),
.Y(n_20171)
);

INVx2_ASAP7_75t_L g20172 ( 
.A(n_19906),
.Y(n_20172)
);

NAND2xp5_ASAP7_75t_L g20173 ( 
.A(n_19922),
.B(n_10139),
.Y(n_20173)
);

INVx2_ASAP7_75t_L g20174 ( 
.A(n_19923),
.Y(n_20174)
);

INVx1_ASAP7_75t_L g20175 ( 
.A(n_19929),
.Y(n_20175)
);

OAI221xp5_ASAP7_75t_L g20176 ( 
.A1(n_19997),
.A2(n_9065),
.B1(n_9924),
.B2(n_9266),
.C(n_9261),
.Y(n_20176)
);

OAI22xp33_ASAP7_75t_L g20177 ( 
.A1(n_19881),
.A2(n_10775),
.B1(n_10785),
.B2(n_10745),
.Y(n_20177)
);

INVx1_ASAP7_75t_SL g20178 ( 
.A(n_19801),
.Y(n_20178)
);

INVx2_ASAP7_75t_L g20179 ( 
.A(n_19928),
.Y(n_20179)
);

INVx1_ASAP7_75t_SL g20180 ( 
.A(n_19839),
.Y(n_20180)
);

INVx1_ASAP7_75t_L g20181 ( 
.A(n_19931),
.Y(n_20181)
);

NAND2xp5_ASAP7_75t_L g20182 ( 
.A(n_19933),
.B(n_10139),
.Y(n_20182)
);

NOR2xp33_ASAP7_75t_L g20183 ( 
.A(n_19924),
.B(n_8497),
.Y(n_20183)
);

INVx2_ASAP7_75t_L g20184 ( 
.A(n_19972),
.Y(n_20184)
);

INVxp67_ASAP7_75t_L g20185 ( 
.A(n_19963),
.Y(n_20185)
);

INVx1_ASAP7_75t_SL g20186 ( 
.A(n_19842),
.Y(n_20186)
);

INVx1_ASAP7_75t_L g20187 ( 
.A(n_19959),
.Y(n_20187)
);

AOI22xp33_ASAP7_75t_SL g20188 ( 
.A1(n_19989),
.A2(n_9468),
.B1(n_9566),
.B2(n_9476),
.Y(n_20188)
);

NAND2xp5_ASAP7_75t_L g20189 ( 
.A(n_19956),
.B(n_19966),
.Y(n_20189)
);

O2A1O1Ixp33_ASAP7_75t_L g20190 ( 
.A1(n_19957),
.A2(n_10775),
.B(n_10785),
.C(n_10745),
.Y(n_20190)
);

OAI21xp5_ASAP7_75t_L g20191 ( 
.A1(n_19886),
.A2(n_10210),
.B(n_10204),
.Y(n_20191)
);

AOI21xp33_ASAP7_75t_SL g20192 ( 
.A1(n_19847),
.A2(n_9261),
.B(n_9065),
.Y(n_20192)
);

INVx1_ASAP7_75t_L g20193 ( 
.A(n_19859),
.Y(n_20193)
);

INVx2_ASAP7_75t_L g20194 ( 
.A(n_19968),
.Y(n_20194)
);

INVx1_ASAP7_75t_L g20195 ( 
.A(n_19960),
.Y(n_20195)
);

AOI21xp33_ASAP7_75t_SL g20196 ( 
.A1(n_19870),
.A2(n_19895),
.B(n_19891),
.Y(n_20196)
);

OAI321xp33_ASAP7_75t_L g20197 ( 
.A1(n_19784),
.A2(n_9994),
.A3(n_9266),
.B1(n_9924),
.B2(n_9261),
.C(n_10311),
.Y(n_20197)
);

INVx1_ASAP7_75t_L g20198 ( 
.A(n_19781),
.Y(n_20198)
);

INVx1_ASAP7_75t_L g20199 ( 
.A(n_19786),
.Y(n_20199)
);

OAI22xp5_ASAP7_75t_L g20200 ( 
.A1(n_19746),
.A2(n_9744),
.B1(n_9636),
.B2(n_9594),
.Y(n_20200)
);

AOI22xp33_ASAP7_75t_L g20201 ( 
.A1(n_19890),
.A2(n_11264),
.B1(n_11265),
.B2(n_10139),
.Y(n_20201)
);

INVx2_ASAP7_75t_SL g20202 ( 
.A(n_19889),
.Y(n_20202)
);

HB1xp67_ASAP7_75t_L g20203 ( 
.A(n_19899),
.Y(n_20203)
);

INVx2_ASAP7_75t_L g20204 ( 
.A(n_19964),
.Y(n_20204)
);

AOI22xp5_ASAP7_75t_L g20205 ( 
.A1(n_19816),
.A2(n_9476),
.B1(n_9629),
.B2(n_9566),
.Y(n_20205)
);

AOI221xp5_ASAP7_75t_L g20206 ( 
.A1(n_19973),
.A2(n_10910),
.B1(n_10936),
.B2(n_10798),
.C(n_10785),
.Y(n_20206)
);

OR2x2_ASAP7_75t_L g20207 ( 
.A(n_19911),
.B(n_10339),
.Y(n_20207)
);

NAND2xp5_ASAP7_75t_L g20208 ( 
.A(n_19980),
.B(n_10139),
.Y(n_20208)
);

INVx1_ASAP7_75t_L g20209 ( 
.A(n_19939),
.Y(n_20209)
);

INVx1_ASAP7_75t_SL g20210 ( 
.A(n_19938),
.Y(n_20210)
);

INVx1_ASAP7_75t_L g20211 ( 
.A(n_19976),
.Y(n_20211)
);

AOI21xp5_ASAP7_75t_L g20212 ( 
.A1(n_19736),
.A2(n_11265),
.B(n_11264),
.Y(n_20212)
);

INVxp67_ASAP7_75t_L g20213 ( 
.A(n_19845),
.Y(n_20213)
);

INVx1_ASAP7_75t_L g20214 ( 
.A(n_19885),
.Y(n_20214)
);

OAI21xp33_ASAP7_75t_L g20215 ( 
.A1(n_20003),
.A2(n_9594),
.B(n_9588),
.Y(n_20215)
);

AND2x4_ASAP7_75t_L g20216 ( 
.A(n_19987),
.B(n_10931),
.Y(n_20216)
);

OR2x2_ASAP7_75t_L g20217 ( 
.A(n_19996),
.B(n_10339),
.Y(n_20217)
);

OR2x2_ASAP7_75t_L g20218 ( 
.A(n_19780),
.B(n_10339),
.Y(n_20218)
);

INVxp67_ASAP7_75t_L g20219 ( 
.A(n_19977),
.Y(n_20219)
);

NAND2xp5_ASAP7_75t_L g20220 ( 
.A(n_19984),
.B(n_10139),
.Y(n_20220)
);

AOI221xp5_ASAP7_75t_L g20221 ( 
.A1(n_19998),
.A2(n_11124),
.B1(n_11105),
.B2(n_10910),
.C(n_10936),
.Y(n_20221)
);

NOR2xp33_ASAP7_75t_L g20222 ( 
.A(n_20013),
.B(n_8497),
.Y(n_20222)
);

OAI211xp5_ASAP7_75t_L g20223 ( 
.A1(n_19813),
.A2(n_9199),
.B(n_9064),
.C(n_9145),
.Y(n_20223)
);

AOI322xp5_ASAP7_75t_L g20224 ( 
.A1(n_19757),
.A2(n_9595),
.A3(n_9578),
.B1(n_9694),
.B2(n_9622),
.C1(n_9493),
.C2(n_10076),
.Y(n_20224)
);

NAND2xp5_ASAP7_75t_L g20225 ( 
.A(n_19848),
.B(n_11264),
.Y(n_20225)
);

NAND2xp5_ASAP7_75t_L g20226 ( 
.A(n_19944),
.B(n_9268),
.Y(n_20226)
);

OR2x2_ASAP7_75t_L g20227 ( 
.A(n_19826),
.B(n_19779),
.Y(n_20227)
);

NAND3xp33_ASAP7_75t_L g20228 ( 
.A(n_19902),
.B(n_9566),
.C(n_9476),
.Y(n_20228)
);

INVx2_ASAP7_75t_L g20229 ( 
.A(n_19877),
.Y(n_20229)
);

AOI21xp33_ASAP7_75t_L g20230 ( 
.A1(n_19947),
.A2(n_11326),
.B(n_11322),
.Y(n_20230)
);

INVx1_ASAP7_75t_L g20231 ( 
.A(n_19985),
.Y(n_20231)
);

INVx1_ASAP7_75t_L g20232 ( 
.A(n_19858),
.Y(n_20232)
);

NAND2xp5_ASAP7_75t_L g20233 ( 
.A(n_19759),
.B(n_9268),
.Y(n_20233)
);

OAI21xp5_ASAP7_75t_SL g20234 ( 
.A1(n_19878),
.A2(n_9266),
.B(n_9261),
.Y(n_20234)
);

OAI221xp5_ASAP7_75t_L g20235 ( 
.A1(n_19983),
.A2(n_9266),
.B1(n_9994),
.B2(n_9924),
.C(n_9549),
.Y(n_20235)
);

INVx1_ASAP7_75t_L g20236 ( 
.A(n_19978),
.Y(n_20236)
);

NAND2xp5_ASAP7_75t_L g20237 ( 
.A(n_19854),
.B(n_19738),
.Y(n_20237)
);

INVx2_ASAP7_75t_L g20238 ( 
.A(n_19873),
.Y(n_20238)
);

INVx1_ASAP7_75t_L g20239 ( 
.A(n_19764),
.Y(n_20239)
);

INVx2_ASAP7_75t_L g20240 ( 
.A(n_19962),
.Y(n_20240)
);

AND2x2_ASAP7_75t_L g20241 ( 
.A(n_19862),
.B(n_19809),
.Y(n_20241)
);

O2A1O1Ixp33_ASAP7_75t_L g20242 ( 
.A1(n_19912),
.A2(n_11133),
.B(n_10910),
.C(n_10798),
.Y(n_20242)
);

NOR2xp33_ASAP7_75t_L g20243 ( 
.A(n_19930),
.B(n_8497),
.Y(n_20243)
);

A2O1A1Ixp33_ASAP7_75t_SL g20244 ( 
.A1(n_19766),
.A2(n_9659),
.B(n_9705),
.C(n_9620),
.Y(n_20244)
);

OAI22xp33_ASAP7_75t_L g20245 ( 
.A1(n_19986),
.A2(n_20009),
.B1(n_19853),
.B2(n_19876),
.Y(n_20245)
);

OAI21xp5_ASAP7_75t_SL g20246 ( 
.A1(n_19829),
.A2(n_9994),
.B(n_9924),
.Y(n_20246)
);

INVx1_ASAP7_75t_L g20247 ( 
.A(n_19846),
.Y(n_20247)
);

OR2x2_ASAP7_75t_L g20248 ( 
.A(n_19871),
.B(n_10339),
.Y(n_20248)
);

INVx2_ASAP7_75t_L g20249 ( 
.A(n_20000),
.Y(n_20249)
);

INVx3_ASAP7_75t_L g20250 ( 
.A(n_19945),
.Y(n_20250)
);

INVx1_ASAP7_75t_SL g20251 ( 
.A(n_19811),
.Y(n_20251)
);

OAI21xp5_ASAP7_75t_L g20252 ( 
.A1(n_19867),
.A2(n_10210),
.B(n_10204),
.Y(n_20252)
);

INVxp67_ASAP7_75t_L g20253 ( 
.A(n_19856),
.Y(n_20253)
);

INVx1_ASAP7_75t_L g20254 ( 
.A(n_19914),
.Y(n_20254)
);

AND2x4_ASAP7_75t_L g20255 ( 
.A(n_19815),
.B(n_9159),
.Y(n_20255)
);

INVx1_ASAP7_75t_L g20256 ( 
.A(n_19999),
.Y(n_20256)
);

INVx1_ASAP7_75t_L g20257 ( 
.A(n_19990),
.Y(n_20257)
);

INVx1_ASAP7_75t_L g20258 ( 
.A(n_19831),
.Y(n_20258)
);

INVx1_ASAP7_75t_L g20259 ( 
.A(n_19869),
.Y(n_20259)
);

INVx3_ASAP7_75t_L g20260 ( 
.A(n_19945),
.Y(n_20260)
);

NAND2xp5_ASAP7_75t_L g20261 ( 
.A(n_19794),
.B(n_9268),
.Y(n_20261)
);

NAND2xp5_ASAP7_75t_L g20262 ( 
.A(n_19988),
.B(n_9268),
.Y(n_20262)
);

AOI222xp33_ASAP7_75t_L g20263 ( 
.A1(n_19950),
.A2(n_10936),
.B1(n_10798),
.B2(n_10947),
.C1(n_10910),
.C2(n_10785),
.Y(n_20263)
);

INVx2_ASAP7_75t_SL g20264 ( 
.A(n_19844),
.Y(n_20264)
);

INVx1_ASAP7_75t_L g20265 ( 
.A(n_19883),
.Y(n_20265)
);

INVx2_ASAP7_75t_L g20266 ( 
.A(n_19974),
.Y(n_20266)
);

AOI211x1_ASAP7_75t_SL g20267 ( 
.A1(n_20007),
.A2(n_10936),
.B(n_10947),
.C(n_10798),
.Y(n_20267)
);

NAND2xp5_ASAP7_75t_SL g20268 ( 
.A(n_19852),
.B(n_9476),
.Y(n_20268)
);

INVx2_ASAP7_75t_L g20269 ( 
.A(n_19974),
.Y(n_20269)
);

NOR2xp33_ASAP7_75t_L g20270 ( 
.A(n_19810),
.B(n_19909),
.Y(n_20270)
);

INVx1_ASAP7_75t_L g20271 ( 
.A(n_19792),
.Y(n_20271)
);

OAI21xp5_ASAP7_75t_L g20272 ( 
.A1(n_19991),
.A2(n_10224),
.B(n_10220),
.Y(n_20272)
);

AOI221xp5_ASAP7_75t_L g20273 ( 
.A1(n_19741),
.A2(n_11128),
.B1(n_11147),
.B2(n_11076),
.C(n_10947),
.Y(n_20273)
);

AND2x4_ASAP7_75t_L g20274 ( 
.A(n_19995),
.B(n_9159),
.Y(n_20274)
);

INVx1_ASAP7_75t_L g20275 ( 
.A(n_19932),
.Y(n_20275)
);

OAI21xp33_ASAP7_75t_L g20276 ( 
.A1(n_19751),
.A2(n_9602),
.B(n_9588),
.Y(n_20276)
);

INVx1_ASAP7_75t_L g20277 ( 
.A(n_19940),
.Y(n_20277)
);

AOI21xp33_ASAP7_75t_L g20278 ( 
.A1(n_19961),
.A2(n_11326),
.B(n_11322),
.Y(n_20278)
);

INVx1_ASAP7_75t_L g20279 ( 
.A(n_19750),
.Y(n_20279)
);

OR2x2_ASAP7_75t_L g20280 ( 
.A(n_20006),
.B(n_10339),
.Y(n_20280)
);

INVx1_ASAP7_75t_L g20281 ( 
.A(n_19749),
.Y(n_20281)
);

OR2x2_ASAP7_75t_L g20282 ( 
.A(n_19979),
.B(n_10339),
.Y(n_20282)
);

NAND2xp5_ASAP7_75t_L g20283 ( 
.A(n_19796),
.B(n_9268),
.Y(n_20283)
);

AOI21xp33_ASAP7_75t_SL g20284 ( 
.A1(n_19769),
.A2(n_9994),
.B(n_9924),
.Y(n_20284)
);

NAND2xp5_ASAP7_75t_L g20285 ( 
.A(n_19768),
.B(n_9268),
.Y(n_20285)
);

AND2x2_ASAP7_75t_L g20286 ( 
.A(n_19875),
.B(n_9452),
.Y(n_20286)
);

INVx1_ASAP7_75t_L g20287 ( 
.A(n_20008),
.Y(n_20287)
);

AOI221xp5_ASAP7_75t_L g20288 ( 
.A1(n_20020),
.A2(n_19840),
.B1(n_19898),
.B2(n_11090),
.C(n_11092),
.Y(n_20288)
);

INVx2_ASAP7_75t_L g20289 ( 
.A(n_20103),
.Y(n_20289)
);

INVx1_ASAP7_75t_L g20290 ( 
.A(n_20120),
.Y(n_20290)
);

OAI221xp5_ASAP7_75t_L g20291 ( 
.A1(n_20100),
.A2(n_19981),
.B1(n_9994),
.B2(n_9924),
.C(n_9568),
.Y(n_20291)
);

NAND2xp5_ASAP7_75t_SL g20292 ( 
.A(n_20048),
.B(n_9476),
.Y(n_20292)
);

AOI21xp5_ASAP7_75t_L g20293 ( 
.A1(n_20025),
.A2(n_10432),
.B(n_10403),
.Y(n_20293)
);

AOI221xp5_ASAP7_75t_L g20294 ( 
.A1(n_20033),
.A2(n_20251),
.B1(n_20032),
.B2(n_20055),
.C(n_20030),
.Y(n_20294)
);

AOI21xp5_ASAP7_75t_L g20295 ( 
.A1(n_20110),
.A2(n_10432),
.B(n_10403),
.Y(n_20295)
);

AOI22xp5_ASAP7_75t_L g20296 ( 
.A1(n_20109),
.A2(n_9629),
.B1(n_9653),
.B2(n_9566),
.Y(n_20296)
);

NOR4xp25_ASAP7_75t_L g20297 ( 
.A(n_20029),
.B(n_10077),
.C(n_10143),
.D(n_10076),
.Y(n_20297)
);

AOI22xp5_ASAP7_75t_L g20298 ( 
.A1(n_20056),
.A2(n_9629),
.B1(n_9653),
.B2(n_9566),
.Y(n_20298)
);

AOI322xp5_ASAP7_75t_L g20299 ( 
.A1(n_20027),
.A2(n_9694),
.A3(n_9622),
.B1(n_9493),
.B2(n_10077),
.C1(n_10143),
.C2(n_10076),
.Y(n_20299)
);

AOI21xp33_ASAP7_75t_L g20300 ( 
.A1(n_20114),
.A2(n_11326),
.B(n_11322),
.Y(n_20300)
);

INVx1_ASAP7_75t_L g20301 ( 
.A(n_20015),
.Y(n_20301)
);

AOI322xp5_ASAP7_75t_L g20302 ( 
.A1(n_20148),
.A2(n_9622),
.A3(n_9694),
.B1(n_10143),
.B2(n_10077),
.C1(n_10076),
.C2(n_10947),
.Y(n_20302)
);

AOI211xp5_ASAP7_75t_L g20303 ( 
.A1(n_20018),
.A2(n_9386),
.B(n_9537),
.C(n_9211),
.Y(n_20303)
);

OAI22xp33_ASAP7_75t_L g20304 ( 
.A1(n_20116),
.A2(n_11090),
.B1(n_11092),
.B2(n_11076),
.Y(n_20304)
);

AOI211xp5_ASAP7_75t_L g20305 ( 
.A1(n_20245),
.A2(n_9386),
.B(n_9537),
.C(n_9211),
.Y(n_20305)
);

AOI21xp5_ASAP7_75t_L g20306 ( 
.A1(n_20022),
.A2(n_10432),
.B(n_10403),
.Y(n_20306)
);

AOI21xp33_ASAP7_75t_L g20307 ( 
.A1(n_20059),
.A2(n_11326),
.B(n_11322),
.Y(n_20307)
);

OAI21xp5_ASAP7_75t_L g20308 ( 
.A1(n_20023),
.A2(n_20091),
.B(n_20043),
.Y(n_20308)
);

O2A1O1Ixp33_ASAP7_75t_L g20309 ( 
.A1(n_20213),
.A2(n_10093),
.B(n_10054),
.C(n_11076),
.Y(n_20309)
);

AOI22xp5_ASAP7_75t_L g20310 ( 
.A1(n_20103),
.A2(n_9629),
.B1(n_9653),
.B2(n_9566),
.Y(n_20310)
);

AOI21xp5_ASAP7_75t_L g20311 ( 
.A1(n_20024),
.A2(n_10432),
.B(n_10403),
.Y(n_20311)
);

OR2x2_ASAP7_75t_L g20312 ( 
.A(n_20135),
.B(n_10546),
.Y(n_20312)
);

INVx1_ASAP7_75t_L g20313 ( 
.A(n_20260),
.Y(n_20313)
);

AOI22xp33_ASAP7_75t_L g20314 ( 
.A1(n_20130),
.A2(n_10991),
.B1(n_9653),
.B2(n_9658),
.Y(n_20314)
);

AOI22xp5_ASAP7_75t_L g20315 ( 
.A1(n_20081),
.A2(n_20113),
.B1(n_20149),
.B2(n_20090),
.Y(n_20315)
);

AOI21xp5_ASAP7_75t_SL g20316 ( 
.A1(n_20266),
.A2(n_10180),
.B(n_9377),
.Y(n_20316)
);

AOI221xp5_ASAP7_75t_L g20317 ( 
.A1(n_20256),
.A2(n_11076),
.B1(n_11101),
.B2(n_11092),
.C(n_11090),
.Y(n_20317)
);

OAI22xp5_ASAP7_75t_L g20318 ( 
.A1(n_20099),
.A2(n_9602),
.B1(n_9618),
.B2(n_9588),
.Y(n_20318)
);

INVx1_ASAP7_75t_L g20319 ( 
.A(n_20260),
.Y(n_20319)
);

INVxp33_ASAP7_75t_L g20320 ( 
.A(n_20021),
.Y(n_20320)
);

OAI21xp5_ASAP7_75t_SL g20321 ( 
.A1(n_20146),
.A2(n_9994),
.B(n_9659),
.Y(n_20321)
);

INVxp67_ASAP7_75t_L g20322 ( 
.A(n_20049),
.Y(n_20322)
);

NOR3xp33_ASAP7_75t_L g20323 ( 
.A(n_20052),
.B(n_8088),
.C(n_8020),
.Y(n_20323)
);

OAI21xp5_ASAP7_75t_L g20324 ( 
.A1(n_20137),
.A2(n_10224),
.B(n_10220),
.Y(n_20324)
);

INVx1_ASAP7_75t_L g20325 ( 
.A(n_20250),
.Y(n_20325)
);

NAND2xp5_ASAP7_75t_SL g20326 ( 
.A(n_20039),
.B(n_9629),
.Y(n_20326)
);

AOI21xp33_ASAP7_75t_SL g20327 ( 
.A1(n_20257),
.A2(n_9994),
.B(n_10403),
.Y(n_20327)
);

OAI21xp5_ASAP7_75t_SL g20328 ( 
.A1(n_20031),
.A2(n_9659),
.B(n_9620),
.Y(n_20328)
);

AOI22xp5_ASAP7_75t_L g20329 ( 
.A1(n_20183),
.A2(n_9653),
.B1(n_9658),
.B2(n_9629),
.Y(n_20329)
);

AOI21xp5_ASAP7_75t_L g20330 ( 
.A1(n_20232),
.A2(n_10432),
.B(n_10403),
.Y(n_20330)
);

AOI22xp5_ASAP7_75t_L g20331 ( 
.A1(n_20134),
.A2(n_9653),
.B1(n_9658),
.B2(n_9629),
.Y(n_20331)
);

AOI221x1_ASAP7_75t_L g20332 ( 
.A1(n_20028),
.A2(n_9602),
.B1(n_9632),
.B2(n_9623),
.C(n_9618),
.Y(n_20332)
);

INVx1_ASAP7_75t_L g20333 ( 
.A(n_20141),
.Y(n_20333)
);

OAI22xp5_ASAP7_75t_L g20334 ( 
.A1(n_20047),
.A2(n_9618),
.B1(n_9632),
.B2(n_9623),
.Y(n_20334)
);

AOI221xp5_ASAP7_75t_L g20335 ( 
.A1(n_20155),
.A2(n_20281),
.B1(n_20196),
.B2(n_20287),
.C(n_20038),
.Y(n_20335)
);

NAND2xp5_ASAP7_75t_SL g20336 ( 
.A(n_20060),
.B(n_9629),
.Y(n_20336)
);

INVx1_ASAP7_75t_L g20337 ( 
.A(n_20126),
.Y(n_20337)
);

OAI22xp5_ASAP7_75t_L g20338 ( 
.A1(n_20050),
.A2(n_20157),
.B1(n_20097),
.B2(n_20143),
.Y(n_20338)
);

OAI22x1_ASAP7_75t_L g20339 ( 
.A1(n_20142),
.A2(n_9145),
.B1(n_9064),
.B2(n_9636),
.Y(n_20339)
);

AOI211xp5_ASAP7_75t_L g20340 ( 
.A1(n_20053),
.A2(n_9537),
.B(n_9766),
.C(n_9717),
.Y(n_20340)
);

INVx1_ASAP7_75t_L g20341 ( 
.A(n_20036),
.Y(n_20341)
);

OAI221xp5_ASAP7_75t_SL g20342 ( 
.A1(n_20045),
.A2(n_20276),
.B1(n_20246),
.B2(n_20062),
.C(n_20019),
.Y(n_20342)
);

AOI22xp5_ASAP7_75t_L g20343 ( 
.A1(n_20243),
.A2(n_9653),
.B1(n_9658),
.B2(n_9629),
.Y(n_20343)
);

OAI211xp5_ASAP7_75t_SL g20344 ( 
.A1(n_20156),
.A2(n_9659),
.B(n_9705),
.C(n_9620),
.Y(n_20344)
);

OAI21xp33_ASAP7_75t_L g20345 ( 
.A1(n_20171),
.A2(n_9623),
.B(n_9618),
.Y(n_20345)
);

AOI21xp5_ASAP7_75t_L g20346 ( 
.A1(n_20239),
.A2(n_10440),
.B(n_10432),
.Y(n_20346)
);

AOI322xp5_ASAP7_75t_L g20347 ( 
.A1(n_20061),
.A2(n_10143),
.A3(n_10077),
.B1(n_11092),
.B2(n_11101),
.C1(n_11105),
.C2(n_11090),
.Y(n_20347)
);

AND2x2_ASAP7_75t_L g20348 ( 
.A(n_20112),
.B(n_20136),
.Y(n_20348)
);

O2A1O1Ixp5_ASAP7_75t_L g20349 ( 
.A1(n_20269),
.A2(n_10311),
.B(n_10254),
.C(n_10266),
.Y(n_20349)
);

O2A1O1Ixp33_ASAP7_75t_SL g20350 ( 
.A1(n_20210),
.A2(n_9124),
.B(n_9038),
.C(n_9482),
.Y(n_20350)
);

NOR2xp33_ASAP7_75t_L g20351 ( 
.A(n_20068),
.B(n_8497),
.Y(n_20351)
);

NAND3xp33_ASAP7_75t_L g20352 ( 
.A(n_20259),
.B(n_9653),
.C(n_9629),
.Y(n_20352)
);

NOR2xp33_ASAP7_75t_L g20353 ( 
.A(n_20044),
.B(n_8497),
.Y(n_20353)
);

AOI222xp33_ASAP7_75t_L g20354 ( 
.A1(n_20258),
.A2(n_11124),
.B1(n_11101),
.B2(n_11125),
.C1(n_11119),
.C2(n_11105),
.Y(n_20354)
);

NAND3xp33_ASAP7_75t_L g20355 ( 
.A(n_20271),
.B(n_9653),
.C(n_9629),
.Y(n_20355)
);

OAI22xp33_ASAP7_75t_SL g20356 ( 
.A1(n_20211),
.A2(n_20265),
.B1(n_20064),
.B2(n_20231),
.Y(n_20356)
);

INVx1_ASAP7_75t_L g20357 ( 
.A(n_20074),
.Y(n_20357)
);

OAI221xp5_ASAP7_75t_L g20358 ( 
.A1(n_20083),
.A2(n_9568),
.B1(n_9613),
.B2(n_9598),
.C(n_9549),
.Y(n_20358)
);

NAND4xp25_ASAP7_75t_L g20359 ( 
.A(n_20133),
.B(n_8088),
.C(n_8460),
.D(n_8020),
.Y(n_20359)
);

OAI21xp5_ASAP7_75t_L g20360 ( 
.A1(n_20041),
.A2(n_10224),
.B(n_10220),
.Y(n_20360)
);

OAI21xp5_ASAP7_75t_SL g20361 ( 
.A1(n_20071),
.A2(n_9659),
.B(n_9620),
.Y(n_20361)
);

INVx1_ASAP7_75t_L g20362 ( 
.A(n_20104),
.Y(n_20362)
);

INVxp67_ASAP7_75t_L g20363 ( 
.A(n_20105),
.Y(n_20363)
);

AOI22xp5_ASAP7_75t_L g20364 ( 
.A1(n_20058),
.A2(n_9653),
.B1(n_9658),
.B2(n_9629),
.Y(n_20364)
);

AOI22xp33_ASAP7_75t_SL g20365 ( 
.A1(n_20016),
.A2(n_9653),
.B1(n_9658),
.B2(n_9629),
.Y(n_20365)
);

INVx1_ASAP7_75t_L g20366 ( 
.A(n_20115),
.Y(n_20366)
);

INVx1_ASAP7_75t_L g20367 ( 
.A(n_20123),
.Y(n_20367)
);

AOI222xp33_ASAP7_75t_L g20368 ( 
.A1(n_20253),
.A2(n_11124),
.B1(n_11101),
.B2(n_11125),
.C1(n_11119),
.C2(n_11105),
.Y(n_20368)
);

NOR3xp33_ASAP7_75t_L g20369 ( 
.A(n_20145),
.B(n_20185),
.C(n_20026),
.Y(n_20369)
);

OAI21xp5_ASAP7_75t_SL g20370 ( 
.A1(n_20160),
.A2(n_9705),
.B(n_9620),
.Y(n_20370)
);

AOI21xp5_ASAP7_75t_L g20371 ( 
.A1(n_20237),
.A2(n_10440),
.B(n_11534),
.Y(n_20371)
);

OAI221xp5_ASAP7_75t_L g20372 ( 
.A1(n_20017),
.A2(n_9568),
.B1(n_9613),
.B2(n_9598),
.C(n_9549),
.Y(n_20372)
);

AOI22xp5_ASAP7_75t_L g20373 ( 
.A1(n_20150),
.A2(n_9658),
.B1(n_9688),
.B2(n_9653),
.Y(n_20373)
);

INVx1_ASAP7_75t_L g20374 ( 
.A(n_20153),
.Y(n_20374)
);

NAND4xp25_ASAP7_75t_SL g20375 ( 
.A(n_20034),
.B(n_20073),
.C(n_20195),
.D(n_20121),
.Y(n_20375)
);

AOI21xp33_ASAP7_75t_L g20376 ( 
.A1(n_20154),
.A2(n_11326),
.B(n_11322),
.Y(n_20376)
);

OAI21xp5_ASAP7_75t_L g20377 ( 
.A1(n_20270),
.A2(n_10249),
.B(n_11252),
.Y(n_20377)
);

AOI221xp5_ASAP7_75t_L g20378 ( 
.A1(n_20200),
.A2(n_11125),
.B1(n_11128),
.B2(n_11124),
.C(n_11119),
.Y(n_20378)
);

OAI22xp33_ASAP7_75t_L g20379 ( 
.A1(n_20280),
.A2(n_11125),
.B1(n_11128),
.B2(n_11119),
.Y(n_20379)
);

OAI21xp33_ASAP7_75t_SL g20380 ( 
.A1(n_20057),
.A2(n_10659),
.B(n_10639),
.Y(n_20380)
);

AOI22xp5_ASAP7_75t_L g20381 ( 
.A1(n_20264),
.A2(n_9658),
.B1(n_9688),
.B2(n_9653),
.Y(n_20381)
);

OAI21xp5_ASAP7_75t_L g20382 ( 
.A1(n_20241),
.A2(n_10249),
.B(n_11381),
.Y(n_20382)
);

OR2x2_ASAP7_75t_L g20383 ( 
.A(n_20107),
.B(n_10546),
.Y(n_20383)
);

AOI21xp5_ASAP7_75t_L g20384 ( 
.A1(n_20178),
.A2(n_10440),
.B(n_11534),
.Y(n_20384)
);

O2A1O1Ixp33_ASAP7_75t_L g20385 ( 
.A1(n_20238),
.A2(n_10093),
.B(n_10054),
.C(n_11128),
.Y(n_20385)
);

INVx1_ASAP7_75t_L g20386 ( 
.A(n_20069),
.Y(n_20386)
);

AOI21xp33_ASAP7_75t_L g20387 ( 
.A1(n_20168),
.A2(n_11326),
.B(n_11322),
.Y(n_20387)
);

NAND2xp5_ASAP7_75t_L g20388 ( 
.A(n_20098),
.B(n_9412),
.Y(n_20388)
);

AOI322xp5_ASAP7_75t_L g20389 ( 
.A1(n_20279),
.A2(n_11149),
.A3(n_11134),
.B1(n_11147),
.B2(n_11133),
.C1(n_9725),
.C2(n_9704),
.Y(n_20389)
);

O2A1O1Ixp33_ASAP7_75t_SL g20390 ( 
.A1(n_20277),
.A2(n_9124),
.B(n_9038),
.C(n_9549),
.Y(n_20390)
);

OAI21xp33_ASAP7_75t_L g20391 ( 
.A1(n_20222),
.A2(n_9632),
.B(n_9623),
.Y(n_20391)
);

AOI322xp5_ASAP7_75t_L g20392 ( 
.A1(n_20167),
.A2(n_11149),
.A3(n_11134),
.B1(n_11147),
.B2(n_11133),
.C1(n_9806),
.C2(n_9704),
.Y(n_20392)
);

INVx1_ASAP7_75t_L g20393 ( 
.A(n_20124),
.Y(n_20393)
);

AOI21xp33_ASAP7_75t_L g20394 ( 
.A1(n_20202),
.A2(n_10440),
.B(n_9971),
.Y(n_20394)
);

INVx1_ASAP7_75t_L g20395 ( 
.A(n_20140),
.Y(n_20395)
);

AOI211x1_ASAP7_75t_L g20396 ( 
.A1(n_20215),
.A2(n_11047),
.B(n_11069),
.C(n_11562),
.Y(n_20396)
);

AOI21xp5_ASAP7_75t_L g20397 ( 
.A1(n_20189),
.A2(n_10440),
.B(n_11534),
.Y(n_20397)
);

OAI21xp33_ASAP7_75t_L g20398 ( 
.A1(n_20095),
.A2(n_9634),
.B(n_9632),
.Y(n_20398)
);

NAND5xp2_ASAP7_75t_L g20399 ( 
.A(n_20175),
.B(n_8762),
.C(n_9289),
.D(n_9027),
.E(n_8783),
.Y(n_20399)
);

NAND2xp5_ASAP7_75t_SL g20400 ( 
.A(n_20054),
.B(n_20067),
.Y(n_20400)
);

AOI221xp5_ASAP7_75t_L g20401 ( 
.A1(n_20072),
.A2(n_11134),
.B1(n_11149),
.B2(n_11147),
.C(n_11133),
.Y(n_20401)
);

INVx1_ASAP7_75t_L g20402 ( 
.A(n_20144),
.Y(n_20402)
);

OAI22xp5_ASAP7_75t_L g20403 ( 
.A1(n_20138),
.A2(n_9634),
.B1(n_11134),
.B2(n_11149),
.Y(n_20403)
);

OAI322xp33_ASAP7_75t_L g20404 ( 
.A1(n_20219),
.A2(n_10260),
.A3(n_10273),
.B1(n_10264),
.B2(n_10294),
.C1(n_10293),
.C2(n_10282),
.Y(n_20404)
);

OAI22xp33_ASAP7_75t_SL g20405 ( 
.A1(n_20065),
.A2(n_9634),
.B1(n_9598),
.B2(n_9613),
.Y(n_20405)
);

NAND2xp5_ASAP7_75t_L g20406 ( 
.A(n_20172),
.B(n_9412),
.Y(n_20406)
);

AOI22xp5_ASAP7_75t_L g20407 ( 
.A1(n_20181),
.A2(n_9688),
.B1(n_9726),
.B2(n_9658),
.Y(n_20407)
);

OAI221xp5_ASAP7_75t_L g20408 ( 
.A1(n_20040),
.A2(n_20234),
.B1(n_20180),
.B2(n_20186),
.C(n_20051),
.Y(n_20408)
);

INVx1_ASAP7_75t_L g20409 ( 
.A(n_20174),
.Y(n_20409)
);

OAI21xp5_ASAP7_75t_SL g20410 ( 
.A1(n_20179),
.A2(n_9705),
.B(n_9620),
.Y(n_20410)
);

OAI221xp5_ASAP7_75t_L g20411 ( 
.A1(n_20184),
.A2(n_9598),
.B1(n_9637),
.B2(n_9613),
.C(n_9568),
.Y(n_20411)
);

OAI221xp5_ASAP7_75t_L g20412 ( 
.A1(n_20247),
.A2(n_9613),
.B1(n_9637),
.B2(n_9598),
.C(n_9537),
.Y(n_20412)
);

OAI211xp5_ASAP7_75t_L g20413 ( 
.A1(n_20236),
.A2(n_9064),
.B(n_9124),
.C(n_9038),
.Y(n_20413)
);

OA33x2_ASAP7_75t_L g20414 ( 
.A1(n_20122),
.A2(n_12372),
.A3(n_12591),
.B1(n_12528),
.B2(n_11690),
.B3(n_11710),
.Y(n_20414)
);

O2A1O1Ixp33_ASAP7_75t_L g20415 ( 
.A1(n_20204),
.A2(n_10093),
.B(n_10054),
.C(n_9719),
.Y(n_20415)
);

OAI21xp5_ASAP7_75t_L g20416 ( 
.A1(n_20076),
.A2(n_10249),
.B(n_11381),
.Y(n_20416)
);

NAND2xp5_ASAP7_75t_L g20417 ( 
.A(n_20084),
.B(n_20092),
.Y(n_20417)
);

INVxp33_ASAP7_75t_L g20418 ( 
.A(n_20203),
.Y(n_20418)
);

AOI222xp33_ASAP7_75t_L g20419 ( 
.A1(n_20268),
.A2(n_9634),
.B1(n_10995),
.B2(n_11015),
.C1(n_10993),
.C2(n_10982),
.Y(n_20419)
);

OAI221xp5_ASAP7_75t_L g20420 ( 
.A1(n_20254),
.A2(n_9637),
.B1(n_9377),
.B2(n_9333),
.C(n_9064),
.Y(n_20420)
);

INVxp67_ASAP7_75t_L g20421 ( 
.A(n_20249),
.Y(n_20421)
);

OAI21xp33_ASAP7_75t_L g20422 ( 
.A1(n_20096),
.A2(n_9637),
.B(n_8484),
.Y(n_20422)
);

OAI22xp5_ASAP7_75t_L g20423 ( 
.A1(n_20205),
.A2(n_10294),
.B1(n_10375),
.B2(n_10273),
.Y(n_20423)
);

O2A1O1Ixp33_ASAP7_75t_SL g20424 ( 
.A1(n_20275),
.A2(n_9637),
.B(n_9806),
.C(n_9725),
.Y(n_20424)
);

INVx1_ASAP7_75t_L g20425 ( 
.A(n_20162),
.Y(n_20425)
);

OAI22xp33_ASAP7_75t_L g20426 ( 
.A1(n_20125),
.A2(n_9688),
.B1(n_9726),
.B2(n_9658),
.Y(n_20426)
);

A2O1A1Ixp33_ASAP7_75t_L g20427 ( 
.A1(n_20229),
.A2(n_10751),
.B(n_10756),
.C(n_10755),
.Y(n_20427)
);

INVx1_ASAP7_75t_SL g20428 ( 
.A(n_20161),
.Y(n_20428)
);

OAI322xp33_ASAP7_75t_L g20429 ( 
.A1(n_20037),
.A2(n_10264),
.A3(n_10282),
.B1(n_10273),
.B2(n_10294),
.C1(n_10293),
.C2(n_10260),
.Y(n_20429)
);

AOI22xp5_ASAP7_75t_L g20430 ( 
.A1(n_20079),
.A2(n_9688),
.B1(n_9726),
.B2(n_9658),
.Y(n_20430)
);

OAI221xp5_ASAP7_75t_L g20431 ( 
.A1(n_20127),
.A2(n_9377),
.B1(n_9333),
.B2(n_9841),
.C(n_9736),
.Y(n_20431)
);

INVx1_ASAP7_75t_L g20432 ( 
.A(n_20194),
.Y(n_20432)
);

OAI221xp5_ASAP7_75t_L g20433 ( 
.A1(n_20151),
.A2(n_9377),
.B1(n_9333),
.B2(n_9841),
.C(n_9736),
.Y(n_20433)
);

AOI21xp5_ASAP7_75t_R g20434 ( 
.A1(n_20128),
.A2(n_9066),
.B(n_9058),
.Y(n_20434)
);

AOI221xp5_ASAP7_75t_SL g20435 ( 
.A1(n_20214),
.A2(n_10282),
.B1(n_10293),
.B2(n_10264),
.C(n_10260),
.Y(n_20435)
);

O2A1O1Ixp5_ASAP7_75t_SL g20436 ( 
.A1(n_20187),
.A2(n_9730),
.B(n_9748),
.C(n_9754),
.Y(n_20436)
);

AND2x2_ASAP7_75t_L g20437 ( 
.A(n_20240),
.B(n_9490),
.Y(n_20437)
);

AOI221xp5_ASAP7_75t_L g20438 ( 
.A1(n_20199),
.A2(n_9658),
.B1(n_9799),
.B2(n_9726),
.C(n_9688),
.Y(n_20438)
);

NAND2xp5_ASAP7_75t_L g20439 ( 
.A(n_20193),
.B(n_9412),
.Y(n_20439)
);

AOI22xp33_ASAP7_75t_L g20440 ( 
.A1(n_20066),
.A2(n_10991),
.B1(n_9688),
.B2(n_9726),
.Y(n_20440)
);

NAND3xp33_ASAP7_75t_L g20441 ( 
.A(n_20198),
.B(n_9688),
.C(n_9658),
.Y(n_20441)
);

INVx1_ASAP7_75t_L g20442 ( 
.A(n_20227),
.Y(n_20442)
);

AOI22xp33_ASAP7_75t_L g20443 ( 
.A1(n_20286),
.A2(n_10991),
.B1(n_9726),
.B2(n_9799),
.Y(n_20443)
);

AOI22xp5_ASAP7_75t_L g20444 ( 
.A1(n_20188),
.A2(n_9726),
.B1(n_9799),
.B2(n_9688),
.Y(n_20444)
);

INVx1_ASAP7_75t_L g20445 ( 
.A(n_20209),
.Y(n_20445)
);

AOI222xp33_ASAP7_75t_L g20446 ( 
.A1(n_20228),
.A2(n_11015),
.B1(n_10993),
.B2(n_11019),
.C1(n_10995),
.C2(n_10982),
.Y(n_20446)
);

OAI31xp33_ASAP7_75t_L g20447 ( 
.A1(n_20166),
.A2(n_9806),
.A3(n_9844),
.B(n_9725),
.Y(n_20447)
);

NAND2xp5_ASAP7_75t_L g20448 ( 
.A(n_20158),
.B(n_9412),
.Y(n_20448)
);

INVx1_ASAP7_75t_L g20449 ( 
.A(n_20118),
.Y(n_20449)
);

OAI21xp33_ASAP7_75t_L g20450 ( 
.A1(n_20164),
.A2(n_8484),
.B(n_8442),
.Y(n_20450)
);

OAI32xp33_ASAP7_75t_L g20451 ( 
.A1(n_20082),
.A2(n_10380),
.A3(n_10399),
.B1(n_10375),
.B2(n_10374),
.Y(n_20451)
);

OAI221xp5_ASAP7_75t_SL g20452 ( 
.A1(n_20173),
.A2(n_9866),
.B1(n_10019),
.B2(n_9844),
.C(n_9806),
.Y(n_20452)
);

AOI211xp5_ASAP7_75t_L g20453 ( 
.A1(n_20182),
.A2(n_9688),
.B(n_9799),
.C(n_9726),
.Y(n_20453)
);

AOI22xp5_ASAP7_75t_L g20454 ( 
.A1(n_20165),
.A2(n_9726),
.B1(n_9799),
.B2(n_9688),
.Y(n_20454)
);

NOR3xp33_ASAP7_75t_L g20455 ( 
.A(n_20119),
.B(n_8088),
.C(n_8020),
.Y(n_20455)
);

AOI22xp5_ASAP7_75t_L g20456 ( 
.A1(n_20063),
.A2(n_9726),
.B1(n_9799),
.B2(n_9688),
.Y(n_20456)
);

OAI22xp33_ASAP7_75t_SL g20457 ( 
.A1(n_20217),
.A2(n_10375),
.B1(n_10380),
.B2(n_10374),
.Y(n_20457)
);

NOR2xp33_ASAP7_75t_L g20458 ( 
.A(n_20262),
.B(n_8504),
.Y(n_20458)
);

INVx1_ASAP7_75t_L g20459 ( 
.A(n_20267),
.Y(n_20459)
);

OAI21xp5_ASAP7_75t_L g20460 ( 
.A1(n_20212),
.A2(n_20147),
.B(n_20163),
.Y(n_20460)
);

AOI211xp5_ASAP7_75t_L g20461 ( 
.A1(n_20192),
.A2(n_9688),
.B(n_9799),
.C(n_9726),
.Y(n_20461)
);

AOI21xp5_ASAP7_75t_L g20462 ( 
.A1(n_20233),
.A2(n_10440),
.B(n_11534),
.Y(n_20462)
);

INVx1_ASAP7_75t_L g20463 ( 
.A(n_20225),
.Y(n_20463)
);

AND2x4_ASAP7_75t_L g20464 ( 
.A(n_20274),
.B(n_11047),
.Y(n_20464)
);

NAND3xp33_ASAP7_75t_L g20465 ( 
.A(n_20201),
.B(n_20106),
.C(n_20284),
.Y(n_20465)
);

NAND2xp5_ASAP7_75t_L g20466 ( 
.A(n_20274),
.B(n_9412),
.Y(n_20466)
);

INVx1_ASAP7_75t_L g20467 ( 
.A(n_20261),
.Y(n_20467)
);

INVx2_ASAP7_75t_L g20468 ( 
.A(n_20207),
.Y(n_20468)
);

AOI321xp33_ASAP7_75t_L g20469 ( 
.A1(n_20235),
.A2(n_8702),
.A3(n_9066),
.B1(n_7779),
.B2(n_7918),
.C(n_9571),
.Y(n_20469)
);

AOI221xp5_ASAP7_75t_L g20470 ( 
.A1(n_20077),
.A2(n_9836),
.B1(n_9799),
.B2(n_9726),
.C(n_10982),
.Y(n_20470)
);

INVx1_ASAP7_75t_L g20471 ( 
.A(n_20282),
.Y(n_20471)
);

OAI21xp5_ASAP7_75t_SL g20472 ( 
.A1(n_20129),
.A2(n_20132),
.B(n_20208),
.Y(n_20472)
);

OAI21xp33_ASAP7_75t_L g20473 ( 
.A1(n_20086),
.A2(n_8484),
.B(n_8442),
.Y(n_20473)
);

NOR2xp67_ASAP7_75t_L g20474 ( 
.A(n_20087),
.B(n_7869),
.Y(n_20474)
);

OAI22xp5_ASAP7_75t_L g20475 ( 
.A1(n_20159),
.A2(n_10380),
.B1(n_10650),
.B2(n_10449),
.Y(n_20475)
);

AOI22xp5_ASAP7_75t_L g20476 ( 
.A1(n_20220),
.A2(n_9799),
.B1(n_9836),
.B2(n_9726),
.Y(n_20476)
);

OAI211xp5_ASAP7_75t_L g20477 ( 
.A1(n_20244),
.A2(n_11534),
.B(n_9744),
.C(n_10311),
.Y(n_20477)
);

OAI21xp5_ASAP7_75t_SL g20478 ( 
.A1(n_20089),
.A2(n_9705),
.B(n_9620),
.Y(n_20478)
);

NOR2xp33_ASAP7_75t_L g20479 ( 
.A(n_20176),
.B(n_8612),
.Y(n_20479)
);

AOI21xp5_ASAP7_75t_L g20480 ( 
.A1(n_20283),
.A2(n_20285),
.B(n_20169),
.Y(n_20480)
);

INVx1_ASAP7_75t_L g20481 ( 
.A(n_20218),
.Y(n_20481)
);

INVx1_ASAP7_75t_L g20482 ( 
.A(n_20226),
.Y(n_20482)
);

INVx1_ASAP7_75t_L g20483 ( 
.A(n_20248),
.Y(n_20483)
);

INVxp67_ASAP7_75t_L g20484 ( 
.A(n_20216),
.Y(n_20484)
);

OAI221xp5_ASAP7_75t_L g20485 ( 
.A1(n_20078),
.A2(n_20094),
.B1(n_20093),
.B2(n_20131),
.C(n_20170),
.Y(n_20485)
);

AOI22xp5_ASAP7_75t_L g20486 ( 
.A1(n_20177),
.A2(n_9836),
.B1(n_9799),
.B2(n_9705),
.Y(n_20486)
);

AOI22xp5_ASAP7_75t_L g20487 ( 
.A1(n_20046),
.A2(n_20255),
.B1(n_20216),
.B2(n_20139),
.Y(n_20487)
);

AOI221xp5_ASAP7_75t_L g20488 ( 
.A1(n_20108),
.A2(n_9799),
.B1(n_9836),
.B2(n_10995),
.C(n_10993),
.Y(n_20488)
);

AOI211xp5_ASAP7_75t_SL g20489 ( 
.A1(n_20197),
.A2(n_20088),
.B(n_20230),
.C(n_20101),
.Y(n_20489)
);

AOI21xp5_ASAP7_75t_L g20490 ( 
.A1(n_20080),
.A2(n_11534),
.B(n_10303),
.Y(n_20490)
);

OAI32xp33_ASAP7_75t_L g20491 ( 
.A1(n_20278),
.A2(n_10374),
.A3(n_10468),
.B1(n_10449),
.B2(n_10399),
.Y(n_20491)
);

OAI321xp33_ASAP7_75t_L g20492 ( 
.A1(n_20252),
.A2(n_9836),
.A3(n_9799),
.B1(n_11564),
.B2(n_11562),
.C(n_11477),
.Y(n_20492)
);

A2O1A1Ixp33_ASAP7_75t_L g20493 ( 
.A1(n_20224),
.A2(n_10751),
.B(n_10756),
.C(n_10755),
.Y(n_20493)
);

A2O1A1Ixp33_ASAP7_75t_L g20494 ( 
.A1(n_20242),
.A2(n_10751),
.B(n_10756),
.C(n_10755),
.Y(n_20494)
);

INVx1_ASAP7_75t_L g20495 ( 
.A(n_20070),
.Y(n_20495)
);

NAND2xp5_ASAP7_75t_L g20496 ( 
.A(n_20255),
.B(n_9412),
.Y(n_20496)
);

BUFx2_ASAP7_75t_L g20497 ( 
.A(n_20191),
.Y(n_20497)
);

OAI222xp33_ASAP7_75t_L g20498 ( 
.A1(n_20117),
.A2(n_9844),
.B1(n_9866),
.B2(n_10019),
.C1(n_11019),
.C2(n_11015),
.Y(n_20498)
);

AOI211xp5_ASAP7_75t_L g20499 ( 
.A1(n_20152),
.A2(n_9799),
.B(n_9836),
.C(n_9524),
.Y(n_20499)
);

AOI221xp5_ASAP7_75t_L g20500 ( 
.A1(n_20190),
.A2(n_9836),
.B1(n_11029),
.B2(n_11024),
.C(n_11019),
.Y(n_20500)
);

AOI221xp5_ASAP7_75t_L g20501 ( 
.A1(n_20223),
.A2(n_9836),
.B1(n_11060),
.B2(n_11029),
.C(n_11024),
.Y(n_20501)
);

OAI21xp33_ASAP7_75t_L g20502 ( 
.A1(n_20042),
.A2(n_8484),
.B(n_8442),
.Y(n_20502)
);

AOI21xp33_ASAP7_75t_L g20503 ( 
.A1(n_20272),
.A2(n_9971),
.B(n_9981),
.Y(n_20503)
);

NAND4xp25_ASAP7_75t_L g20504 ( 
.A(n_20221),
.B(n_8517),
.C(n_8460),
.D(n_8758),
.Y(n_20504)
);

AOI221xp5_ASAP7_75t_SL g20505 ( 
.A1(n_20206),
.A2(n_10468),
.B1(n_10634),
.B2(n_10449),
.C(n_10399),
.Y(n_20505)
);

NAND2xp5_ASAP7_75t_L g20506 ( 
.A(n_20075),
.B(n_9412),
.Y(n_20506)
);

AOI22xp5_ASAP7_75t_L g20507 ( 
.A1(n_20102),
.A2(n_9836),
.B1(n_9705),
.B2(n_9747),
.Y(n_20507)
);

AOI21xp33_ASAP7_75t_SL g20508 ( 
.A1(n_20111),
.A2(n_9971),
.B(n_10054),
.Y(n_20508)
);

AND2x2_ASAP7_75t_L g20509 ( 
.A(n_20035),
.B(n_9490),
.Y(n_20509)
);

AOI22xp5_ASAP7_75t_L g20510 ( 
.A1(n_20273),
.A2(n_9836),
.B1(n_9705),
.B2(n_9747),
.Y(n_20510)
);

INVx2_ASAP7_75t_L g20511 ( 
.A(n_20085),
.Y(n_20511)
);

AOI21xp33_ASAP7_75t_L g20512 ( 
.A1(n_20263),
.A2(n_9971),
.B(n_9981),
.Y(n_20512)
);

INVx1_ASAP7_75t_L g20513 ( 
.A(n_20120),
.Y(n_20513)
);

AOI221xp5_ASAP7_75t_L g20514 ( 
.A1(n_20020),
.A2(n_9836),
.B1(n_11060),
.B2(n_11029),
.C(n_11024),
.Y(n_20514)
);

OAI211xp5_ASAP7_75t_L g20515 ( 
.A1(n_20100),
.A2(n_9744),
.B(n_11069),
.C(n_11047),
.Y(n_20515)
);

NAND2xp5_ASAP7_75t_SL g20516 ( 
.A(n_20048),
.B(n_9836),
.Y(n_20516)
);

NAND2xp33_ASAP7_75t_L g20517 ( 
.A(n_20048),
.B(n_9836),
.Y(n_20517)
);

AOI21xp5_ASAP7_75t_L g20518 ( 
.A1(n_20025),
.A2(n_10303),
.B(n_11209),
.Y(n_20518)
);

OAI22xp5_ASAP7_75t_L g20519 ( 
.A1(n_20055),
.A2(n_10634),
.B1(n_10636),
.B2(n_10468),
.Y(n_20519)
);

AOI21xp33_ASAP7_75t_L g20520 ( 
.A1(n_20030),
.A2(n_9971),
.B(n_9981),
.Y(n_20520)
);

A2O1A1Ixp33_ASAP7_75t_L g20521 ( 
.A1(n_20109),
.A2(n_10757),
.B(n_10663),
.C(n_10621),
.Y(n_20521)
);

AOI211xp5_ASAP7_75t_SL g20522 ( 
.A1(n_20055),
.A2(n_9727),
.B(n_9752),
.C(n_9747),
.Y(n_20522)
);

AOI21xp5_ASAP7_75t_L g20523 ( 
.A1(n_20025),
.A2(n_10303),
.B(n_11209),
.Y(n_20523)
);

XNOR2xp5_ASAP7_75t_L g20524 ( 
.A(n_20024),
.B(n_9333),
.Y(n_20524)
);

BUFx2_ASAP7_75t_L g20525 ( 
.A(n_20135),
.Y(n_20525)
);

NAND2x1_ASAP7_75t_L g20526 ( 
.A(n_20260),
.B(n_9719),
.Y(n_20526)
);

INVx1_ASAP7_75t_L g20527 ( 
.A(n_20120),
.Y(n_20527)
);

AOI32xp33_ASAP7_75t_L g20528 ( 
.A1(n_20027),
.A2(n_9747),
.A3(n_9752),
.B1(n_9727),
.B2(n_9844),
.Y(n_20528)
);

NAND2xp5_ASAP7_75t_SL g20529 ( 
.A(n_20048),
.B(n_9744),
.Y(n_20529)
);

AOI322xp5_ASAP7_75t_L g20530 ( 
.A1(n_20032),
.A2(n_9866),
.A3(n_10019),
.B1(n_11063),
.B2(n_11060),
.C1(n_10636),
.C2(n_10650),
.Y(n_20530)
);

AOI22xp5_ASAP7_75t_L g20531 ( 
.A1(n_20032),
.A2(n_9727),
.B1(n_9752),
.B2(n_9747),
.Y(n_20531)
);

NAND4xp25_ASAP7_75t_L g20532 ( 
.A(n_20100),
.B(n_8517),
.C(n_8460),
.D(n_8758),
.Y(n_20532)
);

INVxp67_ASAP7_75t_SL g20533 ( 
.A(n_20213),
.Y(n_20533)
);

INVx1_ASAP7_75t_L g20534 ( 
.A(n_20120),
.Y(n_20534)
);

INVx1_ASAP7_75t_L g20535 ( 
.A(n_20120),
.Y(n_20535)
);

OAI211xp5_ASAP7_75t_L g20536 ( 
.A1(n_20100),
.A2(n_9744),
.B(n_11069),
.C(n_9062),
.Y(n_20536)
);

AOI211xp5_ASAP7_75t_L g20537 ( 
.A1(n_20020),
.A2(n_9524),
.B(n_8714),
.C(n_8717),
.Y(n_20537)
);

AND2x2_ASAP7_75t_L g20538 ( 
.A(n_20120),
.B(n_9490),
.Y(n_20538)
);

NAND2xp5_ASAP7_75t_L g20539 ( 
.A(n_20015),
.B(n_9412),
.Y(n_20539)
);

A2O1A1O1Ixp25_ASAP7_75t_L g20540 ( 
.A1(n_20025),
.A2(n_9524),
.B(n_8779),
.C(n_11936),
.D(n_12161),
.Y(n_20540)
);

NAND2xp5_ASAP7_75t_L g20541 ( 
.A(n_20015),
.B(n_9310),
.Y(n_20541)
);

AOI22xp5_ASAP7_75t_L g20542 ( 
.A1(n_20032),
.A2(n_9727),
.B1(n_9752),
.B2(n_9747),
.Y(n_20542)
);

AOI22xp33_ASAP7_75t_L g20543 ( 
.A1(n_20120),
.A2(n_10991),
.B1(n_9981),
.B2(n_11209),
.Y(n_20543)
);

OAI221xp5_ASAP7_75t_L g20544 ( 
.A1(n_20100),
.A2(n_9377),
.B1(n_9333),
.B2(n_9841),
.C(n_9736),
.Y(n_20544)
);

INVx1_ASAP7_75t_L g20545 ( 
.A(n_20120),
.Y(n_20545)
);

O2A1O1Ixp5_ASAP7_75t_L g20546 ( 
.A1(n_20043),
.A2(n_10254),
.B(n_10266),
.C(n_10243),
.Y(n_20546)
);

OAI21xp5_ASAP7_75t_L g20547 ( 
.A1(n_20025),
.A2(n_11387),
.B(n_11381),
.Y(n_20547)
);

INVx2_ASAP7_75t_L g20548 ( 
.A(n_20103),
.Y(n_20548)
);

NOR2xp33_ASAP7_75t_L g20549 ( 
.A(n_20015),
.B(n_8612),
.Y(n_20549)
);

AOI22xp33_ASAP7_75t_L g20550 ( 
.A1(n_20120),
.A2(n_10991),
.B1(n_9981),
.B2(n_11209),
.Y(n_20550)
);

OAI211xp5_ASAP7_75t_L g20551 ( 
.A1(n_20100),
.A2(n_9744),
.B(n_9062),
.C(n_9727),
.Y(n_20551)
);

AOI221xp5_ASAP7_75t_L g20552 ( 
.A1(n_20020),
.A2(n_11063),
.B1(n_10636),
.B2(n_10650),
.C(n_10646),
.Y(n_20552)
);

AOI211xp5_ASAP7_75t_SL g20553 ( 
.A1(n_20055),
.A2(n_9747),
.B(n_9752),
.C(n_9727),
.Y(n_20553)
);

AOI322xp5_ASAP7_75t_L g20554 ( 
.A1(n_20032),
.A2(n_9866),
.A3(n_10019),
.B1(n_11063),
.B2(n_10634),
.C1(n_10717),
.C2(n_10660),
.Y(n_20554)
);

OAI22xp5_ASAP7_75t_L g20555 ( 
.A1(n_20055),
.A2(n_10976),
.B1(n_10660),
.B2(n_10717),
.Y(n_20555)
);

O2A1O1Ixp5_ASAP7_75t_SL g20556 ( 
.A1(n_20290),
.A2(n_9730),
.B(n_9748),
.C(n_9754),
.Y(n_20556)
);

XNOR2x1_ASAP7_75t_L g20557 ( 
.A(n_20428),
.B(n_9333),
.Y(n_20557)
);

OAI211xp5_ASAP7_75t_L g20558 ( 
.A1(n_20294),
.A2(n_9744),
.B(n_9748),
.C(n_9730),
.Y(n_20558)
);

AOI221xp5_ASAP7_75t_L g20559 ( 
.A1(n_20356),
.A2(n_10093),
.B1(n_10717),
.B2(n_10660),
.C(n_10646),
.Y(n_20559)
);

NOR2xp33_ASAP7_75t_L g20560 ( 
.A(n_20513),
.B(n_9736),
.Y(n_20560)
);

O2A1O1Ixp33_ASAP7_75t_L g20561 ( 
.A1(n_20527),
.A2(n_9742),
.B(n_9719),
.C(n_9558),
.Y(n_20561)
);

NAND3x1_ASAP7_75t_L g20562 ( 
.A(n_20369),
.B(n_11562),
.C(n_11564),
.Y(n_20562)
);

AOI22xp33_ASAP7_75t_L g20563 ( 
.A1(n_20534),
.A2(n_10991),
.B1(n_11232),
.B2(n_11209),
.Y(n_20563)
);

AOI22xp5_ASAP7_75t_L g20564 ( 
.A1(n_20535),
.A2(n_9747),
.B1(n_9752),
.B2(n_9727),
.Y(n_20564)
);

AOI221xp5_ASAP7_75t_L g20565 ( 
.A1(n_20335),
.A2(n_10646),
.B1(n_10848),
.B2(n_10843),
.C(n_10722),
.Y(n_20565)
);

OAI22xp5_ASAP7_75t_L g20566 ( 
.A1(n_20545),
.A2(n_20322),
.B1(n_20434),
.B2(n_20381),
.Y(n_20566)
);

NAND2xp5_ASAP7_75t_L g20567 ( 
.A(n_20538),
.B(n_9310),
.Y(n_20567)
);

NOR3xp33_ASAP7_75t_L g20568 ( 
.A(n_20417),
.B(n_8517),
.C(n_8460),
.Y(n_20568)
);

INVx2_ASAP7_75t_L g20569 ( 
.A(n_20289),
.Y(n_20569)
);

AOI221xp5_ASAP7_75t_L g20570 ( 
.A1(n_20338),
.A2(n_10722),
.B1(n_10861),
.B2(n_10848),
.C(n_10843),
.Y(n_20570)
);

A2O1A1Ixp33_ASAP7_75t_L g20571 ( 
.A1(n_20549),
.A2(n_10757),
.B(n_10663),
.C(n_10485),
.Y(n_20571)
);

NAND3xp33_ASAP7_75t_SL g20572 ( 
.A(n_20525),
.B(n_8653),
.C(n_8639),
.Y(n_20572)
);

AOI222xp33_ASAP7_75t_L g20573 ( 
.A1(n_20473),
.A2(n_20319),
.B1(n_20313),
.B2(n_20421),
.C1(n_20533),
.C2(n_20288),
.Y(n_20573)
);

AO22x1_ASAP7_75t_L g20574 ( 
.A1(n_20320),
.A2(n_10722),
.B1(n_10848),
.B2(n_10843),
.Y(n_20574)
);

NAND2xp5_ASAP7_75t_L g20575 ( 
.A(n_20548),
.B(n_9310),
.Y(n_20575)
);

INVx2_ASAP7_75t_L g20576 ( 
.A(n_20325),
.Y(n_20576)
);

NOR3xp33_ASAP7_75t_L g20577 ( 
.A(n_20393),
.B(n_8517),
.C(n_8460),
.Y(n_20577)
);

AO22x1_ASAP7_75t_L g20578 ( 
.A1(n_20418),
.A2(n_10861),
.B1(n_10883),
.B2(n_10881),
.Y(n_20578)
);

OAI221xp5_ASAP7_75t_L g20579 ( 
.A1(n_20308),
.A2(n_9997),
.B1(n_10091),
.B2(n_9841),
.C(n_9736),
.Y(n_20579)
);

AOI221xp5_ASAP7_75t_L g20580 ( 
.A1(n_20327),
.A2(n_10861),
.B1(n_10955),
.B2(n_10883),
.C(n_10881),
.Y(n_20580)
);

OAI21xp5_ASAP7_75t_SL g20581 ( 
.A1(n_20363),
.A2(n_9752),
.B(n_9727),
.Y(n_20581)
);

NOR3xp33_ASAP7_75t_L g20582 ( 
.A(n_20395),
.B(n_20409),
.C(n_20402),
.Y(n_20582)
);

NAND2xp5_ASAP7_75t_L g20583 ( 
.A(n_20301),
.B(n_9310),
.Y(n_20583)
);

AOI21xp33_ASAP7_75t_L g20584 ( 
.A1(n_20432),
.A2(n_9971),
.B(n_9981),
.Y(n_20584)
);

AOI221xp5_ASAP7_75t_L g20585 ( 
.A1(n_20359),
.A2(n_10881),
.B1(n_10961),
.B2(n_10955),
.C(n_10883),
.Y(n_20585)
);

O2A1O1Ixp33_ASAP7_75t_L g20586 ( 
.A1(n_20425),
.A2(n_9742),
.B(n_9719),
.C(n_9558),
.Y(n_20586)
);

NOR4xp25_ASAP7_75t_L g20587 ( 
.A(n_20375),
.B(n_8861),
.C(n_10961),
.D(n_10955),
.Y(n_20587)
);

AOI222xp33_ASAP7_75t_L g20588 ( 
.A1(n_20517),
.A2(n_10961),
.B1(n_10976),
.B2(n_9663),
.C1(n_9692),
.C2(n_10663),
.Y(n_20588)
);

AOI21xp5_ASAP7_75t_L g20589 ( 
.A1(n_20484),
.A2(n_10494),
.B(n_10485),
.Y(n_20589)
);

AOI22xp5_ASAP7_75t_L g20590 ( 
.A1(n_20323),
.A2(n_9752),
.B1(n_10976),
.B2(n_8653),
.Y(n_20590)
);

NAND2xp5_ASAP7_75t_L g20591 ( 
.A(n_20386),
.B(n_9310),
.Y(n_20591)
);

NAND4xp25_ASAP7_75t_L g20592 ( 
.A(n_20351),
.B(n_8517),
.C(n_8717),
.D(n_8714),
.Y(n_20592)
);

NAND2xp5_ASAP7_75t_L g20593 ( 
.A(n_20353),
.B(n_9310),
.Y(n_20593)
);

AOI221xp5_ASAP7_75t_L g20594 ( 
.A1(n_20291),
.A2(n_9692),
.B1(n_9663),
.B2(n_9247),
.C(n_9015),
.Y(n_20594)
);

AOI21xp33_ASAP7_75t_L g20595 ( 
.A1(n_20357),
.A2(n_9971),
.B(n_9981),
.Y(n_20595)
);

AOI322xp5_ASAP7_75t_L g20596 ( 
.A1(n_20442),
.A2(n_9692),
.A3(n_9663),
.B1(n_10003),
.B2(n_9945),
.C1(n_9857),
.C2(n_9821),
.Y(n_20596)
);

AOI22xp5_ASAP7_75t_L g20597 ( 
.A1(n_20544),
.A2(n_8639),
.B1(n_10303),
.B2(n_11279),
.Y(n_20597)
);

A2O1A1Ixp33_ASAP7_75t_L g20598 ( 
.A1(n_20528),
.A2(n_20458),
.B(n_20489),
.C(n_20328),
.Y(n_20598)
);

AOI22xp5_ASAP7_75t_L g20599 ( 
.A1(n_20532),
.A2(n_10303),
.B1(n_11282),
.B2(n_11279),
.Y(n_20599)
);

OAI22xp33_ASAP7_75t_L g20600 ( 
.A1(n_20343),
.A2(n_9744),
.B1(n_10032),
.B2(n_9869),
.Y(n_20600)
);

OAI21xp5_ASAP7_75t_L g20601 ( 
.A1(n_20292),
.A2(n_11387),
.B(n_10287),
.Y(n_20601)
);

AOI21xp33_ASAP7_75t_SL g20602 ( 
.A1(n_20362),
.A2(n_9971),
.B(n_10303),
.Y(n_20602)
);

NAND2xp5_ASAP7_75t_L g20603 ( 
.A(n_20366),
.B(n_20367),
.Y(n_20603)
);

A2O1A1Ixp33_ASAP7_75t_L g20604 ( 
.A1(n_20352),
.A2(n_10757),
.B(n_10485),
.C(n_10494),
.Y(n_20604)
);

OAI211xp5_ASAP7_75t_L g20605 ( 
.A1(n_20315),
.A2(n_20374),
.B(n_20408),
.C(n_20472),
.Y(n_20605)
);

NOR3xp33_ASAP7_75t_L g20606 ( 
.A(n_20445),
.B(n_8517),
.C(n_10243),
.Y(n_20606)
);

NAND3xp33_ASAP7_75t_L g20607 ( 
.A(n_20511),
.B(n_9744),
.C(n_9869),
.Y(n_20607)
);

NOR4xp25_ASAP7_75t_L g20608 ( 
.A(n_20342),
.B(n_8861),
.C(n_8703),
.D(n_9710),
.Y(n_20608)
);

NAND4xp25_ASAP7_75t_SL g20609 ( 
.A(n_20551),
.B(n_8703),
.C(n_8717),
.D(n_8714),
.Y(n_20609)
);

OAI221xp5_ASAP7_75t_L g20610 ( 
.A1(n_20314),
.A2(n_9736),
.B1(n_10091),
.B2(n_9997),
.C(n_9841),
.Y(n_20610)
);

AOI22xp33_ASAP7_75t_L g20611 ( 
.A1(n_20437),
.A2(n_11232),
.B1(n_11209),
.B2(n_9981),
.Y(n_20611)
);

O2A1O1Ixp33_ASAP7_75t_L g20612 ( 
.A1(n_20400),
.A2(n_20483),
.B(n_20495),
.C(n_20449),
.Y(n_20612)
);

AOI221xp5_ASAP7_75t_L g20613 ( 
.A1(n_20485),
.A2(n_9692),
.B1(n_9663),
.B2(n_9247),
.C(n_9015),
.Y(n_20613)
);

NAND2xp5_ASAP7_75t_SL g20614 ( 
.A(n_20365),
.B(n_9744),
.Y(n_20614)
);

NAND2xp5_ASAP7_75t_L g20615 ( 
.A(n_20348),
.B(n_9310),
.Y(n_20615)
);

INVx1_ASAP7_75t_L g20616 ( 
.A(n_20341),
.Y(n_20616)
);

OR2x2_ASAP7_75t_L g20617 ( 
.A(n_20383),
.B(n_10546),
.Y(n_20617)
);

AO22x1_ASAP7_75t_L g20618 ( 
.A1(n_20337),
.A2(n_9663),
.B1(n_9692),
.B2(n_9710),
.Y(n_20618)
);

OAI21xp33_ASAP7_75t_L g20619 ( 
.A1(n_20524),
.A2(n_9718),
.B(n_9710),
.Y(n_20619)
);

AOI21xp5_ASAP7_75t_L g20620 ( 
.A1(n_20480),
.A2(n_10494),
.B(n_10483),
.Y(n_20620)
);

AOI32xp33_ASAP7_75t_L g20621 ( 
.A1(n_20459),
.A2(n_9066),
.A3(n_9543),
.B1(n_9553),
.B2(n_9490),
.Y(n_20621)
);

AOI221xp5_ASAP7_75t_L g20622 ( 
.A1(n_20355),
.A2(n_9692),
.B1(n_9663),
.B2(n_9247),
.C(n_9015),
.Y(n_20622)
);

OAI32xp33_ASAP7_75t_L g20623 ( 
.A1(n_20333),
.A2(n_9722),
.A3(n_9718),
.B1(n_9710),
.B2(n_9805),
.Y(n_20623)
);

NAND2xp5_ASAP7_75t_SL g20624 ( 
.A(n_20379),
.B(n_9869),
.Y(n_20624)
);

OAI21xp5_ASAP7_75t_SL g20625 ( 
.A1(n_20465),
.A2(n_9066),
.B(n_9490),
.Y(n_20625)
);

OAI221xp5_ASAP7_75t_L g20626 ( 
.A1(n_20450),
.A2(n_9736),
.B1(n_10091),
.B2(n_9997),
.C(n_9841),
.Y(n_20626)
);

NOR2xp33_ASAP7_75t_L g20627 ( 
.A(n_20516),
.B(n_9736),
.Y(n_20627)
);

AOI22xp5_ASAP7_75t_L g20628 ( 
.A1(n_20479),
.A2(n_11282),
.B1(n_11279),
.B2(n_11296),
.Y(n_20628)
);

OAI21xp33_ASAP7_75t_SL g20629 ( 
.A1(n_20326),
.A2(n_10469),
.B(n_10462),
.Y(n_20629)
);

NAND4xp25_ASAP7_75t_L g20630 ( 
.A(n_20487),
.B(n_9066),
.C(n_8521),
.D(n_8939),
.Y(n_20630)
);

OAI21xp33_ASAP7_75t_L g20631 ( 
.A1(n_20422),
.A2(n_9718),
.B(n_9710),
.Y(n_20631)
);

AND2x2_ASAP7_75t_L g20632 ( 
.A(n_20497),
.B(n_9490),
.Y(n_20632)
);

NOR3xp33_ASAP7_75t_L g20633 ( 
.A(n_20467),
.B(n_10254),
.C(n_10243),
.Y(n_20633)
);

OAI221xp5_ASAP7_75t_L g20634 ( 
.A1(n_20455),
.A2(n_9736),
.B1(n_10091),
.B2(n_9997),
.C(n_9841),
.Y(n_20634)
);

OAI22xp5_ASAP7_75t_L g20635 ( 
.A1(n_20298),
.A2(n_9710),
.B1(n_9722),
.B2(n_9718),
.Y(n_20635)
);

NOR2xp33_ASAP7_75t_L g20636 ( 
.A(n_20471),
.B(n_9736),
.Y(n_20636)
);

OAI211xp5_ASAP7_75t_SL g20637 ( 
.A1(n_20482),
.A2(n_8521),
.B(n_9543),
.C(n_9490),
.Y(n_20637)
);

OAI221xp5_ASAP7_75t_L g20638 ( 
.A1(n_20515),
.A2(n_9841),
.B1(n_10100),
.B2(n_10091),
.C(n_9997),
.Y(n_20638)
);

NOR2xp33_ASAP7_75t_L g20639 ( 
.A(n_20468),
.B(n_9841),
.Y(n_20639)
);

AOI22xp5_ASAP7_75t_L g20640 ( 
.A1(n_20502),
.A2(n_11279),
.B1(n_11282),
.B2(n_11296),
.Y(n_20640)
);

AO221x1_ASAP7_75t_L g20641 ( 
.A1(n_20481),
.A2(n_9015),
.B1(n_9505),
.B2(n_9517),
.C(n_9504),
.Y(n_20641)
);

AOI22xp5_ASAP7_75t_L g20642 ( 
.A1(n_20536),
.A2(n_20509),
.B1(n_20441),
.B2(n_20336),
.Y(n_20642)
);

NAND5xp2_ASAP7_75t_L g20643 ( 
.A(n_20453),
.B(n_9027),
.C(n_9289),
.D(n_9300),
.E(n_9293),
.Y(n_20643)
);

OAI21xp5_ASAP7_75t_SL g20644 ( 
.A1(n_20361),
.A2(n_9066),
.B(n_9490),
.Y(n_20644)
);

INVx1_ASAP7_75t_L g20645 ( 
.A(n_20463),
.Y(n_20645)
);

INVx1_ASAP7_75t_L g20646 ( 
.A(n_20474),
.Y(n_20646)
);

AND2x4_ASAP7_75t_L g20647 ( 
.A(n_20529),
.B(n_9543),
.Y(n_20647)
);

A2O1A1Ixp33_ASAP7_75t_L g20648 ( 
.A1(n_20398),
.A2(n_10495),
.B(n_10496),
.C(n_10483),
.Y(n_20648)
);

OAI221xp5_ASAP7_75t_L g20649 ( 
.A1(n_20410),
.A2(n_9841),
.B1(n_10100),
.B2(n_10091),
.C(n_9997),
.Y(n_20649)
);

NOR2x1_ASAP7_75t_L g20650 ( 
.A(n_20460),
.B(n_9763),
.Y(n_20650)
);

NAND3xp33_ASAP7_75t_SL g20651 ( 
.A(n_20461),
.B(n_9289),
.C(n_9027),
.Y(n_20651)
);

AOI221xp5_ASAP7_75t_L g20652 ( 
.A1(n_20539),
.A2(n_9247),
.B1(n_9722),
.B2(n_9718),
.C(n_9304),
.Y(n_20652)
);

NOR2xp33_ASAP7_75t_L g20653 ( 
.A(n_20312),
.B(n_9997),
.Y(n_20653)
);

NOR2xp33_ASAP7_75t_L g20654 ( 
.A(n_20541),
.B(n_9997),
.Y(n_20654)
);

INVx1_ASAP7_75t_L g20655 ( 
.A(n_20388),
.Y(n_20655)
);

OAI22xp5_ASAP7_75t_L g20656 ( 
.A1(n_20296),
.A2(n_9718),
.B1(n_9722),
.B2(n_9754),
.Y(n_20656)
);

AND2x2_ASAP7_75t_L g20657 ( 
.A(n_20537),
.B(n_9543),
.Y(n_20657)
);

NAND2xp5_ASAP7_75t_SL g20658 ( 
.A(n_20514),
.B(n_9869),
.Y(n_20658)
);

OR2x2_ASAP7_75t_L g20659 ( 
.A(n_20526),
.B(n_10546),
.Y(n_20659)
);

AOI221xp5_ASAP7_75t_L g20660 ( 
.A1(n_20406),
.A2(n_9722),
.B1(n_9304),
.B2(n_9742),
.C(n_9504),
.Y(n_20660)
);

NOR4xp25_ASAP7_75t_L g20661 ( 
.A(n_20391),
.B(n_9722),
.C(n_9754),
.D(n_8662),
.Y(n_20661)
);

AO21x1_ASAP7_75t_L g20662 ( 
.A1(n_20439),
.A2(n_10266),
.B(n_10462),
.Y(n_20662)
);

AOI211xp5_ASAP7_75t_L g20663 ( 
.A1(n_20387),
.A2(n_10839),
.B(n_11248),
.C(n_11245),
.Y(n_20663)
);

NAND4xp25_ASAP7_75t_L g20664 ( 
.A(n_20302),
.B(n_9066),
.C(n_8939),
.D(n_8734),
.Y(n_20664)
);

NOR3xp33_ASAP7_75t_L g20665 ( 
.A(n_20380),
.B(n_10882),
.C(n_10875),
.Y(n_20665)
);

AOI322xp5_ASAP7_75t_L g20666 ( 
.A1(n_20426),
.A2(n_9875),
.A3(n_9857),
.B1(n_9867),
.B2(n_9885),
.C1(n_9821),
.C2(n_9805),
.Y(n_20666)
);

A2O1A1Ixp33_ASAP7_75t_L g20667 ( 
.A1(n_20478),
.A2(n_20523),
.B(n_20518),
.C(n_20321),
.Y(n_20667)
);

NAND4xp25_ASAP7_75t_L g20668 ( 
.A(n_20469),
.B(n_9066),
.C(n_8734),
.D(n_8815),
.Y(n_20668)
);

A2O1A1Ixp33_ASAP7_75t_L g20669 ( 
.A1(n_20293),
.A2(n_10495),
.B(n_10496),
.C(n_10483),
.Y(n_20669)
);

AOI221xp5_ASAP7_75t_L g20670 ( 
.A1(n_20491),
.A2(n_9304),
.B1(n_9742),
.B2(n_9504),
.C(n_9517),
.Y(n_20670)
);

NOR4xp75_ASAP7_75t_SL g20671 ( 
.A(n_20475),
.B(n_9212),
.C(n_9058),
.D(n_8912),
.Y(n_20671)
);

OAI21xp33_ASAP7_75t_L g20672 ( 
.A1(n_20407),
.A2(n_20299),
.B(n_20373),
.Y(n_20672)
);

AOI21xp5_ASAP7_75t_L g20673 ( 
.A1(n_20424),
.A2(n_10496),
.B(n_10495),
.Y(n_20673)
);

AOI21xp33_ASAP7_75t_SL g20674 ( 
.A1(n_20448),
.A2(n_9971),
.B(n_9981),
.Y(n_20674)
);

OAI21xp5_ASAP7_75t_L g20675 ( 
.A1(n_20493),
.A2(n_20547),
.B(n_20540),
.Y(n_20675)
);

AOI22x1_ASAP7_75t_L g20676 ( 
.A1(n_20522),
.A2(n_9558),
.B1(n_9584),
.B2(n_9533),
.Y(n_20676)
);

O2A1O1Ixp33_ASAP7_75t_L g20677 ( 
.A1(n_20405),
.A2(n_9558),
.B(n_9584),
.C(n_9533),
.Y(n_20677)
);

AND2x2_ASAP7_75t_L g20678 ( 
.A(n_20310),
.B(n_9543),
.Y(n_20678)
);

OAI21xp33_ASAP7_75t_L g20679 ( 
.A1(n_20399),
.A2(n_9553),
.B(n_9543),
.Y(n_20679)
);

AOI21xp5_ASAP7_75t_L g20680 ( 
.A1(n_20457),
.A2(n_11232),
.B(n_10421),
.Y(n_20680)
);

NOR3xp33_ASAP7_75t_SL g20681 ( 
.A(n_20504),
.B(n_9062),
.C(n_8592),
.Y(n_20681)
);

AOI21xp5_ASAP7_75t_L g20682 ( 
.A1(n_20390),
.A2(n_11232),
.B(n_10421),
.Y(n_20682)
);

NOR3xp33_ASAP7_75t_L g20683 ( 
.A(n_20520),
.B(n_10882),
.C(n_10875),
.Y(n_20683)
);

OAI221xp5_ASAP7_75t_L g20684 ( 
.A1(n_20499),
.A2(n_9997),
.B1(n_10100),
.B2(n_10091),
.C(n_9377),
.Y(n_20684)
);

OAI21xp33_ASAP7_75t_L g20685 ( 
.A1(n_20345),
.A2(n_9553),
.B(n_9543),
.Y(n_20685)
);

AOI21xp5_ASAP7_75t_L g20686 ( 
.A1(n_20494),
.A2(n_11232),
.B(n_10421),
.Y(n_20686)
);

AOI211xp5_ASAP7_75t_L g20687 ( 
.A1(n_20376),
.A2(n_10839),
.B(n_11248),
.C(n_11245),
.Y(n_20687)
);

AOI22xp5_ASAP7_75t_L g20688 ( 
.A1(n_20501),
.A2(n_11282),
.B1(n_11279),
.B2(n_11296),
.Y(n_20688)
);

NAND2xp5_ASAP7_75t_SL g20689 ( 
.A(n_20438),
.B(n_9869),
.Y(n_20689)
);

OAI211xp5_ASAP7_75t_SL g20690 ( 
.A1(n_20372),
.A2(n_9553),
.B(n_9543),
.C(n_8822),
.Y(n_20690)
);

OAI21xp5_ASAP7_75t_L g20691 ( 
.A1(n_20370),
.A2(n_11387),
.B(n_10287),
.Y(n_20691)
);

AOI21xp5_ASAP7_75t_L g20692 ( 
.A1(n_20466),
.A2(n_11232),
.B(n_10425),
.Y(n_20692)
);

O2A1O1Ixp33_ASAP7_75t_L g20693 ( 
.A1(n_20508),
.A2(n_9584),
.B(n_9533),
.C(n_9505),
.Y(n_20693)
);

A2O1A1Ixp33_ASAP7_75t_L g20694 ( 
.A1(n_20553),
.A2(n_10621),
.B(n_10603),
.C(n_10624),
.Y(n_20694)
);

OAI22xp5_ASAP7_75t_L g20695 ( 
.A1(n_20531),
.A2(n_9805),
.B1(n_9857),
.B2(n_9821),
.Y(n_20695)
);

OAI21xp5_ASAP7_75t_SL g20696 ( 
.A1(n_20542),
.A2(n_9553),
.B(n_9289),
.Y(n_20696)
);

AOI211xp5_ASAP7_75t_L g20697 ( 
.A1(n_20300),
.A2(n_10839),
.B(n_11248),
.C(n_11245),
.Y(n_20697)
);

INVx1_ASAP7_75t_L g20698 ( 
.A(n_20477),
.Y(n_20698)
);

AOI322xp5_ASAP7_75t_L g20699 ( 
.A1(n_20470),
.A2(n_9938),
.A3(n_10003),
.B1(n_9931),
.B2(n_9875),
.C1(n_9940),
.C2(n_9885),
.Y(n_20699)
);

OAI22xp5_ASAP7_75t_L g20700 ( 
.A1(n_20476),
.A2(n_9867),
.B1(n_9885),
.B2(n_9875),
.Y(n_20700)
);

OAI211xp5_ASAP7_75t_L g20701 ( 
.A1(n_20297),
.A2(n_20443),
.B(n_20307),
.C(n_20488),
.Y(n_20701)
);

OAI21xp5_ASAP7_75t_SL g20702 ( 
.A1(n_20364),
.A2(n_9553),
.B(n_9289),
.Y(n_20702)
);

OAI221xp5_ASAP7_75t_L g20703 ( 
.A1(n_20382),
.A2(n_9997),
.B1(n_10100),
.B2(n_10091),
.C(n_9377),
.Y(n_20703)
);

NOR2xp67_ASAP7_75t_L g20704 ( 
.A(n_20492),
.B(n_10051),
.Y(n_20704)
);

AND2x2_ASAP7_75t_L g20705 ( 
.A(n_20329),
.B(n_20331),
.Y(n_20705)
);

NAND2xp5_ASAP7_75t_L g20706 ( 
.A(n_20303),
.B(n_9310),
.Y(n_20706)
);

A2O1A1Ixp33_ASAP7_75t_L g20707 ( 
.A1(n_20371),
.A2(n_10621),
.B(n_10603),
.C(n_10624),
.Y(n_20707)
);

NAND2xp5_ASAP7_75t_L g20708 ( 
.A(n_20505),
.B(n_9314),
.Y(n_20708)
);

INVx1_ASAP7_75t_L g20709 ( 
.A(n_20506),
.Y(n_20709)
);

OAI21xp33_ASAP7_75t_SL g20710 ( 
.A1(n_20436),
.A2(n_10469),
.B(n_10462),
.Y(n_20710)
);

AOI22xp5_ASAP7_75t_L g20711 ( 
.A1(n_20344),
.A2(n_11279),
.B1(n_11282),
.B2(n_11296),
.Y(n_20711)
);

NAND4xp25_ASAP7_75t_SL g20712 ( 
.A(n_20415),
.B(n_8662),
.C(n_9033),
.D(n_9020),
.Y(n_20712)
);

OAI21xp33_ASAP7_75t_L g20713 ( 
.A1(n_20431),
.A2(n_9553),
.B(n_11564),
.Y(n_20713)
);

AOI221xp5_ASAP7_75t_L g20714 ( 
.A1(n_20394),
.A2(n_9304),
.B1(n_9504),
.B2(n_9517),
.C(n_9505),
.Y(n_20714)
);

AOI221xp5_ASAP7_75t_L g20715 ( 
.A1(n_20403),
.A2(n_9517),
.B1(n_9505),
.B2(n_9584),
.C(n_9533),
.Y(n_20715)
);

AOI221x1_ASAP7_75t_L g20716 ( 
.A1(n_20318),
.A2(n_9988),
.B1(n_9992),
.B2(n_9980),
.C(n_9979),
.Y(n_20716)
);

AOI322xp5_ASAP7_75t_L g20717 ( 
.A1(n_20304),
.A2(n_9867),
.A3(n_9940),
.B1(n_9945),
.B2(n_10003),
.C1(n_9938),
.C2(n_9931),
.Y(n_20717)
);

OAI22xp5_ASAP7_75t_L g20718 ( 
.A1(n_20456),
.A2(n_9931),
.B1(n_9940),
.B2(n_9938),
.Y(n_20718)
);

AOI22xp33_ASAP7_75t_L g20719 ( 
.A1(n_20464),
.A2(n_11282),
.B1(n_10206),
.B2(n_10225),
.Y(n_20719)
);

NAND2xp5_ASAP7_75t_L g20720 ( 
.A(n_20464),
.B(n_9314),
.Y(n_20720)
);

OAI211xp5_ASAP7_75t_SL g20721 ( 
.A1(n_20447),
.A2(n_9553),
.B(n_8822),
.C(n_9502),
.Y(n_20721)
);

INVx1_ASAP7_75t_L g20722 ( 
.A(n_20496),
.Y(n_20722)
);

NOR2xp33_ASAP7_75t_L g20723 ( 
.A(n_20433),
.B(n_10091),
.Y(n_20723)
);

AOI311xp33_ASAP7_75t_L g20724 ( 
.A1(n_20411),
.A2(n_9039),
.A3(n_9041),
.B(n_9033),
.C(n_9023),
.Y(n_20724)
);

O2A1O1Ixp33_ASAP7_75t_L g20725 ( 
.A1(n_20350),
.A2(n_20349),
.B(n_20452),
.C(n_20309),
.Y(n_20725)
);

NOR2xp33_ASAP7_75t_SL g20726 ( 
.A(n_20412),
.B(n_9869),
.Y(n_20726)
);

AOI21xp5_ASAP7_75t_L g20727 ( 
.A1(n_20311),
.A2(n_10425),
.B(n_10412),
.Y(n_20727)
);

OAI221xp5_ASAP7_75t_L g20728 ( 
.A1(n_20430),
.A2(n_10091),
.B1(n_10100),
.B2(n_9377),
.C(n_9333),
.Y(n_20728)
);

NOR2xp33_ASAP7_75t_L g20729 ( 
.A(n_20358),
.B(n_10100),
.Y(n_20729)
);

INVx1_ASAP7_75t_SL g20730 ( 
.A(n_20454),
.Y(n_20730)
);

NOR2xp33_ASAP7_75t_L g20731 ( 
.A(n_20316),
.B(n_10100),
.Y(n_20731)
);

OAI33xp33_ASAP7_75t_L g20732 ( 
.A1(n_20519),
.A2(n_9041),
.A3(n_9033),
.B1(n_9045),
.B2(n_9039),
.B3(n_9023),
.Y(n_20732)
);

AOI21xp5_ASAP7_75t_L g20733 ( 
.A1(n_20330),
.A2(n_10425),
.B(n_10412),
.Y(n_20733)
);

AOI221xp5_ASAP7_75t_L g20734 ( 
.A1(n_20555),
.A2(n_9802),
.B1(n_8342),
.B2(n_8448),
.C(n_8277),
.Y(n_20734)
);

NAND4xp25_ASAP7_75t_L g20735 ( 
.A(n_20378),
.B(n_20500),
.C(n_20385),
.D(n_20305),
.Y(n_20735)
);

AOI22xp5_ASAP7_75t_L g20736 ( 
.A1(n_20444),
.A2(n_11300),
.B1(n_11296),
.B2(n_10927),
.Y(n_20736)
);

NAND2xp5_ASAP7_75t_SL g20737 ( 
.A(n_20384),
.B(n_20397),
.Y(n_20737)
);

AOI221xp5_ASAP7_75t_L g20738 ( 
.A1(n_20423),
.A2(n_9802),
.B1(n_8342),
.B2(n_8448),
.C(n_8277),
.Y(n_20738)
);

NAND2xp5_ASAP7_75t_L g20739 ( 
.A(n_20440),
.B(n_9314),
.Y(n_20739)
);

NOR2xp33_ASAP7_75t_L g20740 ( 
.A(n_20420),
.B(n_10100),
.Y(n_20740)
);

OAI221xp5_ASAP7_75t_L g20741 ( 
.A1(n_20377),
.A2(n_10100),
.B1(n_8988),
.B2(n_9289),
.C(n_9027),
.Y(n_20741)
);

AOI221xp5_ASAP7_75t_L g20742 ( 
.A1(n_20503),
.A2(n_9802),
.B1(n_8618),
.B2(n_8453),
.C(n_8015),
.Y(n_20742)
);

NAND4xp25_ASAP7_75t_SL g20743 ( 
.A(n_20552),
.B(n_9033),
.C(n_9039),
.D(n_9023),
.Y(n_20743)
);

INVx1_ASAP7_75t_L g20744 ( 
.A(n_20546),
.Y(n_20744)
);

NAND2xp5_ASAP7_75t_L g20745 ( 
.A(n_20486),
.B(n_9314),
.Y(n_20745)
);

AOI21xp5_ASAP7_75t_L g20746 ( 
.A1(n_20462),
.A2(n_10426),
.B(n_10412),
.Y(n_20746)
);

AND3x1_ASAP7_75t_L g20747 ( 
.A(n_20427),
.B(n_9212),
.C(n_9302),
.Y(n_20747)
);

NAND2xp5_ASAP7_75t_L g20748 ( 
.A(n_20507),
.B(n_9314),
.Y(n_20748)
);

OAI22xp5_ASAP7_75t_L g20749 ( 
.A1(n_20543),
.A2(n_10130),
.B1(n_9945),
.B2(n_10051),
.Y(n_20749)
);

NOR3xp33_ASAP7_75t_L g20750 ( 
.A(n_20413),
.B(n_10882),
.C(n_10875),
.Y(n_20750)
);

AOI21xp5_ASAP7_75t_L g20751 ( 
.A1(n_20346),
.A2(n_10428),
.B(n_10426),
.Y(n_20751)
);

NAND2xp5_ASAP7_75t_L g20752 ( 
.A(n_20295),
.B(n_20306),
.Y(n_20752)
);

NAND2xp5_ASAP7_75t_L g20753 ( 
.A(n_20435),
.B(n_20510),
.Y(n_20753)
);

AOI22xp5_ASAP7_75t_L g20754 ( 
.A1(n_20334),
.A2(n_11300),
.B1(n_11296),
.B2(n_10927),
.Y(n_20754)
);

OR2x2_ASAP7_75t_L g20755 ( 
.A(n_20360),
.B(n_10546),
.Y(n_20755)
);

NOR2xp33_ASAP7_75t_L g20756 ( 
.A(n_20498),
.B(n_10100),
.Y(n_20756)
);

AOI21xp33_ASAP7_75t_L g20757 ( 
.A1(n_20339),
.A2(n_11300),
.B(n_10989),
.Y(n_20757)
);

NOR3xp33_ASAP7_75t_L g20758 ( 
.A(n_20512),
.B(n_20416),
.C(n_20521),
.Y(n_20758)
);

NAND4xp25_ASAP7_75t_SL g20759 ( 
.A(n_20317),
.B(n_9039),
.C(n_9041),
.D(n_9023),
.Y(n_20759)
);

OAI21xp5_ASAP7_75t_L g20760 ( 
.A1(n_20490),
.A2(n_20324),
.B(n_20550),
.Y(n_20760)
);

NOR2xp33_ASAP7_75t_L g20761 ( 
.A(n_20451),
.B(n_10032),
.Y(n_20761)
);

NOR2xp33_ASAP7_75t_L g20762 ( 
.A(n_20404),
.B(n_20429),
.Y(n_20762)
);

NAND2xp5_ASAP7_75t_L g20763 ( 
.A(n_20396),
.B(n_9314),
.Y(n_20763)
);

OAI21xp5_ASAP7_75t_L g20764 ( 
.A1(n_20347),
.A2(n_10287),
.B(n_11570),
.Y(n_20764)
);

AOI21xp5_ASAP7_75t_L g20765 ( 
.A1(n_20340),
.A2(n_10433),
.B(n_10428),
.Y(n_20765)
);

OAI21xp5_ASAP7_75t_L g20766 ( 
.A1(n_20389),
.A2(n_11570),
.B(n_10629),
.Y(n_20766)
);

OAI211xp5_ASAP7_75t_L g20767 ( 
.A1(n_20392),
.A2(n_11477),
.B(n_11087),
.C(n_10051),
.Y(n_20767)
);

INVx1_ASAP7_75t_L g20768 ( 
.A(n_20332),
.Y(n_20768)
);

INVx1_ASAP7_75t_L g20769 ( 
.A(n_20368),
.Y(n_20769)
);

AOI21xp5_ASAP7_75t_L g20770 ( 
.A1(n_20401),
.A2(n_20354),
.B(n_20419),
.Y(n_20770)
);

INVx2_ASAP7_75t_L g20771 ( 
.A(n_20414),
.Y(n_20771)
);

OAI211xp5_ASAP7_75t_L g20772 ( 
.A1(n_20530),
.A2(n_11477),
.B(n_11087),
.C(n_10051),
.Y(n_20772)
);

NOR3xp33_ASAP7_75t_L g20773 ( 
.A(n_20554),
.B(n_10912),
.C(n_10900),
.Y(n_20773)
);

OAI221xp5_ASAP7_75t_L g20774 ( 
.A1(n_20446),
.A2(n_8988),
.B1(n_9289),
.B2(n_9027),
.C(n_10032),
.Y(n_20774)
);

NAND2xp5_ASAP7_75t_L g20775 ( 
.A(n_20538),
.B(n_9314),
.Y(n_20775)
);

INVx1_ASAP7_75t_L g20776 ( 
.A(n_20538),
.Y(n_20776)
);

NOR4xp25_ASAP7_75t_SL g20777 ( 
.A(n_20525),
.B(n_8962),
.C(n_7779),
.D(n_7918),
.Y(n_20777)
);

NOR2xp33_ASAP7_75t_SL g20778 ( 
.A(n_20289),
.B(n_10032),
.Y(n_20778)
);

AOI22xp5_ASAP7_75t_L g20779 ( 
.A1(n_20290),
.A2(n_11300),
.B1(n_10927),
.B2(n_10917),
.Y(n_20779)
);

NOR3xp33_ASAP7_75t_L g20780 ( 
.A(n_20294),
.B(n_10912),
.C(n_10900),
.Y(n_20780)
);

INVx2_ASAP7_75t_L g20781 ( 
.A(n_20289),
.Y(n_20781)
);

AOI221xp5_ASAP7_75t_L g20782 ( 
.A1(n_20356),
.A2(n_9802),
.B1(n_8618),
.B2(n_8453),
.C(n_8015),
.Y(n_20782)
);

INVx2_ASAP7_75t_L g20783 ( 
.A(n_20289),
.Y(n_20783)
);

AOI222xp33_ASAP7_75t_L g20784 ( 
.A1(n_20572),
.A2(n_10469),
.B1(n_10479),
.B2(n_10603),
.C1(n_10629),
.C2(n_10624),
.Y(n_20784)
);

OAI32xp33_ASAP7_75t_L g20785 ( 
.A1(n_20780),
.A2(n_10130),
.A3(n_9043),
.B1(n_9071),
.B2(n_9052),
.Y(n_20785)
);

NOR2xp33_ASAP7_75t_L g20786 ( 
.A(n_20569),
.B(n_10032),
.Y(n_20786)
);

AOI21xp5_ASAP7_75t_L g20787 ( 
.A1(n_20612),
.A2(n_10479),
.B(n_10433),
.Y(n_20787)
);

NOR2xp33_ASAP7_75t_L g20788 ( 
.A(n_20781),
.B(n_10032),
.Y(n_20788)
);

OAI32xp33_ASAP7_75t_L g20789 ( 
.A1(n_20582),
.A2(n_10130),
.A3(n_9043),
.B1(n_9071),
.B2(n_9052),
.Y(n_20789)
);

OAI211xp5_ASAP7_75t_SL g20790 ( 
.A1(n_20573),
.A2(n_9502),
.B(n_9980),
.C(n_9979),
.Y(n_20790)
);

OAI211xp5_ASAP7_75t_L g20791 ( 
.A1(n_20605),
.A2(n_11087),
.B(n_10927),
.C(n_10917),
.Y(n_20791)
);

NOR3xp33_ASAP7_75t_L g20792 ( 
.A(n_20603),
.B(n_10912),
.C(n_10900),
.Y(n_20792)
);

NAND2xp5_ASAP7_75t_L g20793 ( 
.A(n_20560),
.B(n_9314),
.Y(n_20793)
);

AOI221xp5_ASAP7_75t_L g20794 ( 
.A1(n_20566),
.A2(n_10006),
.B1(n_9828),
.B2(n_9763),
.C(n_9571),
.Y(n_20794)
);

NOR3xp33_ASAP7_75t_L g20795 ( 
.A(n_20783),
.B(n_10822),
.C(n_11406),
.Y(n_20795)
);

AOI21xp5_ASAP7_75t_L g20796 ( 
.A1(n_20737),
.A2(n_10479),
.B(n_10428),
.Y(n_20796)
);

O2A1O1Ixp33_ASAP7_75t_L g20797 ( 
.A1(n_20576),
.A2(n_9645),
.B(n_8988),
.C(n_9642),
.Y(n_20797)
);

AND2x2_ASAP7_75t_L g20798 ( 
.A(n_20771),
.B(n_8597),
.Y(n_20798)
);

O2A1O1Ixp33_ASAP7_75t_L g20799 ( 
.A1(n_20598),
.A2(n_9645),
.B(n_8988),
.C(n_9642),
.Y(n_20799)
);

OA22x2_ASAP7_75t_L g20800 ( 
.A1(n_20625),
.A2(n_10946),
.B1(n_10951),
.B2(n_10964),
.Y(n_20800)
);

OAI31xp33_ASAP7_75t_L g20801 ( 
.A1(n_20558),
.A2(n_9027),
.A3(n_9300),
.B(n_9293),
.Y(n_20801)
);

AOI21xp5_ASAP7_75t_L g20802 ( 
.A1(n_20752),
.A2(n_10433),
.B(n_10426),
.Y(n_20802)
);

AOI221xp5_ASAP7_75t_L g20803 ( 
.A1(n_20762),
.A2(n_10006),
.B1(n_9828),
.B2(n_9571),
.C(n_9651),
.Y(n_20803)
);

OAI221xp5_ASAP7_75t_L g20804 ( 
.A1(n_20675),
.A2(n_8988),
.B1(n_9027),
.B2(n_9300),
.C(n_9293),
.Y(n_20804)
);

O2A1O1Ixp33_ASAP7_75t_L g20805 ( 
.A1(n_20616),
.A2(n_9645),
.B(n_8988),
.C(n_9642),
.Y(n_20805)
);

O2A1O1Ixp33_ASAP7_75t_L g20806 ( 
.A1(n_20646),
.A2(n_9645),
.B(n_8988),
.C(n_9642),
.Y(n_20806)
);

OAI21xp33_ASAP7_75t_SL g20807 ( 
.A1(n_20768),
.A2(n_10398),
.B(n_10397),
.Y(n_20807)
);

OAI221xp5_ASAP7_75t_L g20808 ( 
.A1(n_20672),
.A2(n_8988),
.B1(n_9300),
.B2(n_9339),
.C(n_9293),
.Y(n_20808)
);

OAI222xp33_ASAP7_75t_L g20809 ( 
.A1(n_20650),
.A2(n_11506),
.B1(n_11504),
.B2(n_9358),
.C1(n_9300),
.C2(n_9378),
.Y(n_20809)
);

AOI221xp5_ASAP7_75t_L g20810 ( 
.A1(n_20725),
.A2(n_20636),
.B1(n_20579),
.B2(n_20639),
.C(n_20587),
.Y(n_20810)
);

NAND2xp5_ASAP7_75t_L g20811 ( 
.A(n_20731),
.B(n_10546),
.Y(n_20811)
);

AOI22xp5_ASAP7_75t_L g20812 ( 
.A1(n_20756),
.A2(n_10927),
.B1(n_10917),
.B2(n_11300),
.Y(n_20812)
);

OAI211xp5_ASAP7_75t_L g20813 ( 
.A1(n_20769),
.A2(n_10927),
.B(n_10917),
.C(n_10051),
.Y(n_20813)
);

INVx1_ASAP7_75t_L g20814 ( 
.A(n_20557),
.Y(n_20814)
);

OAI221xp5_ASAP7_75t_L g20815 ( 
.A1(n_20778),
.A2(n_8988),
.B1(n_9300),
.B2(n_9339),
.C(n_9293),
.Y(n_20815)
);

OAI21xp5_ASAP7_75t_SL g20816 ( 
.A1(n_20632),
.A2(n_9300),
.B(n_9293),
.Y(n_20816)
);

NOR2xp33_ASAP7_75t_L g20817 ( 
.A(n_20776),
.B(n_10032),
.Y(n_20817)
);

NAND2xp5_ASAP7_75t_L g20818 ( 
.A(n_20627),
.B(n_10546),
.Y(n_20818)
);

INVx1_ASAP7_75t_L g20819 ( 
.A(n_20653),
.Y(n_20819)
);

OAI211xp5_ASAP7_75t_L g20820 ( 
.A1(n_20645),
.A2(n_10917),
.B(n_10051),
.C(n_10032),
.Y(n_20820)
);

AOI21xp5_ASAP7_75t_L g20821 ( 
.A1(n_20760),
.A2(n_10407),
.B(n_10405),
.Y(n_20821)
);

OAI211xp5_ASAP7_75t_L g20822 ( 
.A1(n_20730),
.A2(n_10917),
.B(n_10051),
.C(n_10032),
.Y(n_20822)
);

AOI22xp33_ASAP7_75t_L g20823 ( 
.A1(n_20577),
.A2(n_10206),
.B1(n_10225),
.B2(n_10202),
.Y(n_20823)
);

OAI211xp5_ASAP7_75t_SL g20824 ( 
.A1(n_20744),
.A2(n_9980),
.B(n_9988),
.C(n_9979),
.Y(n_20824)
);

AOI22xp5_ASAP7_75t_L g20825 ( 
.A1(n_20729),
.A2(n_11300),
.B1(n_10989),
.B2(n_10998),
.Y(n_20825)
);

OAI211xp5_ASAP7_75t_SL g20826 ( 
.A1(n_20722),
.A2(n_9980),
.B(n_9988),
.C(n_9979),
.Y(n_20826)
);

NAND3xp33_ASAP7_75t_L g20827 ( 
.A(n_20698),
.B(n_10051),
.C(n_10032),
.Y(n_20827)
);

OAI211xp5_ASAP7_75t_L g20828 ( 
.A1(n_20642),
.A2(n_10051),
.B(n_10032),
.C(n_11504),
.Y(n_20828)
);

O2A1O1Ixp5_ASAP7_75t_SL g20829 ( 
.A1(n_20709),
.A2(n_9041),
.B(n_9053),
.C(n_9045),
.Y(n_20829)
);

AOI221xp5_ASAP7_75t_L g20830 ( 
.A1(n_20608),
.A2(n_10006),
.B1(n_9828),
.B2(n_9571),
.C(n_9651),
.Y(n_20830)
);

AOI22xp5_ASAP7_75t_SL g20831 ( 
.A1(n_20705),
.A2(n_10184),
.B1(n_9513),
.B2(n_9496),
.Y(n_20831)
);

AOI22xp5_ASAP7_75t_L g20832 ( 
.A1(n_20723),
.A2(n_10989),
.B1(n_10998),
.B2(n_10979),
.Y(n_20832)
);

OAI31xp33_ASAP7_75t_L g20833 ( 
.A1(n_20701),
.A2(n_9339),
.A3(n_9358),
.B(n_9293),
.Y(n_20833)
);

AOI22xp5_ASAP7_75t_L g20834 ( 
.A1(n_20568),
.A2(n_10989),
.B1(n_10998),
.B2(n_10979),
.Y(n_20834)
);

AOI211xp5_ASAP7_75t_L g20835 ( 
.A1(n_20607),
.A2(n_10629),
.B(n_11570),
.C(n_10560),
.Y(n_20835)
);

INVxp67_ASAP7_75t_L g20836 ( 
.A(n_20753),
.Y(n_20836)
);

AOI31xp33_ASAP7_75t_L g20837 ( 
.A1(n_20655),
.A2(n_9339),
.A3(n_9378),
.B(n_9358),
.Y(n_20837)
);

OAI211xp5_ASAP7_75t_SL g20838 ( 
.A1(n_20770),
.A2(n_9992),
.B(n_10008),
.C(n_9988),
.Y(n_20838)
);

OAI221xp5_ASAP7_75t_L g20839 ( 
.A1(n_20713),
.A2(n_8988),
.B1(n_9358),
.B2(n_9378),
.C(n_9339),
.Y(n_20839)
);

AOI22xp5_ASAP7_75t_L g20840 ( 
.A1(n_20740),
.A2(n_10989),
.B1(n_10998),
.B2(n_10979),
.Y(n_20840)
);

AOI221xp5_ASAP7_75t_L g20841 ( 
.A1(n_20758),
.A2(n_9575),
.B1(n_9651),
.B2(n_9571),
.C(n_9883),
.Y(n_20841)
);

NOR2xp33_ASAP7_75t_SL g20842 ( 
.A(n_20654),
.B(n_10032),
.Y(n_20842)
);

AOI21xp5_ASAP7_75t_L g20843 ( 
.A1(n_20704),
.A2(n_10407),
.B(n_10405),
.Y(n_20843)
);

OAI21xp33_ASAP7_75t_SL g20844 ( 
.A1(n_20556),
.A2(n_10398),
.B(n_10397),
.Y(n_20844)
);

NAND3xp33_ASAP7_75t_L g20845 ( 
.A(n_20735),
.B(n_10051),
.C(n_10032),
.Y(n_20845)
);

NOR4xp25_ASAP7_75t_L g20846 ( 
.A(n_20667),
.B(n_9042),
.C(n_9052),
.D(n_9043),
.Y(n_20846)
);

AOI211xp5_ASAP7_75t_SL g20847 ( 
.A1(n_20684),
.A2(n_9053),
.B(n_9055),
.C(n_9045),
.Y(n_20847)
);

O2A1O1Ixp33_ASAP7_75t_L g20848 ( 
.A1(n_20689),
.A2(n_9239),
.B(n_9268),
.C(n_8636),
.Y(n_20848)
);

AOI221xp5_ASAP7_75t_L g20849 ( 
.A1(n_20620),
.A2(n_9575),
.B1(n_9651),
.B2(n_9571),
.C(n_9883),
.Y(n_20849)
);

AOI22xp33_ASAP7_75t_L g20850 ( 
.A1(n_20657),
.A2(n_10206),
.B1(n_10225),
.B2(n_10202),
.Y(n_20850)
);

AND2x2_ASAP7_75t_L g20851 ( 
.A(n_20679),
.B(n_8597),
.Y(n_20851)
);

AOI32xp33_ASAP7_75t_L g20852 ( 
.A1(n_20726),
.A2(n_11406),
.A3(n_11417),
.B1(n_11415),
.B2(n_11398),
.Y(n_20852)
);

AOI221xp5_ASAP7_75t_L g20853 ( 
.A1(n_20619),
.A2(n_9575),
.B1(n_9651),
.B2(n_9571),
.C(n_9883),
.Y(n_20853)
);

AOI322xp5_ASAP7_75t_L g20854 ( 
.A1(n_20761),
.A2(n_9355),
.A3(n_9316),
.B1(n_9356),
.B2(n_9366),
.C1(n_9348),
.C2(n_9302),
.Y(n_20854)
);

OAI221xp5_ASAP7_75t_SL g20855 ( 
.A1(n_20581),
.A2(n_10103),
.B1(n_10002),
.B2(n_9900),
.C(n_10121),
.Y(n_20855)
);

AOI21xp33_ASAP7_75t_L g20856 ( 
.A1(n_20575),
.A2(n_10989),
.B(n_10979),
.Y(n_20856)
);

NOR2xp33_ASAP7_75t_L g20857 ( 
.A(n_20668),
.B(n_10032),
.Y(n_20857)
);

NOR2x1p5_ASAP7_75t_L g20858 ( 
.A(n_20583),
.B(n_8734),
.Y(n_20858)
);

AND3x4_ASAP7_75t_L g20859 ( 
.A(n_20665),
.B(n_9575),
.C(n_9571),
.Y(n_20859)
);

AOI22xp5_ASAP7_75t_L g20860 ( 
.A1(n_20606),
.A2(n_10998),
.B1(n_11048),
.B2(n_10979),
.Y(n_20860)
);

OAI211xp5_ASAP7_75t_L g20861 ( 
.A1(n_20591),
.A2(n_10051),
.B(n_11506),
.C(n_11504),
.Y(n_20861)
);

AOI21xp5_ASAP7_75t_L g20862 ( 
.A1(n_20624),
.A2(n_10407),
.B(n_10405),
.Y(n_20862)
);

AOI221xp5_ASAP7_75t_L g20863 ( 
.A1(n_20658),
.A2(n_9575),
.B1(n_9651),
.B2(n_9571),
.C(n_9883),
.Y(n_20863)
);

AOI211xp5_ASAP7_75t_L g20864 ( 
.A1(n_20614),
.A2(n_10560),
.B(n_10551),
.C(n_8636),
.Y(n_20864)
);

OAI31xp33_ASAP7_75t_L g20865 ( 
.A1(n_20767),
.A2(n_9358),
.A3(n_9378),
.B(n_9339),
.Y(n_20865)
);

AOI21xp5_ASAP7_75t_L g20866 ( 
.A1(n_20615),
.A2(n_10411),
.B(n_10390),
.Y(n_20866)
);

NAND3xp33_ASAP7_75t_SL g20867 ( 
.A(n_20777),
.B(n_20750),
.C(n_20773),
.Y(n_20867)
);

AOI211x1_ASAP7_75t_SL g20868 ( 
.A1(n_20690),
.A2(n_9043),
.B(n_9052),
.C(n_9042),
.Y(n_20868)
);

NOR2xp33_ASAP7_75t_L g20869 ( 
.A(n_20664),
.B(n_20617),
.Y(n_20869)
);

AOI21xp5_ASAP7_75t_L g20870 ( 
.A1(n_20727),
.A2(n_10411),
.B(n_10390),
.Y(n_20870)
);

AOI221xp5_ASAP7_75t_L g20871 ( 
.A1(n_20609),
.A2(n_9651),
.B1(n_9575),
.B2(n_9883),
.C(n_9510),
.Y(n_20871)
);

AOI21xp5_ASAP7_75t_L g20872 ( 
.A1(n_20746),
.A2(n_10411),
.B(n_10390),
.Y(n_20872)
);

NOR2xp33_ASAP7_75t_SL g20873 ( 
.A(n_20638),
.B(n_10051),
.Y(n_20873)
);

NAND2xp5_ASAP7_75t_L g20874 ( 
.A(n_20647),
.B(n_10546),
.Y(n_20874)
);

OAI221xp5_ASAP7_75t_SL g20875 ( 
.A1(n_20590),
.A2(n_10103),
.B1(n_10002),
.B2(n_9900),
.C(n_10121),
.Y(n_20875)
);

AOI22xp5_ASAP7_75t_L g20876 ( 
.A1(n_20647),
.A2(n_10998),
.B1(n_11048),
.B2(n_10979),
.Y(n_20876)
);

OAI21xp5_ASAP7_75t_SL g20877 ( 
.A1(n_20644),
.A2(n_20702),
.B(n_20597),
.Y(n_20877)
);

NOR3xp33_ASAP7_75t_L g20878 ( 
.A(n_20721),
.B(n_20634),
.C(n_20637),
.Y(n_20878)
);

AOI22xp5_ASAP7_75t_L g20879 ( 
.A1(n_20610),
.A2(n_11062),
.B1(n_11084),
.B2(n_11048),
.Y(n_20879)
);

AOI221x1_ASAP7_75t_L g20880 ( 
.A1(n_20633),
.A2(n_20683),
.B1(n_20631),
.B2(n_20589),
.C(n_20592),
.Y(n_20880)
);

AOI222xp33_ASAP7_75t_L g20881 ( 
.A1(n_20629),
.A2(n_20651),
.B1(n_20678),
.B2(n_20763),
.C1(n_20772),
.C2(n_20600),
.Y(n_20881)
);

INVx1_ASAP7_75t_L g20882 ( 
.A(n_20659),
.Y(n_20882)
);

NOR3xp33_ASAP7_75t_L g20883 ( 
.A(n_20703),
.B(n_10822),
.C(n_11398),
.Y(n_20883)
);

AOI211xp5_ASAP7_75t_L g20884 ( 
.A1(n_20712),
.A2(n_10560),
.B(n_10551),
.C(n_8636),
.Y(n_20884)
);

AOI221xp5_ASAP7_75t_L g20885 ( 
.A1(n_20661),
.A2(n_20743),
.B1(n_20595),
.B2(n_20759),
.C(n_20584),
.Y(n_20885)
);

AOI221xp5_ASAP7_75t_L g20886 ( 
.A1(n_20765),
.A2(n_9651),
.B1(n_9575),
.B2(n_9883),
.C(n_9510),
.Y(n_20886)
);

AOI222xp33_ASAP7_75t_SL g20887 ( 
.A1(n_20749),
.A2(n_9835),
.B1(n_9070),
.B2(n_9053),
.C1(n_9081),
.C2(n_9055),
.Y(n_20887)
);

AOI21xp5_ASAP7_75t_L g20888 ( 
.A1(n_20733),
.A2(n_20751),
.B(n_20593),
.Y(n_20888)
);

NOR2xp33_ASAP7_75t_L g20889 ( 
.A(n_20630),
.B(n_20755),
.Y(n_20889)
);

OAI211xp5_ASAP7_75t_SL g20890 ( 
.A1(n_20681),
.A2(n_10008),
.B(n_10028),
.C(n_9992),
.Y(n_20890)
);

AOI22xp33_ASAP7_75t_L g20891 ( 
.A1(n_20782),
.A2(n_10206),
.B1(n_10225),
.B2(n_10202),
.Y(n_20891)
);

NAND2xp5_ASAP7_75t_SL g20892 ( 
.A(n_20671),
.B(n_10051),
.Y(n_20892)
);

AOI211xp5_ASAP7_75t_L g20893 ( 
.A1(n_20696),
.A2(n_10551),
.B(n_8636),
.C(n_8660),
.Y(n_20893)
);

NOR3xp33_ASAP7_75t_L g20894 ( 
.A(n_20626),
.B(n_10822),
.C(n_11406),
.Y(n_20894)
);

OAI32xp33_ASAP7_75t_L g20895 ( 
.A1(n_20567),
.A2(n_9042),
.A3(n_9071),
.B1(n_9052),
.B2(n_9043),
.Y(n_20895)
);

OAI211xp5_ASAP7_75t_L g20896 ( 
.A1(n_20621),
.A2(n_10051),
.B(n_11506),
.C(n_10184),
.Y(n_20896)
);

AOI21xp5_ASAP7_75t_L g20897 ( 
.A1(n_20720),
.A2(n_10391),
.B(n_10384),
.Y(n_20897)
);

OAI22xp5_ASAP7_75t_L g20898 ( 
.A1(n_20564),
.A2(n_9053),
.B1(n_9055),
.B2(n_9045),
.Y(n_20898)
);

OAI321xp33_ASAP7_75t_L g20899 ( 
.A1(n_20774),
.A2(n_9454),
.A3(n_9358),
.B1(n_9464),
.B2(n_9378),
.C(n_9339),
.Y(n_20899)
);

AOI211x1_ASAP7_75t_L g20900 ( 
.A1(n_20775),
.A2(n_9070),
.B(n_9081),
.C(n_9055),
.Y(n_20900)
);

AOI211xp5_ASAP7_75t_L g20901 ( 
.A1(n_20649),
.A2(n_8636),
.B(n_8660),
.C(n_8374),
.Y(n_20901)
);

NAND2xp5_ASAP7_75t_L g20902 ( 
.A(n_20708),
.B(n_10557),
.Y(n_20902)
);

AOI21x1_ASAP7_75t_L g20903 ( 
.A1(n_20618),
.A2(n_10951),
.B(n_10946),
.Y(n_20903)
);

INVx2_ASAP7_75t_L g20904 ( 
.A(n_20706),
.Y(n_20904)
);

NAND4xp75_ASAP7_75t_L g20905 ( 
.A(n_20747),
.B(n_10202),
.C(n_10225),
.D(n_10206),
.Y(n_20905)
);

INVx1_ASAP7_75t_L g20906 ( 
.A(n_20745),
.Y(n_20906)
);

AOI22xp5_ASAP7_75t_L g20907 ( 
.A1(n_20685),
.A2(n_11062),
.B1(n_11084),
.B2(n_11048),
.Y(n_20907)
);

O2A1O1Ixp33_ASAP7_75t_L g20908 ( 
.A1(n_20604),
.A2(n_9239),
.B(n_9268),
.C(n_8660),
.Y(n_20908)
);

AOI21xp33_ASAP7_75t_L g20909 ( 
.A1(n_20748),
.A2(n_11062),
.B(n_11048),
.Y(n_20909)
);

AOI311xp33_ASAP7_75t_L g20910 ( 
.A1(n_20741),
.A2(n_9096),
.A3(n_9100),
.B(n_9081),
.C(n_9070),
.Y(n_20910)
);

AOI221xp5_ASAP7_75t_L g20911 ( 
.A1(n_20674),
.A2(n_9651),
.B1(n_9575),
.B2(n_9883),
.C(n_9520),
.Y(n_20911)
);

AOI211xp5_ASAP7_75t_L g20912 ( 
.A1(n_20643),
.A2(n_8660),
.B(n_8374),
.C(n_11398),
.Y(n_20912)
);

NAND2xp33_ASAP7_75t_SL g20913 ( 
.A(n_20739),
.B(n_8248),
.Y(n_20913)
);

OAI21xp33_ASAP7_75t_L g20914 ( 
.A1(n_20728),
.A2(n_9883),
.B(n_9992),
.Y(n_20914)
);

A2O1A1Ixp33_ASAP7_75t_L g20915 ( 
.A1(n_20561),
.A2(n_20669),
.B(n_20648),
.C(n_20586),
.Y(n_20915)
);

AOI22xp5_ASAP7_75t_L g20916 ( 
.A1(n_20562),
.A2(n_20732),
.B1(n_20559),
.B2(n_20594),
.Y(n_20916)
);

AOI22xp5_ASAP7_75t_L g20917 ( 
.A1(n_20565),
.A2(n_11062),
.B1(n_11084),
.B2(n_11048),
.Y(n_20917)
);

AOI221xp5_ASAP7_75t_L g20918 ( 
.A1(n_20623),
.A2(n_9575),
.B1(n_9883),
.B2(n_9520),
.C(n_9510),
.Y(n_20918)
);

AOI322xp5_ASAP7_75t_L g20919 ( 
.A1(n_20710),
.A2(n_9355),
.A3(n_9316),
.B1(n_9356),
.B2(n_9366),
.C1(n_9348),
.C2(n_9302),
.Y(n_20919)
);

AND2x2_ASAP7_75t_L g20920 ( 
.A(n_20724),
.B(n_8597),
.Y(n_20920)
);

NAND4xp25_ASAP7_75t_SL g20921 ( 
.A(n_20663),
.B(n_9081),
.C(n_9096),
.D(n_9070),
.Y(n_20921)
);

NAND2xp5_ASAP7_75t_L g20922 ( 
.A(n_20687),
.B(n_10557),
.Y(n_20922)
);

OAI22xp33_ASAP7_75t_L g20923 ( 
.A1(n_20628),
.A2(n_9100),
.B1(n_9103),
.B2(n_9096),
.Y(n_20923)
);

NAND2xp5_ASAP7_75t_L g20924 ( 
.A(n_20697),
.B(n_10557),
.Y(n_20924)
);

NAND2xp33_ASAP7_75t_R g20925 ( 
.A(n_20602),
.B(n_10184),
.Y(n_20925)
);

A2O1A1Ixp33_ASAP7_75t_SL g20926 ( 
.A1(n_20686),
.A2(n_9043),
.B(n_9052),
.C(n_9042),
.Y(n_20926)
);

AOI221xp5_ASAP7_75t_L g20927 ( 
.A1(n_20757),
.A2(n_9520),
.B1(n_9510),
.B2(n_9146),
.C(n_9183),
.Y(n_20927)
);

AOI21xp5_ASAP7_75t_L g20928 ( 
.A1(n_20694),
.A2(n_10391),
.B(n_10384),
.Y(n_20928)
);

NAND4xp25_ASAP7_75t_L g20929 ( 
.A(n_20742),
.B(n_8745),
.C(n_8815),
.D(n_8734),
.Y(n_20929)
);

NOR2x1_ASAP7_75t_L g20930 ( 
.A(n_20707),
.B(n_20682),
.Y(n_20930)
);

NAND4xp25_ASAP7_75t_SL g20931 ( 
.A(n_20613),
.B(n_9100),
.C(n_9103),
.D(n_9096),
.Y(n_20931)
);

NAND2xp5_ASAP7_75t_L g20932 ( 
.A(n_20736),
.B(n_20692),
.Y(n_20932)
);

OAI211xp5_ASAP7_75t_SL g20933 ( 
.A1(n_20571),
.A2(n_10028),
.B(n_10030),
.C(n_10008),
.Y(n_20933)
);

A2O1A1Ixp33_ASAP7_75t_L g20934 ( 
.A1(n_20673),
.A2(n_20693),
.B(n_20680),
.C(n_20779),
.Y(n_20934)
);

AOI22xp5_ASAP7_75t_L g20935 ( 
.A1(n_20662),
.A2(n_11084),
.B1(n_11062),
.B2(n_11089),
.Y(n_20935)
);

AOI221xp5_ASAP7_75t_L g20936 ( 
.A1(n_20656),
.A2(n_9510),
.B1(n_9520),
.B2(n_9222),
.C(n_9182),
.Y(n_20936)
);

NAND2x1_ASAP7_75t_L g20937 ( 
.A(n_20754),
.B(n_9835),
.Y(n_20937)
);

NOR3xp33_ASAP7_75t_L g20938 ( 
.A(n_20766),
.B(n_11417),
.C(n_11415),
.Y(n_20938)
);

NAND3xp33_ASAP7_75t_SL g20939 ( 
.A(n_20688),
.B(n_9378),
.C(n_9358),
.Y(n_20939)
);

OAI321xp33_ASAP7_75t_L g20940 ( 
.A1(n_20764),
.A2(n_9535),
.A3(n_9454),
.B1(n_9540),
.B2(n_9464),
.C(n_9378),
.Y(n_20940)
);

AOI21xp5_ASAP7_75t_L g20941 ( 
.A1(n_20574),
.A2(n_20578),
.B(n_20691),
.Y(n_20941)
);

INVx2_ASAP7_75t_SL g20942 ( 
.A(n_20641),
.Y(n_20942)
);

OAI321xp33_ASAP7_75t_L g20943 ( 
.A1(n_20718),
.A2(n_9540),
.A3(n_9464),
.B1(n_9643),
.B2(n_9535),
.C(n_9454),
.Y(n_20943)
);

OR2x2_ASAP7_75t_L g20944 ( 
.A(n_20640),
.B(n_10557),
.Y(n_20944)
);

NOR3xp33_ASAP7_75t_L g20945 ( 
.A(n_20570),
.B(n_11417),
.C(n_11415),
.Y(n_20945)
);

INVx2_ASAP7_75t_L g20946 ( 
.A(n_20676),
.Y(n_20946)
);

AOI22xp5_ASAP7_75t_SL g20947 ( 
.A1(n_20700),
.A2(n_10184),
.B1(n_9513),
.B2(n_9496),
.Y(n_20947)
);

AOI322xp5_ASAP7_75t_L g20948 ( 
.A1(n_20563),
.A2(n_9355),
.A3(n_9316),
.B1(n_9356),
.B2(n_9366),
.C1(n_9348),
.C2(n_9302),
.Y(n_20948)
);

NOR2xp33_ASAP7_75t_L g20949 ( 
.A(n_20677),
.B(n_11062),
.Y(n_20949)
);

OAI221xp5_ASAP7_75t_L g20950 ( 
.A1(n_20738),
.A2(n_9454),
.B1(n_9644),
.B2(n_9643),
.C(n_9540),
.Y(n_20950)
);

AOI221xp5_ASAP7_75t_L g20951 ( 
.A1(n_20660),
.A2(n_9520),
.B1(n_9510),
.B2(n_9400),
.C(n_9222),
.Y(n_20951)
);

OAI21xp33_ASAP7_75t_L g20952 ( 
.A1(n_20588),
.A2(n_10028),
.B(n_10008),
.Y(n_20952)
);

OR2x2_ASAP7_75t_L g20953 ( 
.A(n_20599),
.B(n_10557),
.Y(n_20953)
);

O2A1O1Ixp33_ASAP7_75t_L g20954 ( 
.A1(n_20601),
.A2(n_9239),
.B(n_8660),
.C(n_8374),
.Y(n_20954)
);

OA21x2_ASAP7_75t_L g20955 ( 
.A1(n_20716),
.A2(n_10391),
.B(n_10384),
.Y(n_20955)
);

OAI221xp5_ASAP7_75t_L g20956 ( 
.A1(n_20734),
.A2(n_9454),
.B1(n_9643),
.B2(n_9535),
.C(n_9464),
.Y(n_20956)
);

OAI211xp5_ASAP7_75t_L g20957 ( 
.A1(n_20670),
.A2(n_10184),
.B(n_9925),
.C(n_9916),
.Y(n_20957)
);

OAI221xp5_ASAP7_75t_SL g20958 ( 
.A1(n_20711),
.A2(n_10103),
.B1(n_10002),
.B2(n_9900),
.C(n_10121),
.Y(n_20958)
);

NAND3xp33_ASAP7_75t_L g20959 ( 
.A(n_20585),
.B(n_11084),
.C(n_9925),
.Y(n_20959)
);

NAND2xp5_ASAP7_75t_SL g20960 ( 
.A(n_20714),
.B(n_9965),
.Y(n_20960)
);

AOI211x1_ASAP7_75t_L g20961 ( 
.A1(n_20695),
.A2(n_9103),
.B(n_9128),
.C(n_9100),
.Y(n_20961)
);

OAI221xp5_ASAP7_75t_SL g20962 ( 
.A1(n_20719),
.A2(n_10103),
.B1(n_10002),
.B2(n_9900),
.C(n_10121),
.Y(n_20962)
);

NAND2xp5_ASAP7_75t_L g20963 ( 
.A(n_20652),
.B(n_10557),
.Y(n_20963)
);

AOI21x1_ASAP7_75t_L g20964 ( 
.A1(n_20635),
.A2(n_10951),
.B(n_10946),
.Y(n_20964)
);

AOI21xp33_ASAP7_75t_SL g20965 ( 
.A1(n_20611),
.A2(n_9925),
.B(n_9916),
.Y(n_20965)
);

AOI211xp5_ASAP7_75t_L g20966 ( 
.A1(n_20715),
.A2(n_8374),
.B(n_11426),
.C(n_11425),
.Y(n_20966)
);

AOI21xp33_ASAP7_75t_SL g20967 ( 
.A1(n_20622),
.A2(n_9925),
.B(n_9916),
.Y(n_20967)
);

A2O1A1Ixp33_ASAP7_75t_L g20968 ( 
.A1(n_20580),
.A2(n_10398),
.B(n_10397),
.C(n_10320),
.Y(n_20968)
);

OAI211xp5_ASAP7_75t_L g20969 ( 
.A1(n_20596),
.A2(n_20666),
.B(n_20699),
.C(n_20717),
.Y(n_20969)
);

AOI221xp5_ASAP7_75t_L g20970 ( 
.A1(n_20612),
.A2(n_9520),
.B1(n_9510),
.B2(n_9183),
.C(n_9311),
.Y(n_20970)
);

NOR2x1_ASAP7_75t_L g20971 ( 
.A(n_20771),
.B(n_10184),
.Y(n_20971)
);

OAI321xp33_ASAP7_75t_L g20972 ( 
.A1(n_20675),
.A2(n_9540),
.A3(n_9464),
.B1(n_9643),
.B2(n_9535),
.C(n_9454),
.Y(n_20972)
);

AOI21xp5_ASAP7_75t_L g20973 ( 
.A1(n_20612),
.A2(n_10320),
.B(n_10316),
.Y(n_20973)
);

INVx1_ASAP7_75t_L g20974 ( 
.A(n_20569),
.Y(n_20974)
);

NAND2xp5_ASAP7_75t_L g20975 ( 
.A(n_20560),
.B(n_10557),
.Y(n_20975)
);

NAND2x1_ASAP7_75t_L g20976 ( 
.A(n_20650),
.B(n_9835),
.Y(n_20976)
);

NOR2xp33_ASAP7_75t_R g20977 ( 
.A(n_20616),
.B(n_7782),
.Y(n_20977)
);

AO221x1_ASAP7_75t_L g20978 ( 
.A1(n_20566),
.A2(n_8296),
.B1(n_8314),
.B2(n_8273),
.C(n_8248),
.Y(n_20978)
);

NAND3xp33_ASAP7_75t_L g20979 ( 
.A(n_20573),
.B(n_11084),
.C(n_9925),
.Y(n_20979)
);

NAND2xp5_ASAP7_75t_L g20980 ( 
.A(n_20560),
.B(n_10557),
.Y(n_20980)
);

OAI22xp5_ASAP7_75t_L g20981 ( 
.A1(n_20579),
.A2(n_9128),
.B1(n_9132),
.B2(n_9103),
.Y(n_20981)
);

NOR2xp33_ASAP7_75t_L g20982 ( 
.A(n_20569),
.B(n_9916),
.Y(n_20982)
);

AOI211x1_ASAP7_75t_SL g20983 ( 
.A1(n_20566),
.A2(n_9071),
.B(n_9107),
.C(n_9042),
.Y(n_20983)
);

AOI221xp5_ASAP7_75t_SL g20984 ( 
.A1(n_20612),
.A2(n_9133),
.B1(n_9147),
.B2(n_9132),
.C(n_9128),
.Y(n_20984)
);

NAND2xp5_ASAP7_75t_L g20985 ( 
.A(n_20798),
.B(n_20974),
.Y(n_20985)
);

NAND3xp33_ASAP7_75t_SL g20986 ( 
.A(n_20810),
.B(n_9464),
.C(n_9454),
.Y(n_20986)
);

AND2x2_ASAP7_75t_L g20987 ( 
.A(n_20920),
.B(n_20851),
.Y(n_20987)
);

OAI22xp5_ASAP7_75t_L g20988 ( 
.A1(n_20836),
.A2(n_20845),
.B1(n_20979),
.B2(n_20803),
.Y(n_20988)
);

NAND3xp33_ASAP7_75t_L g20989 ( 
.A(n_20869),
.B(n_9925),
.C(n_9916),
.Y(n_20989)
);

INVx1_ASAP7_75t_L g20990 ( 
.A(n_20930),
.Y(n_20990)
);

NOR2x1_ASAP7_75t_L g20991 ( 
.A(n_20882),
.B(n_10184),
.Y(n_20991)
);

NAND2xp5_ASAP7_75t_L g20992 ( 
.A(n_20786),
.B(n_9288),
.Y(n_20992)
);

NOR2xp33_ASAP7_75t_L g20993 ( 
.A(n_20867),
.B(n_9916),
.Y(n_20993)
);

AOI221x1_ASAP7_75t_L g20994 ( 
.A1(n_20814),
.A2(n_10035),
.B1(n_10046),
.B2(n_10030),
.C(n_10028),
.Y(n_20994)
);

NAND3xp33_ASAP7_75t_L g20995 ( 
.A(n_20889),
.B(n_9925),
.C(n_9916),
.Y(n_20995)
);

NAND2xp5_ASAP7_75t_SL g20996 ( 
.A(n_20788),
.B(n_9965),
.Y(n_20996)
);

NAND2xp5_ASAP7_75t_L g20997 ( 
.A(n_20817),
.B(n_9288),
.Y(n_20997)
);

XNOR2xp5_ASAP7_75t_L g20998 ( 
.A(n_20969),
.B(n_8454),
.Y(n_20998)
);

INVxp67_ASAP7_75t_L g20999 ( 
.A(n_20946),
.Y(n_20999)
);

INVx1_ASAP7_75t_L g21000 ( 
.A(n_20916),
.Y(n_21000)
);

INVx1_ASAP7_75t_L g21001 ( 
.A(n_20892),
.Y(n_21001)
);

INVxp67_ASAP7_75t_SL g21002 ( 
.A(n_20942),
.Y(n_21002)
);

AOI21xp5_ASAP7_75t_L g21003 ( 
.A1(n_20843),
.A2(n_10687),
.B(n_10680),
.Y(n_21003)
);

NAND2xp5_ASAP7_75t_L g21004 ( 
.A(n_20881),
.B(n_9288),
.Y(n_21004)
);

NAND2xp5_ASAP7_75t_L g21005 ( 
.A(n_20819),
.B(n_9288),
.Y(n_21005)
);

AND2x2_ASAP7_75t_L g21006 ( 
.A(n_20878),
.B(n_9616),
.Y(n_21006)
);

OAI21xp33_ASAP7_75t_L g21007 ( 
.A1(n_20857),
.A2(n_9182),
.B(n_9146),
.Y(n_21007)
);

NOR2x1_ASAP7_75t_L g21008 ( 
.A(n_20904),
.B(n_10184),
.Y(n_21008)
);

NOR2xp67_ASAP7_75t_L g21009 ( 
.A(n_20941),
.B(n_8735),
.Y(n_21009)
);

NAND4xp25_ASAP7_75t_L g21010 ( 
.A(n_20880),
.B(n_8815),
.C(n_8821),
.D(n_8745),
.Y(n_21010)
);

AOI21xp5_ASAP7_75t_L g21011 ( 
.A1(n_20888),
.A2(n_10687),
.B(n_10680),
.Y(n_21011)
);

NOR2xp67_ASAP7_75t_L g21012 ( 
.A(n_20827),
.B(n_8735),
.Y(n_21012)
);

NAND4xp25_ASAP7_75t_L g21013 ( 
.A(n_20885),
.B(n_8815),
.C(n_8821),
.D(n_8745),
.Y(n_21013)
);

INVx1_ASAP7_75t_L g21014 ( 
.A(n_20932),
.Y(n_21014)
);

HB1xp67_ASAP7_75t_L g21015 ( 
.A(n_20858),
.Y(n_21015)
);

AND2x2_ASAP7_75t_L g21016 ( 
.A(n_20978),
.B(n_9616),
.Y(n_21016)
);

INVx1_ASAP7_75t_L g21017 ( 
.A(n_20934),
.Y(n_21017)
);

NAND2xp5_ASAP7_75t_L g21018 ( 
.A(n_20915),
.B(n_9288),
.Y(n_21018)
);

INVx1_ASAP7_75t_L g21019 ( 
.A(n_20877),
.Y(n_21019)
);

NAND2xp5_ASAP7_75t_L g21020 ( 
.A(n_20983),
.B(n_9288),
.Y(n_21020)
);

AOI22xp5_ASAP7_75t_L g21021 ( 
.A1(n_20842),
.A2(n_11094),
.B1(n_11089),
.B2(n_10296),
.Y(n_21021)
);

NOR3xp33_ASAP7_75t_L g21022 ( 
.A(n_20906),
.B(n_10824),
.C(n_10823),
.Y(n_21022)
);

NOR2x1_ASAP7_75t_L g21023 ( 
.A(n_20976),
.B(n_10184),
.Y(n_21023)
);

AOI222xp33_ASAP7_75t_L g21024 ( 
.A1(n_20807),
.A2(n_10580),
.B1(n_10532),
.B2(n_10534),
.C1(n_10548),
.C2(n_10533),
.Y(n_21024)
);

NAND4xp25_ASAP7_75t_L g21025 ( 
.A(n_20873),
.B(n_8821),
.C(n_8826),
.D(n_8745),
.Y(n_21025)
);

NAND4xp25_ASAP7_75t_L g21026 ( 
.A(n_20913),
.B(n_8826),
.C(n_8821),
.D(n_8997),
.Y(n_21026)
);

INVx1_ASAP7_75t_SL g21027 ( 
.A(n_20811),
.Y(n_21027)
);

NAND2xp5_ASAP7_75t_L g21028 ( 
.A(n_20868),
.B(n_9288),
.Y(n_21028)
);

INVxp67_ASAP7_75t_L g21029 ( 
.A(n_20960),
.Y(n_21029)
);

INVx1_ASAP7_75t_L g21030 ( 
.A(n_20859),
.Y(n_21030)
);

NAND2xp5_ASAP7_75t_L g21031 ( 
.A(n_20949),
.B(n_9288),
.Y(n_21031)
);

AND2x2_ASAP7_75t_L g21032 ( 
.A(n_20977),
.B(n_9616),
.Y(n_21032)
);

INVx1_ASAP7_75t_L g21033 ( 
.A(n_20902),
.Y(n_21033)
);

OAI31xp33_ASAP7_75t_SL g21034 ( 
.A1(n_20971),
.A2(n_10533),
.A3(n_10534),
.B(n_10532),
.Y(n_21034)
);

INVx1_ASAP7_75t_L g21035 ( 
.A(n_20975),
.Y(n_21035)
);

NOR3xp33_ASAP7_75t_SL g21036 ( 
.A(n_20929),
.B(n_8735),
.C(n_8592),
.Y(n_21036)
);

CKINVDCx20_ASAP7_75t_L g21037 ( 
.A(n_20925),
.Y(n_21037)
);

AND2x2_ASAP7_75t_L g21038 ( 
.A(n_20980),
.B(n_9616),
.Y(n_21038)
);

NOR2xp33_ASAP7_75t_L g21039 ( 
.A(n_20914),
.B(n_9916),
.Y(n_21039)
);

OAI22xp5_ASAP7_75t_L g21040 ( 
.A1(n_20825),
.A2(n_9132),
.B1(n_9133),
.B2(n_9128),
.Y(n_21040)
);

NOR3xp33_ASAP7_75t_L g21041 ( 
.A(n_20982),
.B(n_10824),
.C(n_10823),
.Y(n_21041)
);

INVx1_ASAP7_75t_L g21042 ( 
.A(n_20818),
.Y(n_21042)
);

NOR2xp33_ASAP7_75t_L g21043 ( 
.A(n_20937),
.B(n_9916),
.Y(n_21043)
);

INVx1_ASAP7_75t_L g21044 ( 
.A(n_20874),
.Y(n_21044)
);

NAND2xp5_ASAP7_75t_L g21045 ( 
.A(n_20865),
.B(n_9965),
.Y(n_21045)
);

AND2x2_ASAP7_75t_L g21046 ( 
.A(n_20912),
.B(n_9616),
.Y(n_21046)
);

AOI211xp5_ASAP7_75t_L g21047 ( 
.A1(n_20838),
.A2(n_8374),
.B(n_10276),
.C(n_10256),
.Y(n_21047)
);

AOI22xp5_ASAP7_75t_L g21048 ( 
.A1(n_20790),
.A2(n_11094),
.B1(n_11089),
.B2(n_10296),
.Y(n_21048)
);

AND2x2_ASAP7_75t_L g21049 ( 
.A(n_20830),
.B(n_8597),
.Y(n_21049)
);

AOI221xp5_ASAP7_75t_L g21050 ( 
.A1(n_20967),
.A2(n_9520),
.B1(n_9510),
.B2(n_9147),
.C(n_9155),
.Y(n_21050)
);

INVx2_ASAP7_75t_L g21051 ( 
.A(n_20944),
.Y(n_21051)
);

AOI21xp5_ASAP7_75t_L g21052 ( 
.A1(n_20787),
.A2(n_10687),
.B(n_10680),
.Y(n_21052)
);

NAND2xp5_ASAP7_75t_SL g21053 ( 
.A(n_20833),
.B(n_9965),
.Y(n_21053)
);

AOI22xp5_ASAP7_75t_L g21054 ( 
.A1(n_20938),
.A2(n_11094),
.B1(n_11089),
.B2(n_10296),
.Y(n_21054)
);

NAND3xp33_ASAP7_75t_SL g21055 ( 
.A(n_20884),
.B(n_20973),
.C(n_20901),
.Y(n_21055)
);

NAND2xp5_ASAP7_75t_L g21056 ( 
.A(n_20847),
.B(n_9965),
.Y(n_21056)
);

NOR2x1_ASAP7_75t_L g21057 ( 
.A(n_20890),
.B(n_9863),
.Y(n_21057)
);

INVx1_ASAP7_75t_L g21058 ( 
.A(n_20963),
.Y(n_21058)
);

NAND4xp25_ASAP7_75t_L g21059 ( 
.A(n_20910),
.B(n_8826),
.C(n_9047),
.D(n_8997),
.Y(n_21059)
);

NOR2xp67_ASAP7_75t_L g21060 ( 
.A(n_20921),
.B(n_8749),
.Y(n_21060)
);

NOR2x1_ASAP7_75t_L g21061 ( 
.A(n_20931),
.B(n_9863),
.Y(n_21061)
);

INVx1_ASAP7_75t_L g21062 ( 
.A(n_20953),
.Y(n_21062)
);

INVx1_ASAP7_75t_L g21063 ( 
.A(n_20922),
.Y(n_21063)
);

AND2x2_ASAP7_75t_L g21064 ( 
.A(n_20970),
.B(n_9624),
.Y(n_21064)
);

NOR2xp33_ASAP7_75t_L g21065 ( 
.A(n_20958),
.B(n_20924),
.Y(n_21065)
);

NAND3xp33_ASAP7_75t_L g21066 ( 
.A(n_20864),
.B(n_9925),
.C(n_10288),
.Y(n_21066)
);

NAND2xp5_ASAP7_75t_L g21067 ( 
.A(n_20883),
.B(n_9965),
.Y(n_21067)
);

INVx1_ASAP7_75t_L g21068 ( 
.A(n_20793),
.Y(n_21068)
);

NOR2xp33_ASAP7_75t_L g21069 ( 
.A(n_20939),
.B(n_9925),
.Y(n_21069)
);

INVx2_ASAP7_75t_L g21070 ( 
.A(n_20961),
.Y(n_21070)
);

NOR2xp33_ASAP7_75t_SL g21071 ( 
.A(n_20962),
.B(n_20875),
.Y(n_21071)
);

OAI211xp5_ASAP7_75t_L g21072 ( 
.A1(n_20812),
.A2(n_10206),
.B(n_10225),
.C(n_10202),
.Y(n_21072)
);

INVx1_ASAP7_75t_L g21073 ( 
.A(n_20959),
.Y(n_21073)
);

AND2x2_ASAP7_75t_L g21074 ( 
.A(n_20794),
.B(n_20894),
.Y(n_21074)
);

NOR4xp25_ASAP7_75t_L g21075 ( 
.A(n_20952),
.B(n_9133),
.C(n_9147),
.D(n_9132),
.Y(n_21075)
);

NAND2xp5_ASAP7_75t_L g21076 ( 
.A(n_20862),
.B(n_9965),
.Y(n_21076)
);

OR2x2_ASAP7_75t_L g21077 ( 
.A(n_20846),
.B(n_10255),
.Y(n_21077)
);

AOI22xp33_ASAP7_75t_L g21078 ( 
.A1(n_20945),
.A2(n_20839),
.B1(n_20792),
.B2(n_20824),
.Y(n_21078)
);

NAND2x1_ASAP7_75t_SL g21079 ( 
.A(n_20840),
.B(n_20832),
.Y(n_21079)
);

NAND3xp33_ASAP7_75t_L g21080 ( 
.A(n_20966),
.B(n_10296),
.C(n_10288),
.Y(n_21080)
);

INVx2_ASAP7_75t_L g21081 ( 
.A(n_20900),
.Y(n_21081)
);

NAND2xp5_ASAP7_75t_L g21082 ( 
.A(n_20801),
.B(n_11089),
.Y(n_21082)
);

OAI21xp5_ASAP7_75t_SL g21083 ( 
.A1(n_20957),
.A2(n_9535),
.B(n_9464),
.Y(n_21083)
);

INVx1_ASAP7_75t_L g21084 ( 
.A(n_20848),
.Y(n_21084)
);

NOR2xp33_ASAP7_75t_L g21085 ( 
.A(n_20855),
.B(n_11089),
.Y(n_21085)
);

NAND2xp5_ASAP7_75t_L g21086 ( 
.A(n_20893),
.B(n_20802),
.Y(n_21086)
);

AND2x2_ASAP7_75t_L g21087 ( 
.A(n_20984),
.B(n_9624),
.Y(n_21087)
);

NAND2xp5_ASAP7_75t_L g21088 ( 
.A(n_20870),
.B(n_11094),
.Y(n_21088)
);

INVx1_ASAP7_75t_L g21089 ( 
.A(n_20785),
.Y(n_21089)
);

NAND3x1_ASAP7_75t_SL g21090 ( 
.A(n_20863),
.B(n_8353),
.C(n_9813),
.Y(n_21090)
);

NAND2xp5_ASAP7_75t_L g21091 ( 
.A(n_20928),
.B(n_20872),
.Y(n_21091)
);

INVx1_ASAP7_75t_L g21092 ( 
.A(n_20981),
.Y(n_21092)
);

NAND2xp5_ASAP7_75t_L g21093 ( 
.A(n_20796),
.B(n_11094),
.Y(n_21093)
);

AOI21xp5_ASAP7_75t_L g21094 ( 
.A1(n_20926),
.A2(n_20866),
.B(n_20897),
.Y(n_21094)
);

INVx1_ASAP7_75t_L g21095 ( 
.A(n_20896),
.Y(n_21095)
);

NAND2xp5_ASAP7_75t_SL g21096 ( 
.A(n_20940),
.B(n_8248),
.Y(n_21096)
);

INVx1_ASAP7_75t_L g21097 ( 
.A(n_20813),
.Y(n_21097)
);

NAND2xp5_ASAP7_75t_SL g21098 ( 
.A(n_20923),
.B(n_8248),
.Y(n_21098)
);

OAI21xp33_ASAP7_75t_SL g21099 ( 
.A1(n_20829),
.A2(n_10533),
.B(n_10532),
.Y(n_21099)
);

NOR2xp33_ASAP7_75t_L g21100 ( 
.A(n_20828),
.B(n_11094),
.Y(n_21100)
);

AND2x2_ASAP7_75t_L g21101 ( 
.A(n_20886),
.B(n_9624),
.Y(n_21101)
);

A2O1A1Ixp33_ASAP7_75t_L g21102 ( 
.A1(n_20965),
.A2(n_10964),
.B(n_10968),
.C(n_10967),
.Y(n_21102)
);

INVx1_ASAP7_75t_L g21103 ( 
.A(n_20791),
.Y(n_21103)
);

NAND3xp33_ASAP7_75t_L g21104 ( 
.A(n_20887),
.B(n_10296),
.C(n_10288),
.Y(n_21104)
);

NAND4xp25_ASAP7_75t_L g21105 ( 
.A(n_20799),
.B(n_8826),
.C(n_9047),
.D(n_8997),
.Y(n_21105)
);

AOI211x1_ASAP7_75t_SL g21106 ( 
.A1(n_20933),
.A2(n_9071),
.B(n_9107),
.C(n_9042),
.Y(n_21106)
);

NAND3xp33_ASAP7_75t_L g21107 ( 
.A(n_20854),
.B(n_10296),
.C(n_10288),
.Y(n_21107)
);

NAND2xp5_ASAP7_75t_SL g21108 ( 
.A(n_20852),
.B(n_8248),
.Y(n_21108)
);

INVx1_ASAP7_75t_L g21109 ( 
.A(n_20861),
.Y(n_21109)
);

INVx1_ASAP7_75t_L g21110 ( 
.A(n_20903),
.Y(n_21110)
);

AOI221xp5_ASAP7_75t_L g21111 ( 
.A1(n_20909),
.A2(n_9520),
.B1(n_9510),
.B2(n_9147),
.C(n_9162),
.Y(n_21111)
);

NAND2xp5_ASAP7_75t_L g21112 ( 
.A(n_20821),
.B(n_10255),
.Y(n_21112)
);

NOR2xp33_ASAP7_75t_L g21113 ( 
.A(n_20808),
.B(n_7706),
.Y(n_21113)
);

NAND3xp33_ASAP7_75t_L g21114 ( 
.A(n_20835),
.B(n_10302),
.C(n_10288),
.Y(n_21114)
);

NOR2xp33_ASAP7_75t_L g21115 ( 
.A(n_20899),
.B(n_7706),
.Y(n_21115)
);

NOR3xp33_ASAP7_75t_L g21116 ( 
.A(n_20950),
.B(n_10824),
.C(n_10823),
.Y(n_21116)
);

NAND3xp33_ASAP7_75t_SL g21117 ( 
.A(n_20805),
.B(n_9540),
.C(n_9535),
.Y(n_21117)
);

NAND2xp33_ASAP7_75t_SL g21118 ( 
.A(n_20898),
.B(n_20850),
.Y(n_21118)
);

NOR4xp25_ASAP7_75t_SL g21119 ( 
.A(n_20826),
.B(n_8835),
.C(n_10035),
.D(n_10030),
.Y(n_21119)
);

NAND2xp5_ASAP7_75t_L g21120 ( 
.A(n_20822),
.B(n_10255),
.Y(n_21120)
);

NAND2xp5_ASAP7_75t_SL g21121 ( 
.A(n_20806),
.B(n_8248),
.Y(n_21121)
);

OAI32xp33_ASAP7_75t_L g21122 ( 
.A1(n_20844),
.A2(n_9071),
.A3(n_9120),
.B1(n_9114),
.B2(n_9107),
.Y(n_21122)
);

AND2x4_ASAP7_75t_L g21123 ( 
.A(n_20968),
.B(n_9520),
.Y(n_21123)
);

NAND2xp5_ASAP7_75t_L g21124 ( 
.A(n_20954),
.B(n_20908),
.Y(n_21124)
);

INVx1_ASAP7_75t_L g21125 ( 
.A(n_20789),
.Y(n_21125)
);

NOR4xp75_ASAP7_75t_L g21126 ( 
.A(n_20956),
.B(n_9804),
.C(n_9807),
.D(n_9803),
.Y(n_21126)
);

NAND4xp25_ASAP7_75t_L g21127 ( 
.A(n_20841),
.B(n_9047),
.C(n_9048),
.D(n_8997),
.Y(n_21127)
);

INVx1_ASAP7_75t_SL g21128 ( 
.A(n_20955),
.Y(n_21128)
);

NAND2xp5_ASAP7_75t_L g21129 ( 
.A(n_20820),
.B(n_10255),
.Y(n_21129)
);

INVx1_ASAP7_75t_L g21130 ( 
.A(n_20800),
.Y(n_21130)
);

INVxp67_ASAP7_75t_L g21131 ( 
.A(n_20804),
.Y(n_21131)
);

NAND4xp25_ASAP7_75t_L g21132 ( 
.A(n_20797),
.B(n_9047),
.C(n_9048),
.D(n_8997),
.Y(n_21132)
);

INVx1_ASAP7_75t_L g21133 ( 
.A(n_20955),
.Y(n_21133)
);

NAND2xp5_ASAP7_75t_L g21134 ( 
.A(n_20816),
.B(n_10255),
.Y(n_21134)
);

NOR2xp67_ASAP7_75t_L g21135 ( 
.A(n_20972),
.B(n_8749),
.Y(n_21135)
);

INVx1_ASAP7_75t_SL g21136 ( 
.A(n_20947),
.Y(n_21136)
);

OAI211xp5_ASAP7_75t_L g21137 ( 
.A1(n_20856),
.A2(n_10230),
.B(n_10248),
.C(n_10202),
.Y(n_21137)
);

INVx2_ASAP7_75t_L g21138 ( 
.A(n_20964),
.Y(n_21138)
);

NOR3xp33_ASAP7_75t_L g21139 ( 
.A(n_20815),
.B(n_10830),
.C(n_11425),
.Y(n_21139)
);

NAND4xp25_ASAP7_75t_L g21140 ( 
.A(n_20911),
.B(n_9047),
.C(n_9048),
.D(n_8997),
.Y(n_21140)
);

INVx1_ASAP7_75t_L g21141 ( 
.A(n_20895),
.Y(n_21141)
);

AOI21xp5_ASAP7_75t_L g21142 ( 
.A1(n_20943),
.A2(n_10691),
.B(n_10320),
.Y(n_21142)
);

CKINVDCx5p33_ASAP7_75t_R g21143 ( 
.A(n_20879),
.Y(n_21143)
);

NAND2xp5_ASAP7_75t_L g21144 ( 
.A(n_20860),
.B(n_10255),
.Y(n_21144)
);

INVxp67_ASAP7_75t_SL g21145 ( 
.A(n_20834),
.Y(n_21145)
);

INVx2_ASAP7_75t_L g21146 ( 
.A(n_20905),
.Y(n_21146)
);

NAND2xp5_ASAP7_75t_L g21147 ( 
.A(n_20784),
.B(n_10255),
.Y(n_21147)
);

INVx1_ASAP7_75t_L g21148 ( 
.A(n_20998),
.Y(n_21148)
);

NOR4xp25_ASAP7_75t_L g21149 ( 
.A(n_21000),
.B(n_20809),
.C(n_20849),
.D(n_20927),
.Y(n_21149)
);

NAND2xp5_ASAP7_75t_SL g21150 ( 
.A(n_21009),
.B(n_20871),
.Y(n_21150)
);

NOR2xp33_ASAP7_75t_L g21151 ( 
.A(n_21002),
.B(n_20837),
.Y(n_21151)
);

NAND2xp5_ASAP7_75t_L g21152 ( 
.A(n_20990),
.B(n_20795),
.Y(n_21152)
);

NAND3xp33_ASAP7_75t_L g21153 ( 
.A(n_21017),
.B(n_20917),
.C(n_20951),
.Y(n_21153)
);

NOR3xp33_ASAP7_75t_L g21154 ( 
.A(n_20985),
.B(n_20853),
.C(n_20918),
.Y(n_21154)
);

NOR3xp33_ASAP7_75t_L g21155 ( 
.A(n_21019),
.B(n_20936),
.C(n_20876),
.Y(n_21155)
);

OAI211xp5_ASAP7_75t_SL g21156 ( 
.A1(n_20999),
.A2(n_20935),
.B(n_20907),
.C(n_20919),
.Y(n_21156)
);

NOR2xp33_ASAP7_75t_L g21157 ( 
.A(n_21030),
.B(n_20831),
.Y(n_21157)
);

NAND3xp33_ASAP7_75t_L g21158 ( 
.A(n_21065),
.B(n_20823),
.C(n_20891),
.Y(n_21158)
);

NAND3xp33_ASAP7_75t_L g21159 ( 
.A(n_21014),
.B(n_20948),
.C(n_10248),
.Y(n_21159)
);

O2A1O1Ixp5_ASAP7_75t_SL g21160 ( 
.A1(n_21001),
.A2(n_9133),
.B(n_9162),
.C(n_9155),
.Y(n_21160)
);

NAND3xp33_ASAP7_75t_SL g21161 ( 
.A(n_21128),
.B(n_21143),
.C(n_21027),
.Y(n_21161)
);

NOR4xp25_ASAP7_75t_L g21162 ( 
.A(n_21103),
.B(n_10035),
.C(n_10046),
.D(n_10030),
.Y(n_21162)
);

NAND3xp33_ASAP7_75t_L g21163 ( 
.A(n_21130),
.B(n_10248),
.C(n_10230),
.Y(n_21163)
);

NAND2xp5_ASAP7_75t_SL g21164 ( 
.A(n_20987),
.B(n_8248),
.Y(n_21164)
);

AND2x2_ASAP7_75t_L g21165 ( 
.A(n_21049),
.B(n_9624),
.Y(n_21165)
);

AOI21xp5_ASAP7_75t_L g21166 ( 
.A1(n_21091),
.A2(n_10691),
.B(n_10548),
.Y(n_21166)
);

OAI21xp33_ASAP7_75t_L g21167 ( 
.A1(n_21071),
.A2(n_9162),
.B(n_9155),
.Y(n_21167)
);

NOR3xp33_ASAP7_75t_L g21168 ( 
.A(n_21058),
.B(n_10830),
.C(n_10580),
.Y(n_21168)
);

NAND4xp25_ASAP7_75t_L g21169 ( 
.A(n_20993),
.B(n_7731),
.C(n_7745),
.D(n_7738),
.Y(n_21169)
);

NOR3xp33_ASAP7_75t_L g21170 ( 
.A(n_20988),
.B(n_10830),
.C(n_10580),
.Y(n_21170)
);

OAI21xp5_ASAP7_75t_L g21171 ( 
.A1(n_21131),
.A2(n_21004),
.B(n_21018),
.Y(n_21171)
);

OAI211xp5_ASAP7_75t_L g21172 ( 
.A1(n_21145),
.A2(n_10248),
.B(n_10267),
.C(n_10230),
.Y(n_21172)
);

OR2x2_ASAP7_75t_L g21173 ( 
.A(n_21010),
.B(n_10255),
.Y(n_21173)
);

AOI221xp5_ASAP7_75t_L g21174 ( 
.A1(n_21118),
.A2(n_9165),
.B1(n_9173),
.B2(n_9162),
.C(n_9155),
.Y(n_21174)
);

NAND4xp75_ASAP7_75t_L g21175 ( 
.A(n_21062),
.B(n_10248),
.C(n_10267),
.D(n_10230),
.Y(n_21175)
);

NOR3xp33_ASAP7_75t_L g21176 ( 
.A(n_21029),
.B(n_11426),
.C(n_11425),
.Y(n_21176)
);

NOR3xp33_ASAP7_75t_L g21177 ( 
.A(n_21015),
.B(n_11438),
.C(n_11426),
.Y(n_21177)
);

OAI211xp5_ASAP7_75t_L g21178 ( 
.A1(n_21141),
.A2(n_10248),
.B(n_10267),
.C(n_10230),
.Y(n_21178)
);

HB1xp67_ASAP7_75t_L g21179 ( 
.A(n_21133),
.Y(n_21179)
);

NAND4xp25_ASAP7_75t_L g21180 ( 
.A(n_21013),
.B(n_7738),
.C(n_7745),
.D(n_7724),
.Y(n_21180)
);

NAND4xp25_ASAP7_75t_L g21181 ( 
.A(n_21136),
.B(n_21089),
.C(n_21125),
.D(n_21074),
.Y(n_21181)
);

NAND4xp25_ASAP7_75t_L g21182 ( 
.A(n_21092),
.B(n_9047),
.C(n_9048),
.D(n_8997),
.Y(n_21182)
);

INVx1_ASAP7_75t_L g21183 ( 
.A(n_21070),
.Y(n_21183)
);

NAND3xp33_ASAP7_75t_L g21184 ( 
.A(n_21146),
.B(n_10267),
.C(n_10230),
.Y(n_21184)
);

NOR4xp25_ASAP7_75t_L g21185 ( 
.A(n_21110),
.B(n_10046),
.C(n_10050),
.D(n_10035),
.Y(n_21185)
);

OAI211xp5_ASAP7_75t_L g21186 ( 
.A1(n_21095),
.A2(n_21073),
.B(n_21051),
.C(n_21063),
.Y(n_21186)
);

NAND2xp5_ASAP7_75t_L g21187 ( 
.A(n_21078),
.B(n_9909),
.Y(n_21187)
);

AND4x1_ASAP7_75t_L g21188 ( 
.A(n_21042),
.B(n_9813),
.C(n_9852),
.D(n_8353),
.Y(n_21188)
);

NOR3xp33_ASAP7_75t_L g21189 ( 
.A(n_21035),
.B(n_11439),
.C(n_11438),
.Y(n_21189)
);

NOR3xp33_ASAP7_75t_L g21190 ( 
.A(n_21033),
.B(n_11439),
.C(n_11438),
.Y(n_21190)
);

NAND3xp33_ASAP7_75t_L g21191 ( 
.A(n_21044),
.B(n_10267),
.C(n_10288),
.Y(n_21191)
);

NAND4xp75_ASAP7_75t_L g21192 ( 
.A(n_21068),
.B(n_10267),
.C(n_11335),
.D(n_10302),
.Y(n_21192)
);

NAND3xp33_ASAP7_75t_L g21193 ( 
.A(n_21084),
.B(n_10302),
.C(n_11335),
.Y(n_21193)
);

NOR2xp67_ASAP7_75t_L g21194 ( 
.A(n_21138),
.B(n_8749),
.Y(n_21194)
);

OAI31xp33_ASAP7_75t_L g21195 ( 
.A1(n_21081),
.A2(n_9540),
.A3(n_9643),
.B(n_9535),
.Y(n_21195)
);

AOI321xp33_ASAP7_75t_L g21196 ( 
.A1(n_21094),
.A2(n_9048),
.A3(n_8997),
.B1(n_9109),
.B2(n_9089),
.C(n_9047),
.Y(n_21196)
);

NAND4xp25_ASAP7_75t_L g21197 ( 
.A(n_21055),
.B(n_9089),
.C(n_9048),
.D(n_9047),
.Y(n_21197)
);

NOR2x1_ASAP7_75t_L g21198 ( 
.A(n_21109),
.B(n_9863),
.Y(n_21198)
);

NAND4xp25_ASAP7_75t_L g21199 ( 
.A(n_21086),
.B(n_21124),
.C(n_21097),
.D(n_21135),
.Y(n_21199)
);

NOR3xp33_ASAP7_75t_L g21200 ( 
.A(n_20996),
.B(n_11449),
.C(n_11448),
.Y(n_21200)
);

NOR3xp33_ASAP7_75t_L g21201 ( 
.A(n_21053),
.B(n_11449),
.C(n_11448),
.Y(n_21201)
);

NOR3xp33_ASAP7_75t_L g21202 ( 
.A(n_21037),
.B(n_11449),
.C(n_11448),
.Y(n_21202)
);

NAND4xp25_ASAP7_75t_L g21203 ( 
.A(n_21006),
.B(n_21025),
.C(n_21085),
.D(n_21105),
.Y(n_21203)
);

OAI211xp5_ASAP7_75t_SL g21204 ( 
.A1(n_21108),
.A2(n_10050),
.B(n_10057),
.C(n_10046),
.Y(n_21204)
);

AOI211xp5_ASAP7_75t_SL g21205 ( 
.A1(n_21067),
.A2(n_21045),
.B(n_21147),
.C(n_21076),
.Y(n_21205)
);

NAND5xp2_ASAP7_75t_L g21206 ( 
.A(n_21083),
.B(n_9643),
.C(n_9709),
.D(n_9644),
.E(n_9540),
.Y(n_21206)
);

NAND2xp5_ASAP7_75t_L g21207 ( 
.A(n_21079),
.B(n_9909),
.Y(n_21207)
);

INVx2_ASAP7_75t_L g21208 ( 
.A(n_21077),
.Y(n_21208)
);

NOR3xp33_ASAP7_75t_L g21209 ( 
.A(n_21121),
.B(n_11467),
.C(n_11439),
.Y(n_21209)
);

AOI211xp5_ASAP7_75t_L g21210 ( 
.A1(n_21122),
.A2(n_21026),
.B(n_21060),
.C(n_21115),
.Y(n_21210)
);

NOR2xp33_ASAP7_75t_L g21211 ( 
.A(n_21132),
.B(n_11335),
.Y(n_21211)
);

OR3x1_ASAP7_75t_L g21212 ( 
.A(n_20986),
.B(n_10057),
.C(n_10050),
.Y(n_21212)
);

NAND2xp5_ASAP7_75t_L g21213 ( 
.A(n_21012),
.B(n_9909),
.Y(n_21213)
);

NAND2xp5_ASAP7_75t_L g21214 ( 
.A(n_21123),
.B(n_21057),
.Y(n_21214)
);

NOR2x1_ASAP7_75t_L g21215 ( 
.A(n_21061),
.B(n_9863),
.Y(n_21215)
);

AOI21xp5_ASAP7_75t_L g21216 ( 
.A1(n_21003),
.A2(n_10691),
.B(n_10548),
.Y(n_21216)
);

NAND2xp5_ASAP7_75t_SL g21217 ( 
.A(n_21023),
.B(n_8248),
.Y(n_21217)
);

AOI221xp5_ASAP7_75t_L g21218 ( 
.A1(n_21075),
.A2(n_9176),
.B1(n_9193),
.B2(n_9173),
.C(n_9165),
.Y(n_21218)
);

AOI211x1_ASAP7_75t_L g21219 ( 
.A1(n_21098),
.A2(n_9173),
.B(n_9176),
.C(n_9165),
.Y(n_21219)
);

NAND3xp33_ASAP7_75t_L g21220 ( 
.A(n_21050),
.B(n_10302),
.C(n_11335),
.Y(n_21220)
);

AOI311xp33_ASAP7_75t_L g21221 ( 
.A1(n_21116),
.A2(n_9176),
.A3(n_9193),
.B(n_9173),
.C(n_9165),
.Y(n_21221)
);

NAND2xp5_ASAP7_75t_SL g21222 ( 
.A(n_21123),
.B(n_8248),
.Y(n_21222)
);

NAND2xp5_ASAP7_75t_L g21223 ( 
.A(n_21038),
.B(n_9909),
.Y(n_21223)
);

NOR2xp67_ASAP7_75t_L g21224 ( 
.A(n_21066),
.B(n_8749),
.Y(n_21224)
);

NOR3xp33_ASAP7_75t_L g21225 ( 
.A(n_21090),
.B(n_11479),
.C(n_11467),
.Y(n_21225)
);

OAI21xp33_ASAP7_75t_L g21226 ( 
.A1(n_21144),
.A2(n_9193),
.B(n_9176),
.Y(n_21226)
);

NAND2xp5_ASAP7_75t_L g21227 ( 
.A(n_21032),
.B(n_9909),
.Y(n_21227)
);

NOR4xp75_ASAP7_75t_L g21228 ( 
.A(n_21005),
.B(n_9807),
.C(n_9804),
.D(n_9803),
.Y(n_21228)
);

OAI211xp5_ASAP7_75t_SL g21229 ( 
.A1(n_21056),
.A2(n_10057),
.B(n_10064),
.C(n_10050),
.Y(n_21229)
);

NAND3xp33_ASAP7_75t_SL g21230 ( 
.A(n_21111),
.B(n_9644),
.C(n_9643),
.Y(n_21230)
);

INVx1_ASAP7_75t_L g21231 ( 
.A(n_21112),
.Y(n_21231)
);

NOR3x1_ASAP7_75t_L g21232 ( 
.A(n_21117),
.B(n_10967),
.C(n_10964),
.Y(n_21232)
);

NAND2xp5_ASAP7_75t_L g21233 ( 
.A(n_21113),
.B(n_9909),
.Y(n_21233)
);

O2A1O1Ixp33_ASAP7_75t_L g21234 ( 
.A1(n_21096),
.A2(n_9239),
.B(n_9709),
.C(n_9644),
.Y(n_21234)
);

NAND2xp5_ASAP7_75t_SL g21235 ( 
.A(n_20991),
.B(n_8273),
.Y(n_21235)
);

AOI211x1_ASAP7_75t_L g21236 ( 
.A1(n_21052),
.A2(n_9194),
.B(n_9197),
.C(n_9193),
.Y(n_21236)
);

NAND3xp33_ASAP7_75t_L g21237 ( 
.A(n_21139),
.B(n_10302),
.C(n_11335),
.Y(n_21237)
);

OR2x2_ASAP7_75t_L g21238 ( 
.A(n_21127),
.B(n_11535),
.Y(n_21238)
);

OAI222xp33_ASAP7_75t_R g21239 ( 
.A1(n_21040),
.A2(n_8513),
.B1(n_8284),
.B2(n_8202),
.C1(n_8322),
.C2(n_8212),
.Y(n_21239)
);

A2O1A1Ixp33_ASAP7_75t_L g21240 ( 
.A1(n_21100),
.A2(n_10967),
.B(n_10969),
.C(n_10968),
.Y(n_21240)
);

NOR2x1_ASAP7_75t_L g21241 ( 
.A(n_21120),
.B(n_9863),
.Y(n_21241)
);

AOI211xp5_ASAP7_75t_L g21242 ( 
.A1(n_21129),
.A2(n_10276),
.B(n_10279),
.C(n_10256),
.Y(n_21242)
);

OAI21xp33_ASAP7_75t_L g21243 ( 
.A1(n_21007),
.A2(n_9197),
.B(n_9194),
.Y(n_21243)
);

NAND2xp5_ASAP7_75t_L g21244 ( 
.A(n_21134),
.B(n_9909),
.Y(n_21244)
);

AOI221xp5_ASAP7_75t_L g21245 ( 
.A1(n_21031),
.A2(n_9207),
.B1(n_9215),
.B2(n_9197),
.C(n_9194),
.Y(n_21245)
);

OAI21xp33_ASAP7_75t_L g21246 ( 
.A1(n_21140),
.A2(n_9197),
.B(n_9194),
.Y(n_21246)
);

OAI222xp33_ASAP7_75t_R g21247 ( 
.A1(n_21054),
.A2(n_8284),
.B1(n_8202),
.B2(n_8322),
.C1(n_8212),
.C2(n_8623),
.Y(n_21247)
);

NAND2xp5_ASAP7_75t_L g21248 ( 
.A(n_21046),
.B(n_9909),
.Y(n_21248)
);

NOR2x1_ASAP7_75t_L g21249 ( 
.A(n_21008),
.B(n_9863),
.Y(n_21249)
);

INVx1_ASAP7_75t_L g21250 ( 
.A(n_21088),
.Y(n_21250)
);

O2A1O1Ixp33_ASAP7_75t_L g21251 ( 
.A1(n_21093),
.A2(n_9239),
.B(n_9709),
.C(n_9644),
.Y(n_21251)
);

O2A1O1Ixp33_ASAP7_75t_L g21252 ( 
.A1(n_21082),
.A2(n_9239),
.B(n_9709),
.C(n_9644),
.Y(n_21252)
);

NAND3xp33_ASAP7_75t_L g21253 ( 
.A(n_21080),
.B(n_10302),
.C(n_11335),
.Y(n_21253)
);

OAI211xp5_ASAP7_75t_L g21254 ( 
.A1(n_21011),
.A2(n_9215),
.B(n_9216),
.C(n_9207),
.Y(n_21254)
);

NAND3xp33_ASAP7_75t_L g21255 ( 
.A(n_21041),
.B(n_9909),
.C(n_9309),
.Y(n_21255)
);

AOI211xp5_ASAP7_75t_L g21256 ( 
.A1(n_21043),
.A2(n_10276),
.B(n_10279),
.C(n_10256),
.Y(n_21256)
);

NAND4xp75_ASAP7_75t_L g21257 ( 
.A(n_21064),
.B(n_11114),
.C(n_11146),
.D(n_11108),
.Y(n_21257)
);

NOR3xp33_ASAP7_75t_L g21258 ( 
.A(n_20992),
.B(n_11479),
.C(n_11467),
.Y(n_21258)
);

AOI21xp5_ASAP7_75t_L g21259 ( 
.A1(n_20997),
.A2(n_21028),
.B(n_21020),
.Y(n_21259)
);

INVx1_ASAP7_75t_L g21260 ( 
.A(n_21106),
.Y(n_21260)
);

NAND3xp33_ASAP7_75t_L g21261 ( 
.A(n_20989),
.B(n_9309),
.C(n_9276),
.Y(n_21261)
);

AO221x1_ASAP7_75t_L g21262 ( 
.A1(n_21119),
.A2(n_8314),
.B1(n_8349),
.B2(n_8296),
.C(n_8273),
.Y(n_21262)
);

INVx1_ASAP7_75t_L g21263 ( 
.A(n_21087),
.Y(n_21263)
);

NAND3xp33_ASAP7_75t_SL g21264 ( 
.A(n_21047),
.B(n_9709),
.C(n_9644),
.Y(n_21264)
);

AOI211xp5_ASAP7_75t_L g21265 ( 
.A1(n_21059),
.A2(n_10279),
.B(n_11483),
.C(n_11479),
.Y(n_21265)
);

NOR4xp25_ASAP7_75t_L g21266 ( 
.A(n_21137),
.B(n_10064),
.C(n_10069),
.D(n_10057),
.Y(n_21266)
);

NOR4xp25_ASAP7_75t_L g21267 ( 
.A(n_21072),
.B(n_21102),
.C(n_21114),
.D(n_20995),
.Y(n_21267)
);

NAND4xp25_ASAP7_75t_L g21268 ( 
.A(n_21039),
.B(n_9047),
.C(n_9048),
.D(n_8997),
.Y(n_21268)
);

NOR2xp33_ASAP7_75t_L g21269 ( 
.A(n_21101),
.B(n_7860),
.Y(n_21269)
);

AOI311xp33_ASAP7_75t_L g21270 ( 
.A1(n_21069),
.A2(n_9216),
.A3(n_9221),
.B(n_9215),
.C(n_9207),
.Y(n_21270)
);

NAND3xp33_ASAP7_75t_L g21271 ( 
.A(n_21034),
.B(n_21022),
.C(n_21016),
.Y(n_21271)
);

AND2x2_ASAP7_75t_L g21272 ( 
.A(n_21036),
.B(n_9624),
.Y(n_21272)
);

NAND5xp2_ASAP7_75t_L g21273 ( 
.A(n_21021),
.B(n_9712),
.C(n_9834),
.D(n_9819),
.E(n_9709),
.Y(n_21273)
);

NAND2xp5_ASAP7_75t_SL g21274 ( 
.A(n_21099),
.B(n_8273),
.Y(n_21274)
);

NAND2xp5_ASAP7_75t_L g21275 ( 
.A(n_21142),
.B(n_9024),
.Y(n_21275)
);

AOI221xp5_ASAP7_75t_L g21276 ( 
.A1(n_21107),
.A2(n_21104),
.B1(n_21048),
.B2(n_21126),
.C(n_20994),
.Y(n_21276)
);

NOR4xp25_ASAP7_75t_L g21277 ( 
.A(n_21024),
.B(n_10069),
.C(n_10075),
.D(n_10064),
.Y(n_21277)
);

INVxp67_ASAP7_75t_L g21278 ( 
.A(n_20987),
.Y(n_21278)
);

NAND4xp25_ASAP7_75t_SL g21279 ( 
.A(n_21000),
.B(n_9215),
.C(n_9216),
.D(n_9207),
.Y(n_21279)
);

NAND2xp5_ASAP7_75t_SL g21280 ( 
.A(n_21000),
.B(n_8273),
.Y(n_21280)
);

AOI211xp5_ASAP7_75t_L g21281 ( 
.A1(n_20988),
.A2(n_11493),
.B(n_11505),
.C(n_11483),
.Y(n_21281)
);

INVx1_ASAP7_75t_L g21282 ( 
.A(n_20998),
.Y(n_21282)
);

NAND4xp25_ASAP7_75t_L g21283 ( 
.A(n_21071),
.B(n_9089),
.C(n_9109),
.D(n_9048),
.Y(n_21283)
);

AOI21xp33_ASAP7_75t_L g21284 ( 
.A1(n_21000),
.A2(n_9679),
.B(n_10316),
.Y(n_21284)
);

NAND2xp5_ASAP7_75t_SL g21285 ( 
.A(n_21000),
.B(n_8273),
.Y(n_21285)
);

AND2x2_ASAP7_75t_L g21286 ( 
.A(n_20987),
.B(n_9633),
.Y(n_21286)
);

AOI221x1_ASAP7_75t_L g21287 ( 
.A1(n_21000),
.A2(n_10075),
.B1(n_10085),
.B2(n_10069),
.C(n_10064),
.Y(n_21287)
);

NOR5xp2_ASAP7_75t_L g21288 ( 
.A(n_20999),
.B(n_7857),
.C(n_7997),
.D(n_7825),
.E(n_7732),
.Y(n_21288)
);

NAND2xp5_ASAP7_75t_L g21289 ( 
.A(n_20998),
.B(n_9024),
.Y(n_21289)
);

AOI211xp5_ASAP7_75t_L g21290 ( 
.A1(n_20988),
.A2(n_11493),
.B(n_11505),
.C(n_11483),
.Y(n_21290)
);

NOR3xp33_ASAP7_75t_SL g21291 ( 
.A(n_21143),
.B(n_10075),
.C(n_10069),
.Y(n_21291)
);

NAND4xp25_ASAP7_75t_L g21292 ( 
.A(n_21071),
.B(n_9089),
.C(n_9109),
.D(n_9048),
.Y(n_21292)
);

NAND3xp33_ASAP7_75t_SL g21293 ( 
.A(n_21128),
.B(n_9712),
.C(n_9709),
.Y(n_21293)
);

NAND3xp33_ASAP7_75t_SL g21294 ( 
.A(n_21128),
.B(n_9819),
.C(n_9712),
.Y(n_21294)
);

NAND3xp33_ASAP7_75t_SL g21295 ( 
.A(n_21128),
.B(n_9819),
.C(n_9712),
.Y(n_21295)
);

NOR3xp33_ASAP7_75t_L g21296 ( 
.A(n_21000),
.B(n_11508),
.C(n_11505),
.Y(n_21296)
);

NOR3xp33_ASAP7_75t_L g21297 ( 
.A(n_21000),
.B(n_11511),
.C(n_11508),
.Y(n_21297)
);

O2A1O1Ixp33_ASAP7_75t_L g21298 ( 
.A1(n_21000),
.A2(n_9239),
.B(n_9819),
.C(n_9712),
.Y(n_21298)
);

INVxp67_ASAP7_75t_L g21299 ( 
.A(n_20987),
.Y(n_21299)
);

NAND2xp5_ASAP7_75t_L g21300 ( 
.A(n_20998),
.B(n_9024),
.Y(n_21300)
);

INVx1_ASAP7_75t_L g21301 ( 
.A(n_21179),
.Y(n_21301)
);

INVx2_ASAP7_75t_L g21302 ( 
.A(n_21183),
.Y(n_21302)
);

INVx1_ASAP7_75t_L g21303 ( 
.A(n_21214),
.Y(n_21303)
);

AND2x2_ASAP7_75t_L g21304 ( 
.A(n_21278),
.B(n_10053),
.Y(n_21304)
);

NAND2xp5_ASAP7_75t_L g21305 ( 
.A(n_21299),
.B(n_10534),
.Y(n_21305)
);

NOR2xp33_ASAP7_75t_SL g21306 ( 
.A(n_21181),
.B(n_7782),
.Y(n_21306)
);

NAND2xp5_ASAP7_75t_SL g21307 ( 
.A(n_21149),
.B(n_9146),
.Y(n_21307)
);

INVxp67_ASAP7_75t_L g21308 ( 
.A(n_21151),
.Y(n_21308)
);

INVxp67_ASAP7_75t_L g21309 ( 
.A(n_21157),
.Y(n_21309)
);

INVx1_ASAP7_75t_L g21310 ( 
.A(n_21194),
.Y(n_21310)
);

INVx1_ASAP7_75t_L g21311 ( 
.A(n_21150),
.Y(n_21311)
);

BUFx2_ASAP7_75t_L g21312 ( 
.A(n_21148),
.Y(n_21312)
);

INVx1_ASAP7_75t_SL g21313 ( 
.A(n_21152),
.Y(n_21313)
);

NAND2xp33_ASAP7_75t_SL g21314 ( 
.A(n_21282),
.B(n_8796),
.Y(n_21314)
);

NOR2xp33_ASAP7_75t_L g21315 ( 
.A(n_21283),
.B(n_9900),
.Y(n_21315)
);

NAND2xp5_ASAP7_75t_L g21316 ( 
.A(n_21154),
.B(n_9679),
.Y(n_21316)
);

AOI21xp5_ASAP7_75t_L g21317 ( 
.A1(n_21161),
.A2(n_10322),
.B(n_10316),
.Y(n_21317)
);

INVx2_ASAP7_75t_L g21318 ( 
.A(n_21249),
.Y(n_21318)
);

XOR2x2_ASAP7_75t_L g21319 ( 
.A(n_21153),
.B(n_9712),
.Y(n_21319)
);

NOR2xp33_ASAP7_75t_L g21320 ( 
.A(n_21292),
.B(n_9900),
.Y(n_21320)
);

NAND2xp5_ASAP7_75t_L g21321 ( 
.A(n_21263),
.B(n_9679),
.Y(n_21321)
);

HB1xp67_ASAP7_75t_L g21322 ( 
.A(n_21208),
.Y(n_21322)
);

INVxp67_ASAP7_75t_SL g21323 ( 
.A(n_21155),
.Y(n_21323)
);

AND2x2_ASAP7_75t_L g21324 ( 
.A(n_21272),
.B(n_10053),
.Y(n_21324)
);

INVx1_ASAP7_75t_L g21325 ( 
.A(n_21271),
.Y(n_21325)
);

INVxp67_ASAP7_75t_L g21326 ( 
.A(n_21158),
.Y(n_21326)
);

OAI221xp5_ASAP7_75t_L g21327 ( 
.A1(n_21167),
.A2(n_9834),
.B1(n_9819),
.B2(n_9712),
.C(n_9900),
.Y(n_21327)
);

OAI221xp5_ASAP7_75t_L g21328 ( 
.A1(n_21276),
.A2(n_9834),
.B1(n_9819),
.B2(n_10002),
.C(n_9900),
.Y(n_21328)
);

NAND2xp5_ASAP7_75t_L g21329 ( 
.A(n_21260),
.B(n_9679),
.Y(n_21329)
);

INVx1_ASAP7_75t_L g21330 ( 
.A(n_21280),
.Y(n_21330)
);

BUFx6f_ASAP7_75t_L g21331 ( 
.A(n_21231),
.Y(n_21331)
);

NAND4xp25_ASAP7_75t_L g21332 ( 
.A(n_21203),
.B(n_9109),
.C(n_9113),
.D(n_9089),
.Y(n_21332)
);

AND2x2_ASAP7_75t_L g21333 ( 
.A(n_21171),
.B(n_10053),
.Y(n_21333)
);

INVx1_ASAP7_75t_L g21334 ( 
.A(n_21285),
.Y(n_21334)
);

NAND2xp5_ASAP7_75t_L g21335 ( 
.A(n_21210),
.B(n_9679),
.Y(n_21335)
);

INVx1_ASAP7_75t_L g21336 ( 
.A(n_21222),
.Y(n_21336)
);

INVx2_ASAP7_75t_SL g21337 ( 
.A(n_21241),
.Y(n_21337)
);

INVxp67_ASAP7_75t_L g21338 ( 
.A(n_21199),
.Y(n_21338)
);

INVx1_ASAP7_75t_L g21339 ( 
.A(n_21250),
.Y(n_21339)
);

NAND2xp5_ASAP7_75t_SL g21340 ( 
.A(n_21187),
.B(n_9146),
.Y(n_21340)
);

NAND2xp5_ASAP7_75t_L g21341 ( 
.A(n_21224),
.B(n_9679),
.Y(n_21341)
);

NAND2xp5_ASAP7_75t_SL g21342 ( 
.A(n_21267),
.B(n_9146),
.Y(n_21342)
);

INVx1_ASAP7_75t_L g21343 ( 
.A(n_21186),
.Y(n_21343)
);

NAND3xp33_ASAP7_75t_L g21344 ( 
.A(n_21205),
.B(n_9114),
.C(n_9107),
.Y(n_21344)
);

OAI221xp5_ASAP7_75t_L g21345 ( 
.A1(n_21207),
.A2(n_21159),
.B1(n_21156),
.B2(n_21226),
.C(n_21215),
.Y(n_21345)
);

INVxp67_ASAP7_75t_SL g21346 ( 
.A(n_21259),
.Y(n_21346)
);

INVx1_ASAP7_75t_L g21347 ( 
.A(n_21217),
.Y(n_21347)
);

INVx1_ASAP7_75t_L g21348 ( 
.A(n_21235),
.Y(n_21348)
);

NOR3xp33_ASAP7_75t_L g21349 ( 
.A(n_21268),
.B(n_10326),
.C(n_10322),
.Y(n_21349)
);

NAND2xp5_ASAP7_75t_L g21350 ( 
.A(n_21246),
.B(n_21164),
.Y(n_21350)
);

INVxp67_ASAP7_75t_L g21351 ( 
.A(n_21274),
.Y(n_21351)
);

INVx1_ASAP7_75t_L g21352 ( 
.A(n_21212),
.Y(n_21352)
);

NAND2xp5_ASAP7_75t_L g21353 ( 
.A(n_21291),
.B(n_9679),
.Y(n_21353)
);

NAND2xp5_ASAP7_75t_SL g21354 ( 
.A(n_21225),
.B(n_9146),
.Y(n_21354)
);

OR2x2_ASAP7_75t_L g21355 ( 
.A(n_21238),
.B(n_10968),
.Y(n_21355)
);

AOI21xp5_ASAP7_75t_L g21356 ( 
.A1(n_21275),
.A2(n_10334),
.B(n_10326),
.Y(n_21356)
);

NAND3xp33_ASAP7_75t_L g21357 ( 
.A(n_21269),
.B(n_9114),
.C(n_9107),
.Y(n_21357)
);

NOR2x1_ASAP7_75t_L g21358 ( 
.A(n_21198),
.B(n_9569),
.Y(n_21358)
);

AND2x2_ASAP7_75t_L g21359 ( 
.A(n_21165),
.B(n_10053),
.Y(n_21359)
);

OR2x2_ASAP7_75t_L g21360 ( 
.A(n_21197),
.B(n_10969),
.Y(n_21360)
);

OAI21xp5_ASAP7_75t_L g21361 ( 
.A1(n_21289),
.A2(n_10326),
.B(n_10322),
.Y(n_21361)
);

NAND2xp5_ASAP7_75t_L g21362 ( 
.A(n_21257),
.B(n_9679),
.Y(n_21362)
);

INVx1_ASAP7_75t_SL g21363 ( 
.A(n_21173),
.Y(n_21363)
);

NAND2xp5_ASAP7_75t_L g21364 ( 
.A(n_21211),
.B(n_9679),
.Y(n_21364)
);

INVx1_ASAP7_75t_L g21365 ( 
.A(n_21244),
.Y(n_21365)
);

NAND2xp5_ASAP7_75t_L g21366 ( 
.A(n_21300),
.B(n_10053),
.Y(n_21366)
);

BUFx4f_ASAP7_75t_SL g21367 ( 
.A(n_21247),
.Y(n_21367)
);

OR2x2_ASAP7_75t_L g21368 ( 
.A(n_21230),
.B(n_10969),
.Y(n_21368)
);

INVxp33_ASAP7_75t_L g21369 ( 
.A(n_21248),
.Y(n_21369)
);

INVx1_ASAP7_75t_L g21370 ( 
.A(n_21261),
.Y(n_21370)
);

NAND3xp33_ASAP7_75t_SL g21371 ( 
.A(n_21170),
.B(n_9834),
.C(n_9819),
.Y(n_21371)
);

OR2x2_ASAP7_75t_L g21372 ( 
.A(n_21264),
.B(n_10984),
.Y(n_21372)
);

INVx1_ASAP7_75t_L g21373 ( 
.A(n_21237),
.Y(n_21373)
);

NAND2xp5_ASAP7_75t_L g21374 ( 
.A(n_21243),
.B(n_10053),
.Y(n_21374)
);

CKINVDCx5p33_ASAP7_75t_R g21375 ( 
.A(n_21213),
.Y(n_21375)
);

INVx1_ASAP7_75t_L g21376 ( 
.A(n_21255),
.Y(n_21376)
);

AOI21xp5_ASAP7_75t_L g21377 ( 
.A1(n_21216),
.A2(n_10334),
.B(n_10336),
.Y(n_21377)
);

INVxp67_ASAP7_75t_L g21378 ( 
.A(n_21279),
.Y(n_21378)
);

INVx1_ASAP7_75t_L g21379 ( 
.A(n_21236),
.Y(n_21379)
);

NAND3xp33_ASAP7_75t_L g21380 ( 
.A(n_21284),
.B(n_9114),
.C(n_9107),
.Y(n_21380)
);

BUFx3_ASAP7_75t_L g21381 ( 
.A(n_21233),
.Y(n_21381)
);

XOR2x2_ASAP7_75t_L g21382 ( 
.A(n_21188),
.B(n_9834),
.Y(n_21382)
);

NAND2xp5_ASAP7_75t_L g21383 ( 
.A(n_21232),
.B(n_10053),
.Y(n_21383)
);

NOR2xp33_ASAP7_75t_SL g21384 ( 
.A(n_21293),
.B(n_7782),
.Y(n_21384)
);

NAND2xp5_ASAP7_75t_L g21385 ( 
.A(n_21201),
.B(n_10053),
.Y(n_21385)
);

XNOR2xp5_ASAP7_75t_L g21386 ( 
.A(n_21266),
.B(n_8454),
.Y(n_21386)
);

INVx1_ASAP7_75t_SL g21387 ( 
.A(n_21227),
.Y(n_21387)
);

INVx1_ASAP7_75t_L g21388 ( 
.A(n_21262),
.Y(n_21388)
);

NOR2xp67_ASAP7_75t_L g21389 ( 
.A(n_21294),
.B(n_8749),
.Y(n_21389)
);

INVx1_ASAP7_75t_L g21390 ( 
.A(n_21204),
.Y(n_21390)
);

INVx2_ASAP7_75t_SL g21391 ( 
.A(n_21223),
.Y(n_21391)
);

INVx1_ASAP7_75t_SL g21392 ( 
.A(n_21286),
.Y(n_21392)
);

NAND3xp33_ASAP7_75t_L g21393 ( 
.A(n_21265),
.B(n_9120),
.C(n_9114),
.Y(n_21393)
);

INVx1_ASAP7_75t_L g21394 ( 
.A(n_21219),
.Y(n_21394)
);

CKINVDCx20_ASAP7_75t_R g21395 ( 
.A(n_21295),
.Y(n_21395)
);

NAND2xp5_ASAP7_75t_L g21396 ( 
.A(n_21166),
.B(n_10053),
.Y(n_21396)
);

HB1xp67_ASAP7_75t_L g21397 ( 
.A(n_21277),
.Y(n_21397)
);

NAND2xp5_ASAP7_75t_L g21398 ( 
.A(n_21209),
.B(n_10053),
.Y(n_21398)
);

OAI21xp5_ASAP7_75t_L g21399 ( 
.A1(n_21220),
.A2(n_10334),
.B(n_10984),
.Y(n_21399)
);

INVx2_ASAP7_75t_L g21400 ( 
.A(n_21253),
.Y(n_21400)
);

INVx1_ASAP7_75t_L g21401 ( 
.A(n_21229),
.Y(n_21401)
);

AND2x2_ASAP7_75t_L g21402 ( 
.A(n_21270),
.B(n_10053),
.Y(n_21402)
);

NOR2xp67_ASAP7_75t_L g21403 ( 
.A(n_21206),
.B(n_8749),
.Y(n_21403)
);

XNOR2xp5_ASAP7_75t_L g21404 ( 
.A(n_21182),
.B(n_8454),
.Y(n_21404)
);

OAI221xp5_ASAP7_75t_L g21405 ( 
.A1(n_21196),
.A2(n_9834),
.B1(n_10002),
.B2(n_10103),
.C(n_9900),
.Y(n_21405)
);

NOR3xp33_ASAP7_75t_L g21406 ( 
.A(n_21234),
.B(n_10351),
.C(n_10341),
.Y(n_21406)
);

NAND2xp5_ASAP7_75t_L g21407 ( 
.A(n_21242),
.B(n_11108),
.Y(n_21407)
);

NOR2xp67_ASAP7_75t_SL g21408 ( 
.A(n_21254),
.B(n_8405),
.Y(n_21408)
);

INVx1_ASAP7_75t_L g21409 ( 
.A(n_21193),
.Y(n_21409)
);

INVx2_ASAP7_75t_SL g21410 ( 
.A(n_21163),
.Y(n_21410)
);

AND2x2_ASAP7_75t_L g21411 ( 
.A(n_21221),
.B(n_9863),
.Y(n_21411)
);

NAND3xp33_ASAP7_75t_L g21412 ( 
.A(n_21296),
.B(n_9120),
.C(n_9114),
.Y(n_21412)
);

NAND2xp5_ASAP7_75t_L g21413 ( 
.A(n_21168),
.B(n_21162),
.Y(n_21413)
);

OR2x2_ASAP7_75t_L g21414 ( 
.A(n_21273),
.B(n_10984),
.Y(n_21414)
);

OR2x2_ASAP7_75t_L g21415 ( 
.A(n_21185),
.B(n_10990),
.Y(n_21415)
);

AND2x2_ASAP7_75t_L g21416 ( 
.A(n_21297),
.B(n_9863),
.Y(n_21416)
);

NAND2xp5_ASAP7_75t_L g21417 ( 
.A(n_21252),
.B(n_21240),
.Y(n_21417)
);

AND2x4_ASAP7_75t_SL g21418 ( 
.A(n_21200),
.B(n_8203),
.Y(n_21418)
);

OR2x2_ASAP7_75t_L g21419 ( 
.A(n_21258),
.B(n_10990),
.Y(n_21419)
);

NAND2xp5_ASAP7_75t_SL g21420 ( 
.A(n_21251),
.B(n_9146),
.Y(n_21420)
);

INVx1_ASAP7_75t_L g21421 ( 
.A(n_21184),
.Y(n_21421)
);

INVxp67_ASAP7_75t_L g21422 ( 
.A(n_21191),
.Y(n_21422)
);

INVx1_ASAP7_75t_L g21423 ( 
.A(n_21298),
.Y(n_21423)
);

OAI32xp33_ASAP7_75t_L g21424 ( 
.A1(n_21202),
.A2(n_21190),
.A3(n_21189),
.B1(n_21177),
.B2(n_21176),
.Y(n_21424)
);

INVx2_ASAP7_75t_L g21425 ( 
.A(n_21175),
.Y(n_21425)
);

NOR2xp33_ASAP7_75t_L g21426 ( 
.A(n_21169),
.B(n_9900),
.Y(n_21426)
);

OAI21xp5_ASAP7_75t_L g21427 ( 
.A1(n_21195),
.A2(n_11023),
.B(n_10990),
.Y(n_21427)
);

NAND2xp5_ASAP7_75t_L g21428 ( 
.A(n_21256),
.B(n_11108),
.Y(n_21428)
);

AND2x2_ASAP7_75t_L g21429 ( 
.A(n_21281),
.B(n_9633),
.Y(n_21429)
);

INVxp67_ASAP7_75t_L g21430 ( 
.A(n_21192),
.Y(n_21430)
);

CKINVDCx16_ASAP7_75t_R g21431 ( 
.A(n_21239),
.Y(n_21431)
);

OAI31xp33_ASAP7_75t_SL g21432 ( 
.A1(n_21172),
.A2(n_10509),
.A3(n_10518),
.B(n_10507),
.Y(n_21432)
);

OR2x2_ASAP7_75t_L g21433 ( 
.A(n_21180),
.B(n_11023),
.Y(n_21433)
);

INVx1_ASAP7_75t_L g21434 ( 
.A(n_21178),
.Y(n_21434)
);

NAND2xp5_ASAP7_75t_L g21435 ( 
.A(n_21307),
.B(n_21290),
.Y(n_21435)
);

NAND3xp33_ASAP7_75t_L g21436 ( 
.A(n_21301),
.B(n_21160),
.C(n_21287),
.Y(n_21436)
);

INVx1_ASAP7_75t_L g21437 ( 
.A(n_21397),
.Y(n_21437)
);

AOI22xp33_ASAP7_75t_SL g21438 ( 
.A1(n_21306),
.A2(n_21288),
.B1(n_21228),
.B2(n_21174),
.Y(n_21438)
);

NOR2xp67_ASAP7_75t_L g21439 ( 
.A(n_21351),
.B(n_21245),
.Y(n_21439)
);

NAND4xp25_ASAP7_75t_L g21440 ( 
.A(n_21311),
.B(n_21218),
.C(n_9109),
.D(n_9113),
.Y(n_21440)
);

OAI22xp5_ASAP7_75t_L g21441 ( 
.A1(n_21326),
.A2(n_10085),
.B1(n_10095),
.B2(n_10075),
.Y(n_21441)
);

NOR2xp33_ASAP7_75t_L g21442 ( 
.A(n_21343),
.B(n_9900),
.Y(n_21442)
);

NOR2xp67_ASAP7_75t_L g21443 ( 
.A(n_21345),
.B(n_8933),
.Y(n_21443)
);

NOR3xp33_ASAP7_75t_L g21444 ( 
.A(n_21323),
.B(n_10341),
.C(n_10336),
.Y(n_21444)
);

NOR3xp33_ASAP7_75t_L g21445 ( 
.A(n_21309),
.B(n_10341),
.C(n_10336),
.Y(n_21445)
);

AND4x1_ASAP7_75t_L g21446 ( 
.A(n_21325),
.B(n_9852),
.C(n_9813),
.D(n_8892),
.Y(n_21446)
);

NAND2xp5_ASAP7_75t_L g21447 ( 
.A(n_21304),
.B(n_7706),
.Y(n_21447)
);

NOR3xp33_ASAP7_75t_L g21448 ( 
.A(n_21308),
.B(n_10351),
.C(n_10507),
.Y(n_21448)
);

NOR2xp33_ASAP7_75t_L g21449 ( 
.A(n_21431),
.B(n_21367),
.Y(n_21449)
);

AND2x2_ASAP7_75t_L g21450 ( 
.A(n_21324),
.B(n_11493),
.Y(n_21450)
);

NOR3xp33_ASAP7_75t_L g21451 ( 
.A(n_21302),
.B(n_10351),
.C(n_10507),
.Y(n_21451)
);

NAND2xp5_ASAP7_75t_L g21452 ( 
.A(n_21342),
.B(n_7706),
.Y(n_21452)
);

NOR3xp33_ASAP7_75t_L g21453 ( 
.A(n_21303),
.B(n_21338),
.C(n_21339),
.Y(n_21453)
);

NOR2x1_ASAP7_75t_L g21454 ( 
.A(n_21318),
.B(n_9569),
.Y(n_21454)
);

AOI22xp5_ASAP7_75t_L g21455 ( 
.A1(n_21314),
.A2(n_21333),
.B1(n_21319),
.B2(n_21313),
.Y(n_21455)
);

AND2x4_ASAP7_75t_L g21456 ( 
.A(n_21403),
.B(n_9146),
.Y(n_21456)
);

AOI211xp5_ASAP7_75t_L g21457 ( 
.A1(n_21369),
.A2(n_10579),
.B(n_10562),
.C(n_11023),
.Y(n_21457)
);

NAND4xp75_ASAP7_75t_L g21458 ( 
.A(n_21391),
.B(n_11114),
.C(n_11146),
.D(n_11108),
.Y(n_21458)
);

NAND4xp75_ASAP7_75t_L g21459 ( 
.A(n_21365),
.B(n_11114),
.C(n_11146),
.D(n_11108),
.Y(n_21459)
);

AND2x2_ASAP7_75t_SL g21460 ( 
.A(n_21312),
.B(n_8768),
.Y(n_21460)
);

HB1xp67_ASAP7_75t_L g21461 ( 
.A(n_21352),
.Y(n_21461)
);

NOR3xp33_ASAP7_75t_L g21462 ( 
.A(n_21322),
.B(n_10518),
.C(n_10509),
.Y(n_21462)
);

AOI21xp5_ASAP7_75t_L g21463 ( 
.A1(n_21337),
.A2(n_10518),
.B(n_10509),
.Y(n_21463)
);

NAND3xp33_ASAP7_75t_L g21464 ( 
.A(n_21331),
.B(n_21430),
.C(n_21375),
.Y(n_21464)
);

OAI211xp5_ASAP7_75t_L g21465 ( 
.A1(n_21346),
.A2(n_21363),
.B(n_21392),
.C(n_21378),
.Y(n_21465)
);

NAND3xp33_ASAP7_75t_L g21466 ( 
.A(n_21331),
.B(n_9221),
.C(n_9216),
.Y(n_21466)
);

AOI211x1_ASAP7_75t_L g21467 ( 
.A1(n_21424),
.A2(n_9227),
.B(n_9235),
.C(n_9221),
.Y(n_21467)
);

NOR2x1_ASAP7_75t_L g21468 ( 
.A(n_21310),
.B(n_9569),
.Y(n_21468)
);

OA22x2_ASAP7_75t_L g21469 ( 
.A1(n_21388),
.A2(n_11039),
.B1(n_11030),
.B2(n_11040),
.Y(n_21469)
);

OAI211xp5_ASAP7_75t_L g21470 ( 
.A1(n_21336),
.A2(n_9227),
.B(n_9234),
.C(n_9221),
.Y(n_21470)
);

NOR2x1_ASAP7_75t_L g21471 ( 
.A(n_21348),
.B(n_9569),
.Y(n_21471)
);

NOR2x1_ASAP7_75t_L g21472 ( 
.A(n_21347),
.B(n_9572),
.Y(n_21472)
);

NAND4xp25_ASAP7_75t_L g21473 ( 
.A(n_21316),
.B(n_9109),
.C(n_9113),
.D(n_9089),
.Y(n_21473)
);

OR2x2_ASAP7_75t_L g21474 ( 
.A(n_21383),
.B(n_11030),
.Y(n_21474)
);

AND5x1_ASAP7_75t_L g21475 ( 
.A(n_21384),
.B(n_8893),
.C(n_8925),
.D(n_8885),
.E(n_12839),
.Y(n_21475)
);

NAND3xp33_ASAP7_75t_SL g21476 ( 
.A(n_21387),
.B(n_9834),
.C(n_8699),
.Y(n_21476)
);

NOR3x2_ASAP7_75t_L g21477 ( 
.A(n_21331),
.B(n_12897),
.C(n_7907),
.Y(n_21477)
);

INVxp67_ASAP7_75t_SL g21478 ( 
.A(n_21422),
.Y(n_21478)
);

AOI211xp5_ASAP7_75t_SL g21479 ( 
.A1(n_21434),
.A2(n_10095),
.B(n_10107),
.C(n_10085),
.Y(n_21479)
);

NAND3xp33_ASAP7_75t_SL g21480 ( 
.A(n_21395),
.B(n_8699),
.C(n_8796),
.Y(n_21480)
);

OAI211xp5_ASAP7_75t_L g21481 ( 
.A1(n_21425),
.A2(n_21330),
.B(n_21334),
.C(n_21373),
.Y(n_21481)
);

NOR2x1p5_ASAP7_75t_L g21482 ( 
.A(n_21381),
.B(n_21370),
.Y(n_21482)
);

NOR2x1_ASAP7_75t_L g21483 ( 
.A(n_21421),
.B(n_9572),
.Y(n_21483)
);

INVx1_ASAP7_75t_L g21484 ( 
.A(n_21413),
.Y(n_21484)
);

NAND4xp25_ASAP7_75t_L g21485 ( 
.A(n_21379),
.B(n_9109),
.C(n_9113),
.D(n_9089),
.Y(n_21485)
);

NAND4xp25_ASAP7_75t_L g21486 ( 
.A(n_21376),
.B(n_9109),
.C(n_9113),
.D(n_9089),
.Y(n_21486)
);

NOR4xp75_ASAP7_75t_L g21487 ( 
.A(n_21410),
.B(n_9807),
.C(n_9804),
.D(n_9803),
.Y(n_21487)
);

NAND4xp25_ASAP7_75t_L g21488 ( 
.A(n_21401),
.B(n_9109),
.C(n_9113),
.D(n_9089),
.Y(n_21488)
);

NOR2x1p5_ASAP7_75t_L g21489 ( 
.A(n_21400),
.B(n_7981),
.Y(n_21489)
);

NOR3xp33_ASAP7_75t_L g21490 ( 
.A(n_21423),
.B(n_21409),
.C(n_21417),
.Y(n_21490)
);

HB1xp67_ASAP7_75t_L g21491 ( 
.A(n_21394),
.Y(n_21491)
);

AND2x2_ASAP7_75t_L g21492 ( 
.A(n_21402),
.B(n_11516),
.Y(n_21492)
);

NAND4xp75_ASAP7_75t_L g21493 ( 
.A(n_21335),
.B(n_11114),
.C(n_11146),
.D(n_11108),
.Y(n_21493)
);

AND2x2_ASAP7_75t_SL g21494 ( 
.A(n_21390),
.B(n_8768),
.Y(n_21494)
);

NOR2x1_ASAP7_75t_L g21495 ( 
.A(n_21358),
.B(n_9572),
.Y(n_21495)
);

NAND2xp5_ASAP7_75t_L g21496 ( 
.A(n_21418),
.B(n_21389),
.Y(n_21496)
);

NOR3xp33_ASAP7_75t_L g21497 ( 
.A(n_21350),
.B(n_10519),
.C(n_11508),
.Y(n_21497)
);

NOR3xp33_ASAP7_75t_L g21498 ( 
.A(n_21356),
.B(n_10519),
.C(n_11511),
.Y(n_21498)
);

NOR2x1p5_ASAP7_75t_L g21499 ( 
.A(n_21305),
.B(n_21366),
.Y(n_21499)
);

NOR2x1_ASAP7_75t_L g21500 ( 
.A(n_21321),
.B(n_21355),
.Y(n_21500)
);

NOR3xp33_ASAP7_75t_L g21501 ( 
.A(n_21329),
.B(n_10519),
.C(n_11511),
.Y(n_21501)
);

NOR3xp33_ASAP7_75t_L g21502 ( 
.A(n_21396),
.B(n_11516),
.C(n_11515),
.Y(n_21502)
);

NAND3xp33_ASAP7_75t_SL g21503 ( 
.A(n_21317),
.B(n_8699),
.C(n_8881),
.Y(n_21503)
);

NAND2x1p5_ASAP7_75t_L g21504 ( 
.A(n_21340),
.B(n_11515),
.Y(n_21504)
);

INVx1_ASAP7_75t_L g21505 ( 
.A(n_21408),
.Y(n_21505)
);

NAND2xp5_ASAP7_75t_L g21506 ( 
.A(n_21315),
.B(n_7706),
.Y(n_21506)
);

NOR3xp33_ASAP7_75t_SL g21507 ( 
.A(n_21385),
.B(n_10095),
.C(n_10085),
.Y(n_21507)
);

NOR2x1p5_ASAP7_75t_L g21508 ( 
.A(n_21398),
.B(n_7992),
.Y(n_21508)
);

INVx1_ASAP7_75t_L g21509 ( 
.A(n_21382),
.Y(n_21509)
);

NAND3x1_ASAP7_75t_L g21510 ( 
.A(n_21349),
.B(n_9154),
.C(n_9130),
.Y(n_21510)
);

NAND4xp25_ASAP7_75t_L g21511 ( 
.A(n_21320),
.B(n_9129),
.C(n_9113),
.D(n_8915),
.Y(n_21511)
);

NAND4xp75_ASAP7_75t_L g21512 ( 
.A(n_21354),
.B(n_11146),
.C(n_11160),
.D(n_11114),
.Y(n_21512)
);

NOR2xp67_ASAP7_75t_L g21513 ( 
.A(n_21362),
.B(n_8933),
.Y(n_21513)
);

INVx1_ASAP7_75t_L g21514 ( 
.A(n_21407),
.Y(n_21514)
);

NOR2x1_ASAP7_75t_L g21515 ( 
.A(n_21420),
.B(n_9572),
.Y(n_21515)
);

INVx1_ASAP7_75t_L g21516 ( 
.A(n_21416),
.Y(n_21516)
);

NOR4xp75_ASAP7_75t_L g21517 ( 
.A(n_21374),
.B(n_9807),
.C(n_9804),
.D(n_9803),
.Y(n_21517)
);

NAND2xp5_ASAP7_75t_L g21518 ( 
.A(n_21406),
.B(n_7706),
.Y(n_21518)
);

INVx3_ASAP7_75t_L g21519 ( 
.A(n_21372),
.Y(n_21519)
);

NOR2x1_ASAP7_75t_L g21520 ( 
.A(n_21415),
.B(n_9572),
.Y(n_21520)
);

INVx2_ASAP7_75t_SL g21521 ( 
.A(n_21359),
.Y(n_21521)
);

NAND3xp33_ASAP7_75t_SL g21522 ( 
.A(n_21364),
.B(n_8699),
.C(n_8881),
.Y(n_21522)
);

NOR2xp33_ASAP7_75t_L g21523 ( 
.A(n_21426),
.B(n_10002),
.Y(n_21523)
);

NAND4xp25_ASAP7_75t_L g21524 ( 
.A(n_21332),
.B(n_9129),
.C(n_9113),
.D(n_8915),
.Y(n_21524)
);

NOR2x1_ASAP7_75t_L g21525 ( 
.A(n_21371),
.B(n_9572),
.Y(n_21525)
);

AOI211xp5_ASAP7_75t_L g21526 ( 
.A1(n_21386),
.A2(n_10579),
.B(n_10562),
.C(n_11030),
.Y(n_21526)
);

NOR3x1_ASAP7_75t_L g21527 ( 
.A(n_21428),
.B(n_11039),
.C(n_11040),
.Y(n_21527)
);

NOR2x1_ASAP7_75t_L g21528 ( 
.A(n_21344),
.B(n_21341),
.Y(n_21528)
);

NAND3x1_ASAP7_75t_L g21529 ( 
.A(n_21411),
.B(n_9154),
.C(n_9130),
.Y(n_21529)
);

NAND4xp75_ASAP7_75t_L g21530 ( 
.A(n_21377),
.B(n_11146),
.C(n_11160),
.D(n_11114),
.Y(n_21530)
);

INVx1_ASAP7_75t_L g21531 ( 
.A(n_21433),
.Y(n_21531)
);

INVxp67_ASAP7_75t_SL g21532 ( 
.A(n_21404),
.Y(n_21532)
);

NOR2xp67_ASAP7_75t_L g21533 ( 
.A(n_21368),
.B(n_8973),
.Y(n_21533)
);

NAND4xp25_ASAP7_75t_L g21534 ( 
.A(n_21361),
.B(n_9129),
.C(n_9113),
.D(n_8924),
.Y(n_21534)
);

NAND2xp5_ASAP7_75t_SL g21535 ( 
.A(n_21414),
.B(n_9146),
.Y(n_21535)
);

NAND2xp5_ASAP7_75t_L g21536 ( 
.A(n_21360),
.B(n_7706),
.Y(n_21536)
);

AND5x1_ASAP7_75t_L g21537 ( 
.A(n_21432),
.B(n_8893),
.C(n_8925),
.D(n_8885),
.E(n_8924),
.Y(n_21537)
);

AOI211x1_ASAP7_75t_L g21538 ( 
.A1(n_21353),
.A2(n_9234),
.B(n_9235),
.C(n_9227),
.Y(n_21538)
);

NAND3xp33_ASAP7_75t_L g21539 ( 
.A(n_21429),
.B(n_9234),
.C(n_9227),
.Y(n_21539)
);

INVxp67_ASAP7_75t_L g21540 ( 
.A(n_21419),
.Y(n_21540)
);

NOR3xp33_ASAP7_75t_L g21541 ( 
.A(n_21328),
.B(n_11516),
.C(n_11515),
.Y(n_21541)
);

AND2x2_ASAP7_75t_L g21542 ( 
.A(n_21399),
.B(n_11160),
.Y(n_21542)
);

NAND3xp33_ASAP7_75t_SL g21543 ( 
.A(n_21405),
.B(n_8699),
.C(n_8928),
.Y(n_21543)
);

NAND3xp33_ASAP7_75t_SL g21544 ( 
.A(n_21393),
.B(n_8928),
.C(n_10095),
.Y(n_21544)
);

NOR2x1_ASAP7_75t_L g21545 ( 
.A(n_21412),
.B(n_9572),
.Y(n_21545)
);

NOR2xp33_ASAP7_75t_L g21546 ( 
.A(n_21449),
.B(n_21327),
.Y(n_21546)
);

AOI22xp5_ASAP7_75t_L g21547 ( 
.A1(n_21453),
.A2(n_21357),
.B1(n_21380),
.B2(n_21427),
.Y(n_21547)
);

AOI22xp5_ASAP7_75t_L g21548 ( 
.A1(n_21442),
.A2(n_11165),
.B1(n_11201),
.B2(n_11160),
.Y(n_21548)
);

NAND2xp5_ASAP7_75t_L g21549 ( 
.A(n_21437),
.B(n_7706),
.Y(n_21549)
);

NOR2x1p5_ASAP7_75t_L g21550 ( 
.A(n_21532),
.B(n_7992),
.Y(n_21550)
);

NAND2xp5_ASAP7_75t_L g21551 ( 
.A(n_21491),
.B(n_7706),
.Y(n_21551)
);

INVx1_ASAP7_75t_L g21552 ( 
.A(n_21461),
.Y(n_21552)
);

INVx1_ASAP7_75t_L g21553 ( 
.A(n_21435),
.Y(n_21553)
);

INVx1_ASAP7_75t_L g21554 ( 
.A(n_21436),
.Y(n_21554)
);

NAND3xp33_ASAP7_75t_L g21555 ( 
.A(n_21490),
.B(n_11165),
.C(n_11160),
.Y(n_21555)
);

AND2x4_ASAP7_75t_SL g21556 ( 
.A(n_21455),
.B(n_8206),
.Y(n_21556)
);

NOR2x1_ASAP7_75t_L g21557 ( 
.A(n_21464),
.B(n_9572),
.Y(n_21557)
);

AOI22xp5_ASAP7_75t_L g21558 ( 
.A1(n_21465),
.A2(n_11165),
.B1(n_11201),
.B2(n_11160),
.Y(n_21558)
);

INVx1_ASAP7_75t_L g21559 ( 
.A(n_21443),
.Y(n_21559)
);

INVx1_ASAP7_75t_L g21560 ( 
.A(n_21505),
.Y(n_21560)
);

AOI22xp5_ASAP7_75t_L g21561 ( 
.A1(n_21482),
.A2(n_11201),
.B1(n_11165),
.B2(n_9183),
.Y(n_21561)
);

INVx2_ASAP7_75t_L g21562 ( 
.A(n_21489),
.Y(n_21562)
);

AND2x4_ASAP7_75t_L g21563 ( 
.A(n_21456),
.B(n_9182),
.Y(n_21563)
);

NAND2xp5_ASAP7_75t_L g21564 ( 
.A(n_21478),
.B(n_21513),
.Y(n_21564)
);

INVx1_ASAP7_75t_L g21565 ( 
.A(n_21529),
.Y(n_21565)
);

INVx1_ASAP7_75t_L g21566 ( 
.A(n_21496),
.Y(n_21566)
);

NAND2xp5_ASAP7_75t_L g21567 ( 
.A(n_21439),
.B(n_7762),
.Y(n_21567)
);

NAND2xp5_ASAP7_75t_L g21568 ( 
.A(n_21521),
.B(n_7762),
.Y(n_21568)
);

INVx2_ASAP7_75t_L g21569 ( 
.A(n_21499),
.Y(n_21569)
);

INVx1_ASAP7_75t_L g21570 ( 
.A(n_21528),
.Y(n_21570)
);

NAND2xp5_ASAP7_75t_L g21571 ( 
.A(n_21533),
.B(n_7762),
.Y(n_21571)
);

NOR2x1_ASAP7_75t_L g21572 ( 
.A(n_21481),
.B(n_9239),
.Y(n_21572)
);

INVx1_ASAP7_75t_L g21573 ( 
.A(n_21500),
.Y(n_21573)
);

OR2x2_ASAP7_75t_L g21574 ( 
.A(n_21535),
.B(n_11039),
.Y(n_21574)
);

AOI22xp5_ASAP7_75t_L g21575 ( 
.A1(n_21484),
.A2(n_11201),
.B1(n_11165),
.B2(n_9183),
.Y(n_21575)
);

INVx2_ASAP7_75t_L g21576 ( 
.A(n_21508),
.Y(n_21576)
);

INVx1_ASAP7_75t_L g21577 ( 
.A(n_21519),
.Y(n_21577)
);

INVx1_ASAP7_75t_L g21578 ( 
.A(n_21519),
.Y(n_21578)
);

AOI22xp5_ASAP7_75t_L g21579 ( 
.A1(n_21509),
.A2(n_11201),
.B1(n_11165),
.B2(n_9183),
.Y(n_21579)
);

INVx1_ASAP7_75t_L g21580 ( 
.A(n_21514),
.Y(n_21580)
);

INVx1_ASAP7_75t_SL g21581 ( 
.A(n_21516),
.Y(n_21581)
);

INVx1_ASAP7_75t_L g21582 ( 
.A(n_21531),
.Y(n_21582)
);

AOI22xp5_ASAP7_75t_L g21583 ( 
.A1(n_21543),
.A2(n_11201),
.B1(n_9183),
.B2(n_9198),
.Y(n_21583)
);

INVx1_ASAP7_75t_L g21584 ( 
.A(n_21540),
.Y(n_21584)
);

INVx1_ASAP7_75t_L g21585 ( 
.A(n_21438),
.Y(n_21585)
);

AND3x2_ASAP7_75t_L g21586 ( 
.A(n_21526),
.B(n_9183),
.C(n_9182),
.Y(n_21586)
);

INVx2_ASAP7_75t_L g21587 ( 
.A(n_21515),
.Y(n_21587)
);

INVx1_ASAP7_75t_L g21588 ( 
.A(n_21456),
.Y(n_21588)
);

NOR2x2_ASAP7_75t_L g21589 ( 
.A(n_21493),
.B(n_10002),
.Y(n_21589)
);

INVx1_ASAP7_75t_L g21590 ( 
.A(n_21506),
.Y(n_21590)
);

INVx2_ASAP7_75t_L g21591 ( 
.A(n_21474),
.Y(n_21591)
);

AOI22xp5_ASAP7_75t_L g21592 ( 
.A1(n_21544),
.A2(n_9183),
.B1(n_9198),
.B2(n_9182),
.Y(n_21592)
);

AOI22xp5_ASAP7_75t_L g21593 ( 
.A1(n_21523),
.A2(n_9183),
.B1(n_9198),
.B2(n_9182),
.Y(n_21593)
);

AOI22xp5_ASAP7_75t_L g21594 ( 
.A1(n_21480),
.A2(n_9198),
.B1(n_9217),
.B2(n_9182),
.Y(n_21594)
);

INVxp67_ASAP7_75t_L g21595 ( 
.A(n_21492),
.Y(n_21595)
);

NAND2xp5_ASAP7_75t_SL g21596 ( 
.A(n_21452),
.B(n_9182),
.Y(n_21596)
);

INVx1_ASAP7_75t_L g21597 ( 
.A(n_21539),
.Y(n_21597)
);

NAND2xp5_ASAP7_75t_L g21598 ( 
.A(n_21507),
.B(n_7762),
.Y(n_21598)
);

INVx1_ASAP7_75t_SL g21599 ( 
.A(n_21536),
.Y(n_21599)
);

AOI22xp5_ASAP7_75t_L g21600 ( 
.A1(n_21522),
.A2(n_9198),
.B1(n_9217),
.B2(n_9182),
.Y(n_21600)
);

INVx2_ASAP7_75t_L g21601 ( 
.A(n_21520),
.Y(n_21601)
);

NOR2x1_ASAP7_75t_L g21602 ( 
.A(n_21495),
.B(n_8990),
.Y(n_21602)
);

BUFx6f_ASAP7_75t_L g21603 ( 
.A(n_21503),
.Y(n_21603)
);

AOI22xp33_ASAP7_75t_L g21604 ( 
.A1(n_21440),
.A2(n_21541),
.B1(n_21447),
.B2(n_21511),
.Y(n_21604)
);

NOR2xp67_ASAP7_75t_L g21605 ( 
.A(n_21518),
.B(n_8973),
.Y(n_21605)
);

OR2x2_ASAP7_75t_L g21606 ( 
.A(n_21524),
.B(n_11040),
.Y(n_21606)
);

HB1xp67_ASAP7_75t_L g21607 ( 
.A(n_21525),
.Y(n_21607)
);

NOR2x1p5_ASAP7_75t_L g21608 ( 
.A(n_21473),
.B(n_21534),
.Y(n_21608)
);

INVx1_ASAP7_75t_L g21609 ( 
.A(n_21545),
.Y(n_21609)
);

NAND2xp5_ASAP7_75t_L g21610 ( 
.A(n_21538),
.B(n_7762),
.Y(n_21610)
);

INVx1_ASAP7_75t_L g21611 ( 
.A(n_21466),
.Y(n_21611)
);

INVx2_ASAP7_75t_L g21612 ( 
.A(n_21527),
.Y(n_21612)
);

AOI22xp5_ASAP7_75t_L g21613 ( 
.A1(n_21510),
.A2(n_9217),
.B1(n_9222),
.B2(n_9198),
.Y(n_21613)
);

INVx1_ASAP7_75t_L g21614 ( 
.A(n_21467),
.Y(n_21614)
);

INVx1_ASAP7_75t_L g21615 ( 
.A(n_21483),
.Y(n_21615)
);

INVx1_ASAP7_75t_L g21616 ( 
.A(n_21542),
.Y(n_21616)
);

OAI22xp5_ASAP7_75t_L g21617 ( 
.A1(n_21512),
.A2(n_10123),
.B1(n_10107),
.B2(n_9235),
.Y(n_21617)
);

INVx1_ASAP7_75t_L g21618 ( 
.A(n_21454),
.Y(n_21618)
);

OR2x2_ASAP7_75t_L g21619 ( 
.A(n_21485),
.B(n_11042),
.Y(n_21619)
);

AOI22xp5_ASAP7_75t_L g21620 ( 
.A1(n_21450),
.A2(n_9217),
.B1(n_9222),
.B2(n_9198),
.Y(n_21620)
);

INVx1_ASAP7_75t_L g21621 ( 
.A(n_21471),
.Y(n_21621)
);

NAND2xp5_ASAP7_75t_SL g21622 ( 
.A(n_21468),
.B(n_9198),
.Y(n_21622)
);

INVx1_ASAP7_75t_L g21623 ( 
.A(n_21472),
.Y(n_21623)
);

AOI22xp5_ASAP7_75t_L g21624 ( 
.A1(n_21502),
.A2(n_9217),
.B1(n_9222),
.B2(n_9198),
.Y(n_21624)
);

INVx1_ASAP7_75t_L g21625 ( 
.A(n_21530),
.Y(n_21625)
);

INVx1_ASAP7_75t_SL g21626 ( 
.A(n_21458),
.Y(n_21626)
);

AOI22xp5_ASAP7_75t_L g21627 ( 
.A1(n_21498),
.A2(n_9222),
.B1(n_9241),
.B2(n_9217),
.Y(n_21627)
);

NAND2xp5_ASAP7_75t_L g21628 ( 
.A(n_21479),
.B(n_7762),
.Y(n_21628)
);

INVx1_ASAP7_75t_L g21629 ( 
.A(n_21504),
.Y(n_21629)
);

AOI22xp5_ASAP7_75t_L g21630 ( 
.A1(n_21488),
.A2(n_9222),
.B1(n_9241),
.B2(n_9217),
.Y(n_21630)
);

INVx1_ASAP7_75t_L g21631 ( 
.A(n_21470),
.Y(n_21631)
);

INVxp67_ASAP7_75t_L g21632 ( 
.A(n_21459),
.Y(n_21632)
);

NOR2x1_ASAP7_75t_L g21633 ( 
.A(n_21476),
.B(n_8990),
.Y(n_21633)
);

AO22x2_ASAP7_75t_L g21634 ( 
.A1(n_21441),
.A2(n_9138),
.B1(n_9151),
.B2(n_9120),
.Y(n_21634)
);

INVx1_ASAP7_75t_L g21635 ( 
.A(n_21444),
.Y(n_21635)
);

INVx1_ASAP7_75t_L g21636 ( 
.A(n_21445),
.Y(n_21636)
);

INVx1_ASAP7_75t_L g21637 ( 
.A(n_21486),
.Y(n_21637)
);

INVx1_ASAP7_75t_L g21638 ( 
.A(n_21446),
.Y(n_21638)
);

INVxp67_ASAP7_75t_SL g21639 ( 
.A(n_21537),
.Y(n_21639)
);

INVx5_ASAP7_75t_L g21640 ( 
.A(n_21569),
.Y(n_21640)
);

AND4x1_ASAP7_75t_L g21641 ( 
.A(n_21552),
.B(n_21451),
.C(n_21448),
.D(n_21463),
.Y(n_21641)
);

AND4x2_ASAP7_75t_L g21642 ( 
.A(n_21572),
.B(n_21475),
.C(n_21517),
.D(n_21469),
.Y(n_21642)
);

OAI22x1_ASAP7_75t_SL g21643 ( 
.A1(n_21585),
.A2(n_21477),
.B1(n_21487),
.B2(n_21460),
.Y(n_21643)
);

OAI211xp5_ASAP7_75t_L g21644 ( 
.A1(n_21573),
.A2(n_21501),
.B(n_21497),
.C(n_21462),
.Y(n_21644)
);

NOR2x1_ASAP7_75t_L g21645 ( 
.A(n_21588),
.B(n_21494),
.Y(n_21645)
);

OAI22xp33_ASAP7_75t_L g21646 ( 
.A1(n_21570),
.A2(n_21457),
.B1(n_9235),
.B2(n_9238),
.Y(n_21646)
);

NOR3xp33_ASAP7_75t_L g21647 ( 
.A(n_21554),
.B(n_10579),
.C(n_10562),
.Y(n_21647)
);

HB1xp67_ASAP7_75t_L g21648 ( 
.A(n_21562),
.Y(n_21648)
);

O2A1O1Ixp5_ASAP7_75t_L g21649 ( 
.A1(n_21612),
.A2(n_9120),
.B(n_9151),
.C(n_9138),
.Y(n_21649)
);

NOR3xp33_ASAP7_75t_SL g21650 ( 
.A(n_21546),
.B(n_10107),
.C(n_10123),
.Y(n_21650)
);

NAND2xp5_ASAP7_75t_L g21651 ( 
.A(n_21556),
.B(n_9991),
.Y(n_21651)
);

AOI211x1_ASAP7_75t_L g21652 ( 
.A1(n_21567),
.A2(n_10123),
.B(n_10107),
.C(n_9238),
.Y(n_21652)
);

NAND3xp33_ASAP7_75t_SL g21653 ( 
.A(n_21581),
.B(n_10123),
.C(n_7999),
.Y(n_21653)
);

AOI21xp5_ASAP7_75t_L g21654 ( 
.A1(n_21564),
.A2(n_10297),
.B(n_10290),
.Y(n_21654)
);

INVx1_ASAP7_75t_L g21655 ( 
.A(n_21614),
.Y(n_21655)
);

NOR2x1_ASAP7_75t_L g21656 ( 
.A(n_21577),
.B(n_8990),
.Y(n_21656)
);

OAI221xp5_ASAP7_75t_SL g21657 ( 
.A1(n_21604),
.A2(n_9257),
.B1(n_9276),
.B2(n_9238),
.C(n_9234),
.Y(n_21657)
);

AND2x2_ASAP7_75t_L g21658 ( 
.A(n_21576),
.B(n_10002),
.Y(n_21658)
);

HB1xp67_ASAP7_75t_L g21659 ( 
.A(n_21629),
.Y(n_21659)
);

NAND4xp75_ASAP7_75t_L g21660 ( 
.A(n_21578),
.B(n_11363),
.C(n_11373),
.D(n_11347),
.Y(n_21660)
);

NAND3xp33_ASAP7_75t_L g21661 ( 
.A(n_21560),
.B(n_9257),
.C(n_9238),
.Y(n_21661)
);

NOR2x1_ASAP7_75t_L g21662 ( 
.A(n_21601),
.B(n_8990),
.Y(n_21662)
);

NOR2xp67_ASAP7_75t_L g21663 ( 
.A(n_21595),
.B(n_8973),
.Y(n_21663)
);

NAND4xp75_ASAP7_75t_L g21664 ( 
.A(n_21553),
.B(n_11363),
.C(n_11373),
.D(n_11347),
.Y(n_21664)
);

NAND3xp33_ASAP7_75t_L g21665 ( 
.A(n_21603),
.B(n_21582),
.C(n_21580),
.Y(n_21665)
);

AND2x4_ASAP7_75t_L g21666 ( 
.A(n_21563),
.B(n_9466),
.Y(n_21666)
);

INVx5_ASAP7_75t_L g21667 ( 
.A(n_21603),
.Y(n_21667)
);

NOR3xp33_ASAP7_75t_SL g21668 ( 
.A(n_21584),
.B(n_7709),
.C(n_7704),
.Y(n_21668)
);

NAND2xp5_ASAP7_75t_L g21669 ( 
.A(n_21559),
.B(n_9991),
.Y(n_21669)
);

OR2x2_ASAP7_75t_L g21670 ( 
.A(n_21596),
.B(n_11042),
.Y(n_21670)
);

NOR2xp33_ASAP7_75t_R g21671 ( 
.A(n_21566),
.B(n_8814),
.Y(n_21671)
);

NAND2x1p5_ASAP7_75t_L g21672 ( 
.A(n_21599),
.B(n_8716),
.Y(n_21672)
);

AOI221xp5_ASAP7_75t_L g21673 ( 
.A1(n_21632),
.A2(n_9410),
.B1(n_9463),
.B2(n_9357),
.C(n_9307),
.Y(n_21673)
);

NOR3xp33_ASAP7_75t_L g21674 ( 
.A(n_21616),
.B(n_10297),
.C(n_10290),
.Y(n_21674)
);

INVx2_ASAP7_75t_SL g21675 ( 
.A(n_21550),
.Y(n_21675)
);

AND3x4_ASAP7_75t_L g21676 ( 
.A(n_21591),
.B(n_8740),
.C(n_8716),
.Y(n_21676)
);

NAND4xp25_ASAP7_75t_L g21677 ( 
.A(n_21637),
.B(n_9129),
.C(n_8949),
.D(n_8959),
.Y(n_21677)
);

XNOR2xp5_ASAP7_75t_L g21678 ( 
.A(n_21608),
.B(n_8454),
.Y(n_21678)
);

AND2x4_ASAP7_75t_L g21679 ( 
.A(n_21638),
.B(n_9466),
.Y(n_21679)
);

OAI22xp5_ASAP7_75t_SL g21680 ( 
.A1(n_21626),
.A2(n_8768),
.B1(n_9101),
.B2(n_9079),
.Y(n_21680)
);

AOI221xp5_ASAP7_75t_SL g21681 ( 
.A1(n_21631),
.A2(n_9360),
.B1(n_9480),
.B2(n_9317),
.C(n_9257),
.Y(n_21681)
);

OAI211xp5_ASAP7_75t_L g21682 ( 
.A1(n_21547),
.A2(n_21625),
.B(n_21635),
.C(n_21590),
.Y(n_21682)
);

NOR3xp33_ASAP7_75t_SL g21683 ( 
.A(n_21565),
.B(n_7709),
.C(n_7704),
.Y(n_21683)
);

INVx1_ASAP7_75t_L g21684 ( 
.A(n_21549),
.Y(n_21684)
);

NAND2xp5_ASAP7_75t_L g21685 ( 
.A(n_21639),
.B(n_9991),
.Y(n_21685)
);

OR2x2_ASAP7_75t_L g21686 ( 
.A(n_21551),
.B(n_11042),
.Y(n_21686)
);

AND3x2_ASAP7_75t_L g21687 ( 
.A(n_21607),
.B(n_9222),
.C(n_9217),
.Y(n_21687)
);

AND2x4_ASAP7_75t_L g21688 ( 
.A(n_21568),
.B(n_9466),
.Y(n_21688)
);

OR3x2_ASAP7_75t_L g21689 ( 
.A(n_21636),
.B(n_9154),
.C(n_9130),
.Y(n_21689)
);

NOR3xp33_ASAP7_75t_L g21690 ( 
.A(n_21609),
.B(n_10297),
.C(n_10290),
.Y(n_21690)
);

INVx1_ASAP7_75t_L g21691 ( 
.A(n_21597),
.Y(n_21691)
);

NAND2x1p5_ASAP7_75t_L g21692 ( 
.A(n_21615),
.B(n_8716),
.Y(n_21692)
);

INVx1_ASAP7_75t_L g21693 ( 
.A(n_21611),
.Y(n_21693)
);

OR2x2_ASAP7_75t_L g21694 ( 
.A(n_21622),
.B(n_11053),
.Y(n_21694)
);

NOR4xp75_ASAP7_75t_L g21695 ( 
.A(n_21571),
.B(n_8835),
.C(n_9154),
.D(n_9130),
.Y(n_21695)
);

OR2x2_ASAP7_75t_L g21696 ( 
.A(n_21606),
.B(n_11053),
.Y(n_21696)
);

OR2x2_ASAP7_75t_L g21697 ( 
.A(n_21619),
.B(n_11053),
.Y(n_21697)
);

AND3x4_ASAP7_75t_L g21698 ( 
.A(n_21587),
.B(n_8740),
.C(n_8716),
.Y(n_21698)
);

AND3x1_ASAP7_75t_L g21699 ( 
.A(n_21621),
.B(n_9316),
.C(n_9302),
.Y(n_21699)
);

AND3x4_ASAP7_75t_L g21700 ( 
.A(n_21605),
.B(n_8740),
.C(n_8716),
.Y(n_21700)
);

INVx1_ASAP7_75t_L g21701 ( 
.A(n_21623),
.Y(n_21701)
);

NAND2xp5_ASAP7_75t_L g21702 ( 
.A(n_21586),
.B(n_9991),
.Y(n_21702)
);

NAND2xp5_ASAP7_75t_L g21703 ( 
.A(n_21618),
.B(n_9991),
.Y(n_21703)
);

XOR2x2_ASAP7_75t_L g21704 ( 
.A(n_21555),
.B(n_9713),
.Y(n_21704)
);

NAND4xp75_ASAP7_75t_L g21705 ( 
.A(n_21557),
.B(n_21633),
.C(n_21583),
.D(n_21602),
.Y(n_21705)
);

INVx2_ASAP7_75t_L g21706 ( 
.A(n_21589),
.Y(n_21706)
);

NAND2x1_ASAP7_75t_L g21707 ( 
.A(n_21574),
.B(n_8675),
.Y(n_21707)
);

NAND4xp75_ASAP7_75t_L g21708 ( 
.A(n_21598),
.B(n_11363),
.C(n_11373),
.D(n_11347),
.Y(n_21708)
);

INVx1_ASAP7_75t_L g21709 ( 
.A(n_21610),
.Y(n_21709)
);

NAND2x1p5_ASAP7_75t_L g21710 ( 
.A(n_21628),
.B(n_8716),
.Y(n_21710)
);

NAND4xp75_ASAP7_75t_L g21711 ( 
.A(n_21558),
.B(n_11363),
.C(n_11373),
.D(n_11347),
.Y(n_21711)
);

AO22x2_ASAP7_75t_L g21712 ( 
.A1(n_21617),
.A2(n_9138),
.B1(n_9151),
.B2(n_9120),
.Y(n_21712)
);

NOR3xp33_ASAP7_75t_L g21713 ( 
.A(n_21561),
.B(n_10300),
.C(n_11262),
.Y(n_21713)
);

NAND2xp5_ASAP7_75t_SL g21714 ( 
.A(n_21548),
.B(n_9222),
.Y(n_21714)
);

OAI222xp33_ASAP7_75t_L g21715 ( 
.A1(n_21575),
.A2(n_9284),
.B1(n_9276),
.B2(n_9286),
.C1(n_9281),
.C2(n_9257),
.Y(n_21715)
);

OR5x1_ASAP7_75t_L g21716 ( 
.A(n_21634),
.B(n_11129),
.C(n_11139),
.D(n_11127),
.E(n_11122),
.Y(n_21716)
);

XNOR2x1_ASAP7_75t_L g21717 ( 
.A(n_21593),
.B(n_8454),
.Y(n_21717)
);

NAND3xp33_ASAP7_75t_L g21718 ( 
.A(n_21579),
.B(n_9281),
.C(n_9276),
.Y(n_21718)
);

INVx1_ASAP7_75t_SL g21719 ( 
.A(n_21634),
.Y(n_21719)
);

INVx2_ASAP7_75t_L g21720 ( 
.A(n_21613),
.Y(n_21720)
);

INVx1_ASAP7_75t_L g21721 ( 
.A(n_21600),
.Y(n_21721)
);

NOR2x1_ASAP7_75t_L g21722 ( 
.A(n_21594),
.B(n_8990),
.Y(n_21722)
);

INVx2_ASAP7_75t_L g21723 ( 
.A(n_21592),
.Y(n_21723)
);

INVxp67_ASAP7_75t_SL g21724 ( 
.A(n_21630),
.Y(n_21724)
);

AND2x4_ASAP7_75t_L g21725 ( 
.A(n_21620),
.B(n_9466),
.Y(n_21725)
);

OAI221xp5_ASAP7_75t_L g21726 ( 
.A1(n_21624),
.A2(n_9286),
.B1(n_9292),
.B2(n_9284),
.C(n_9281),
.Y(n_21726)
);

AND2x4_ASAP7_75t_L g21727 ( 
.A(n_21627),
.B(n_9466),
.Y(n_21727)
);

INVx2_ASAP7_75t_L g21728 ( 
.A(n_21589),
.Y(n_21728)
);

INVx1_ASAP7_75t_L g21729 ( 
.A(n_21552),
.Y(n_21729)
);

NAND2xp5_ASAP7_75t_L g21730 ( 
.A(n_21552),
.B(n_7762),
.Y(n_21730)
);

AND2x2_ASAP7_75t_L g21731 ( 
.A(n_21552),
.B(n_10002),
.Y(n_21731)
);

HB1xp67_ASAP7_75t_L g21732 ( 
.A(n_21573),
.Y(n_21732)
);

NOR4xp25_ASAP7_75t_L g21733 ( 
.A(n_21552),
.B(n_9284),
.C(n_9286),
.D(n_9281),
.Y(n_21733)
);

NOR2xp33_ASAP7_75t_L g21734 ( 
.A(n_21552),
.B(n_10002),
.Y(n_21734)
);

NOR3xp33_ASAP7_75t_SL g21735 ( 
.A(n_21552),
.B(n_9286),
.C(n_9284),
.Y(n_21735)
);

CKINVDCx20_ASAP7_75t_R g21736 ( 
.A(n_21585),
.Y(n_21736)
);

NOR3xp33_ASAP7_75t_L g21737 ( 
.A(n_21665),
.B(n_11255),
.C(n_10300),
.Y(n_21737)
);

NOR3xp33_ASAP7_75t_L g21738 ( 
.A(n_21682),
.B(n_11255),
.C(n_10300),
.Y(n_21738)
);

AOI221xp5_ASAP7_75t_L g21739 ( 
.A1(n_21732),
.A2(n_9305),
.B1(n_9306),
.B2(n_9303),
.C(n_9292),
.Y(n_21739)
);

INVx1_ASAP7_75t_L g21740 ( 
.A(n_21729),
.Y(n_21740)
);

NAND2xp5_ASAP7_75t_L g21741 ( 
.A(n_21667),
.B(n_9251),
.Y(n_21741)
);

AOI22x1_ASAP7_75t_L g21742 ( 
.A1(n_21659),
.A2(n_9151),
.B1(n_9160),
.B2(n_9138),
.Y(n_21742)
);

OAI211xp5_ASAP7_75t_SL g21743 ( 
.A1(n_21645),
.A2(n_9303),
.B(n_9305),
.C(n_9292),
.Y(n_21743)
);

NOR2xp33_ASAP7_75t_L g21744 ( 
.A(n_21667),
.B(n_10103),
.Y(n_21744)
);

OR2x2_ASAP7_75t_L g21745 ( 
.A(n_21672),
.B(n_11122),
.Y(n_21745)
);

NOR3xp33_ASAP7_75t_L g21746 ( 
.A(n_21655),
.B(n_11255),
.C(n_11262),
.Y(n_21746)
);

O2A1O1Ixp33_ASAP7_75t_L g21747 ( 
.A1(n_21648),
.A2(n_21701),
.B(n_21691),
.C(n_21693),
.Y(n_21747)
);

OAI221xp5_ASAP7_75t_L g21748 ( 
.A1(n_21644),
.A2(n_9305),
.B1(n_9306),
.B2(n_9303),
.C(n_9292),
.Y(n_21748)
);

INVxp67_ASAP7_75t_L g21749 ( 
.A(n_21675),
.Y(n_21749)
);

AOI21xp5_ASAP7_75t_L g21750 ( 
.A1(n_21724),
.A2(n_10103),
.B(n_11519),
.Y(n_21750)
);

AND2x2_ASAP7_75t_L g21751 ( 
.A(n_21667),
.B(n_10103),
.Y(n_21751)
);

OAI21xp5_ASAP7_75t_SL g21752 ( 
.A1(n_21721),
.A2(n_9241),
.B(n_9217),
.Y(n_21752)
);

INVx1_ASAP7_75t_L g21753 ( 
.A(n_21736),
.Y(n_21753)
);

AND2x4_ASAP7_75t_L g21754 ( 
.A(n_21731),
.B(n_9466),
.Y(n_21754)
);

NOR2xp67_ASAP7_75t_L g21755 ( 
.A(n_21640),
.B(n_8202),
.Y(n_21755)
);

NAND3xp33_ASAP7_75t_L g21756 ( 
.A(n_21640),
.B(n_9305),
.C(n_9303),
.Y(n_21756)
);

NAND2xp5_ASAP7_75t_SL g21757 ( 
.A(n_21640),
.B(n_9241),
.Y(n_21757)
);

CKINVDCx20_ASAP7_75t_R g21758 ( 
.A(n_21723),
.Y(n_21758)
);

AO22x2_ASAP7_75t_L g21759 ( 
.A1(n_21706),
.A2(n_9138),
.B1(n_9160),
.B2(n_9151),
.Y(n_21759)
);

OAI21xp5_ASAP7_75t_SL g21760 ( 
.A1(n_21720),
.A2(n_9265),
.B(n_9241),
.Y(n_21760)
);

AOI22xp33_ASAP7_75t_SL g21761 ( 
.A1(n_21728),
.A2(n_11525),
.B1(n_11528),
.B2(n_11519),
.Y(n_21761)
);

NAND2xp5_ASAP7_75t_L g21762 ( 
.A(n_21734),
.B(n_9251),
.Y(n_21762)
);

NAND4xp25_ASAP7_75t_L g21763 ( 
.A(n_21709),
.B(n_9129),
.C(n_8949),
.D(n_8959),
.Y(n_21763)
);

AOI31xp33_ASAP7_75t_L g21764 ( 
.A1(n_21684),
.A2(n_7999),
.A3(n_8000),
.B(n_7995),
.Y(n_21764)
);

AOI221xp5_ASAP7_75t_L g21765 ( 
.A1(n_21643),
.A2(n_9309),
.B1(n_9313),
.B2(n_9307),
.C(n_9306),
.Y(n_21765)
);

NOR3xp33_ASAP7_75t_L g21766 ( 
.A(n_21719),
.B(n_21705),
.C(n_21730),
.Y(n_21766)
);

AND4x1_ASAP7_75t_L g21767 ( 
.A(n_21685),
.B(n_8966),
.C(n_8892),
.D(n_9852),
.Y(n_21767)
);

NOR3x1_ASAP7_75t_L g21768 ( 
.A(n_21669),
.B(n_11127),
.C(n_11122),
.Y(n_21768)
);

INVx4_ASAP7_75t_L g21769 ( 
.A(n_21692),
.Y(n_21769)
);

AOI221xp5_ASAP7_75t_L g21770 ( 
.A1(n_21646),
.A2(n_9309),
.B1(n_9313),
.B2(n_9307),
.C(n_9306),
.Y(n_21770)
);

BUFx6f_ASAP7_75t_L g21771 ( 
.A(n_21707),
.Y(n_21771)
);

NAND2xp5_ASAP7_75t_L g21772 ( 
.A(n_21679),
.B(n_9251),
.Y(n_21772)
);

AND3x4_ASAP7_75t_L g21773 ( 
.A(n_21641),
.B(n_21650),
.C(n_21642),
.Y(n_21773)
);

NOR3xp33_ASAP7_75t_L g21774 ( 
.A(n_21703),
.B(n_11267),
.C(n_11262),
.Y(n_21774)
);

NAND4xp75_ASAP7_75t_L g21775 ( 
.A(n_21663),
.B(n_11363),
.C(n_11373),
.D(n_11347),
.Y(n_21775)
);

OR2x2_ASAP7_75t_L g21776 ( 
.A(n_21710),
.B(n_21717),
.Y(n_21776)
);

NOR3xp33_ASAP7_75t_L g21777 ( 
.A(n_21658),
.B(n_21651),
.C(n_21714),
.Y(n_21777)
);

INVx1_ASAP7_75t_L g21778 ( 
.A(n_21704),
.Y(n_21778)
);

NOR3xp33_ASAP7_75t_L g21779 ( 
.A(n_21702),
.B(n_11270),
.C(n_11267),
.Y(n_21779)
);

OR2x2_ASAP7_75t_L g21780 ( 
.A(n_21666),
.B(n_11127),
.Y(n_21780)
);

OAI21xp5_ASAP7_75t_SL g21781 ( 
.A1(n_21678),
.A2(n_9265),
.B(n_9241),
.Y(n_21781)
);

INVx1_ASAP7_75t_L g21782 ( 
.A(n_21700),
.Y(n_21782)
);

NOR2x1_ASAP7_75t_L g21783 ( 
.A(n_21653),
.B(n_8990),
.Y(n_21783)
);

NAND2xp5_ASAP7_75t_L g21784 ( 
.A(n_21727),
.B(n_9251),
.Y(n_21784)
);

OAI322xp33_ASAP7_75t_L g21785 ( 
.A1(n_21696),
.A2(n_9322),
.A3(n_9313),
.B1(n_9324),
.B2(n_9338),
.C1(n_9317),
.C2(n_9307),
.Y(n_21785)
);

NAND2xp5_ASAP7_75t_L g21786 ( 
.A(n_21688),
.B(n_9251),
.Y(n_21786)
);

OR2x2_ASAP7_75t_L g21787 ( 
.A(n_21697),
.B(n_11129),
.Y(n_21787)
);

NAND2xp5_ASAP7_75t_L g21788 ( 
.A(n_21725),
.B(n_21671),
.Y(n_21788)
);

O2A1O1Ixp33_ASAP7_75t_L g21789 ( 
.A1(n_21694),
.A2(n_10103),
.B(n_9151),
.C(n_9160),
.Y(n_21789)
);

AND2x4_ASAP7_75t_L g21790 ( 
.A(n_21683),
.B(n_9466),
.Y(n_21790)
);

AOI21xp5_ASAP7_75t_L g21791 ( 
.A1(n_21654),
.A2(n_10103),
.B(n_11519),
.Y(n_21791)
);

AOI221xp5_ASAP7_75t_L g21792 ( 
.A1(n_21699),
.A2(n_9322),
.B1(n_9324),
.B2(n_9317),
.C(n_9313),
.Y(n_21792)
);

OAI22xp5_ASAP7_75t_L g21793 ( 
.A1(n_21661),
.A2(n_9322),
.B1(n_9324),
.B2(n_9317),
.Y(n_21793)
);

AOI21xp5_ASAP7_75t_L g21794 ( 
.A1(n_21722),
.A2(n_10103),
.B(n_11525),
.Y(n_21794)
);

NOR2x1_ASAP7_75t_L g21795 ( 
.A(n_21718),
.B(n_21670),
.Y(n_21795)
);

NAND2xp5_ASAP7_75t_L g21796 ( 
.A(n_21668),
.B(n_9251),
.Y(n_21796)
);

OAI221xp5_ASAP7_75t_L g21797 ( 
.A1(n_21735),
.A2(n_9338),
.B1(n_9340),
.B2(n_9324),
.C(n_9322),
.Y(n_21797)
);

AND2x4_ASAP7_75t_L g21798 ( 
.A(n_21687),
.B(n_9466),
.Y(n_21798)
);

BUFx6f_ASAP7_75t_L g21799 ( 
.A(n_21698),
.Y(n_21799)
);

NAND3xp33_ASAP7_75t_SL g21800 ( 
.A(n_21676),
.B(n_8000),
.C(n_7995),
.Y(n_21800)
);

NAND3x1_ASAP7_75t_SL g21801 ( 
.A(n_21649),
.B(n_21656),
.C(n_21662),
.Y(n_21801)
);

AOI21xp5_ASAP7_75t_L g21802 ( 
.A1(n_21686),
.A2(n_11528),
.B(n_11525),
.Y(n_21802)
);

AND2x2_ASAP7_75t_L g21803 ( 
.A(n_21713),
.B(n_11528),
.Y(n_21803)
);

OAI22xp5_ASAP7_75t_L g21804 ( 
.A1(n_21712),
.A2(n_9340),
.B1(n_9342),
.B2(n_9338),
.Y(n_21804)
);

INVx1_ASAP7_75t_L g21805 ( 
.A(n_21712),
.Y(n_21805)
);

AND2x2_ASAP7_75t_L g21806 ( 
.A(n_21690),
.B(n_11531),
.Y(n_21806)
);

OR2x2_ASAP7_75t_L g21807 ( 
.A(n_21733),
.B(n_11129),
.Y(n_21807)
);

NOR2x1_ASAP7_75t_L g21808 ( 
.A(n_21708),
.B(n_8990),
.Y(n_21808)
);

AO211x2_ASAP7_75t_L g21809 ( 
.A1(n_21677),
.A2(n_9338),
.B(n_9342),
.C(n_9340),
.Y(n_21809)
);

NOR4xp75_ASAP7_75t_L g21810 ( 
.A(n_21711),
.B(n_8036),
.C(n_8039),
.D(n_8026),
.Y(n_21810)
);

NAND3xp33_ASAP7_75t_L g21811 ( 
.A(n_21652),
.B(n_9342),
.C(n_9340),
.Y(n_21811)
);

AOI222xp33_ASAP7_75t_L g21812 ( 
.A1(n_21726),
.A2(n_9311),
.B1(n_9241),
.B2(n_9326),
.C1(n_9312),
.C2(n_9265),
.Y(n_21812)
);

NOR3xp33_ASAP7_75t_L g21813 ( 
.A(n_21657),
.B(n_11270),
.C(n_11267),
.Y(n_21813)
);

NOR2x1p5_ASAP7_75t_L g21814 ( 
.A(n_21664),
.B(n_8814),
.Y(n_21814)
);

AND4x1_ASAP7_75t_L g21815 ( 
.A(n_21747),
.B(n_21674),
.C(n_21673),
.D(n_21647),
.Y(n_21815)
);

AND2x2_ASAP7_75t_L g21816 ( 
.A(n_21751),
.B(n_21681),
.Y(n_21816)
);

INVx1_ASAP7_75t_L g21817 ( 
.A(n_21740),
.Y(n_21817)
);

AND2x4_ASAP7_75t_L g21818 ( 
.A(n_21757),
.B(n_21695),
.Y(n_21818)
);

INVx1_ASAP7_75t_L g21819 ( 
.A(n_21753),
.Y(n_21819)
);

INVx3_ASAP7_75t_L g21820 ( 
.A(n_21769),
.Y(n_21820)
);

INVx2_ASAP7_75t_SL g21821 ( 
.A(n_21771),
.Y(n_21821)
);

INVx1_ASAP7_75t_L g21822 ( 
.A(n_21758),
.Y(n_21822)
);

XNOR2x1_ASAP7_75t_L g21823 ( 
.A(n_21773),
.B(n_21660),
.Y(n_21823)
);

NOR2x1_ASAP7_75t_L g21824 ( 
.A(n_21771),
.B(n_21715),
.Y(n_21824)
);

NAND2x1p5_ASAP7_75t_L g21825 ( 
.A(n_21782),
.B(n_21689),
.Y(n_21825)
);

AND2x4_ASAP7_75t_L g21826 ( 
.A(n_21741),
.B(n_21716),
.Y(n_21826)
);

BUFx3_ASAP7_75t_L g21827 ( 
.A(n_21788),
.Y(n_21827)
);

NOR2xp33_ASAP7_75t_L g21828 ( 
.A(n_21749),
.B(n_21680),
.Y(n_21828)
);

INVx1_ASAP7_75t_L g21829 ( 
.A(n_21776),
.Y(n_21829)
);

NOR2x1p5_ASAP7_75t_L g21830 ( 
.A(n_21799),
.B(n_8814),
.Y(n_21830)
);

INVx2_ASAP7_75t_L g21831 ( 
.A(n_21799),
.Y(n_21831)
);

NAND2xp5_ASAP7_75t_L g21832 ( 
.A(n_21744),
.B(n_9251),
.Y(n_21832)
);

NOR3xp33_ASAP7_75t_L g21833 ( 
.A(n_21766),
.B(n_11056),
.C(n_11054),
.Y(n_21833)
);

NOR2xp33_ASAP7_75t_L g21834 ( 
.A(n_21778),
.B(n_21795),
.Y(n_21834)
);

INVx2_ASAP7_75t_L g21835 ( 
.A(n_21814),
.Y(n_21835)
);

INVx2_ASAP7_75t_L g21836 ( 
.A(n_21805),
.Y(n_21836)
);

XOR2xp5_ASAP7_75t_L g21837 ( 
.A(n_21762),
.B(n_8454),
.Y(n_21837)
);

NOR2x1_ASAP7_75t_L g21838 ( 
.A(n_21808),
.B(n_8990),
.Y(n_21838)
);

AOI21x1_ASAP7_75t_L g21839 ( 
.A1(n_21794),
.A2(n_9034),
.B(n_9021),
.Y(n_21839)
);

INVx1_ASAP7_75t_L g21840 ( 
.A(n_21801),
.Y(n_21840)
);

NAND5xp2_ASAP7_75t_L g21841 ( 
.A(n_21777),
.B(n_8966),
.C(n_8914),
.D(n_8895),
.E(n_9021),
.Y(n_21841)
);

INVx2_ASAP7_75t_L g21842 ( 
.A(n_21798),
.Y(n_21842)
);

XNOR2xp5_ASAP7_75t_L g21843 ( 
.A(n_21810),
.B(n_8860),
.Y(n_21843)
);

NAND4xp75_ASAP7_75t_L g21844 ( 
.A(n_21755),
.B(n_11363),
.C(n_11373),
.D(n_11347),
.Y(n_21844)
);

INVx2_ASAP7_75t_L g21845 ( 
.A(n_21790),
.Y(n_21845)
);

NAND2xp5_ASAP7_75t_L g21846 ( 
.A(n_21754),
.B(n_9251),
.Y(n_21846)
);

BUFx2_ASAP7_75t_L g21847 ( 
.A(n_21784),
.Y(n_21847)
);

XNOR2xp5_ASAP7_75t_L g21848 ( 
.A(n_21772),
.B(n_21786),
.Y(n_21848)
);

OAI22xp33_ASAP7_75t_R g21849 ( 
.A1(n_21787),
.A2(n_8212),
.B1(n_8284),
.B2(n_8202),
.Y(n_21849)
);

INVx1_ASAP7_75t_L g21850 ( 
.A(n_21796),
.Y(n_21850)
);

INVx3_ASAP7_75t_L g21851 ( 
.A(n_21780),
.Y(n_21851)
);

XOR2x1_ASAP7_75t_L g21852 ( 
.A(n_21809),
.B(n_9241),
.Y(n_21852)
);

INVx3_ASAP7_75t_L g21853 ( 
.A(n_21745),
.Y(n_21853)
);

OAI21x1_ASAP7_75t_L g21854 ( 
.A1(n_21783),
.A2(n_7907),
.B(n_8983),
.Y(n_21854)
);

AOI22xp5_ASAP7_75t_L g21855 ( 
.A1(n_21760),
.A2(n_9241),
.B1(n_9311),
.B2(n_9265),
.Y(n_21855)
);

NAND2x1p5_ASAP7_75t_L g21856 ( 
.A(n_21791),
.B(n_8740),
.Y(n_21856)
);

NOR3xp33_ASAP7_75t_SL g21857 ( 
.A(n_21752),
.B(n_8036),
.C(n_8026),
.Y(n_21857)
);

INVx2_ASAP7_75t_L g21858 ( 
.A(n_21807),
.Y(n_21858)
);

INVx1_ASAP7_75t_L g21859 ( 
.A(n_21764),
.Y(n_21859)
);

INVx1_ASAP7_75t_L g21860 ( 
.A(n_21806),
.Y(n_21860)
);

OR3x2_ASAP7_75t_L g21861 ( 
.A(n_21763),
.B(n_9383),
.C(n_9363),
.Y(n_21861)
);

AND2x2_ASAP7_75t_L g21862 ( 
.A(n_21803),
.B(n_11531),
.Y(n_21862)
);

OR2x2_ASAP7_75t_L g21863 ( 
.A(n_21800),
.B(n_11171),
.Y(n_21863)
);

INVx1_ASAP7_75t_L g21864 ( 
.A(n_21756),
.Y(n_21864)
);

NAND2xp33_ASAP7_75t_L g21865 ( 
.A(n_21813),
.B(n_9835),
.Y(n_21865)
);

INVxp67_ASAP7_75t_SL g21866 ( 
.A(n_21789),
.Y(n_21866)
);

INVx2_ASAP7_75t_L g21867 ( 
.A(n_21775),
.Y(n_21867)
);

AND3x4_ASAP7_75t_L g21868 ( 
.A(n_21779),
.B(n_8744),
.C(n_8740),
.Y(n_21868)
);

OAI22xp5_ASAP7_75t_L g21869 ( 
.A1(n_21797),
.A2(n_9352),
.B1(n_9357),
.B2(n_9342),
.Y(n_21869)
);

NOR2x1_ASAP7_75t_L g21870 ( 
.A(n_21743),
.B(n_8999),
.Y(n_21870)
);

OAI22xp33_ASAP7_75t_L g21871 ( 
.A1(n_21781),
.A2(n_21793),
.B1(n_21750),
.B2(n_21770),
.Y(n_21871)
);

OAI22x1_ASAP7_75t_L g21872 ( 
.A1(n_21767),
.A2(n_9160),
.B1(n_9166),
.B2(n_9138),
.Y(n_21872)
);

NOR2x1_ASAP7_75t_L g21873 ( 
.A(n_21811),
.B(n_8999),
.Y(n_21873)
);

OAI22xp5_ASAP7_75t_L g21874 ( 
.A1(n_21817),
.A2(n_21738),
.B1(n_21748),
.B2(n_21737),
.Y(n_21874)
);

AOI221xp5_ASAP7_75t_L g21875 ( 
.A1(n_21871),
.A2(n_21804),
.B1(n_21774),
.B2(n_21792),
.C(n_21802),
.Y(n_21875)
);

AOI322xp5_ASAP7_75t_L g21876 ( 
.A1(n_21840),
.A2(n_21765),
.A3(n_21739),
.B1(n_21746),
.B2(n_21761),
.C1(n_21768),
.C2(n_21742),
.Y(n_21876)
);

OAI211xp5_ASAP7_75t_L g21877 ( 
.A1(n_21822),
.A2(n_21812),
.B(n_21759),
.C(n_21785),
.Y(n_21877)
);

OAI22xp5_ASAP7_75t_SL g21878 ( 
.A1(n_21819),
.A2(n_21759),
.B1(n_8878),
.B2(n_8675),
.Y(n_21878)
);

NOR3xp33_ASAP7_75t_L g21879 ( 
.A(n_21820),
.B(n_8983),
.C(n_11072),
.Y(n_21879)
);

OAI322xp33_ASAP7_75t_L g21880 ( 
.A1(n_21836),
.A2(n_9363),
.A3(n_9357),
.B1(n_9371),
.B2(n_9375),
.C1(n_9360),
.C2(n_9352),
.Y(n_21880)
);

NOR2x1p5_ASAP7_75t_L g21881 ( 
.A(n_21827),
.B(n_8814),
.Y(n_21881)
);

INVx1_ASAP7_75t_L g21882 ( 
.A(n_21842),
.Y(n_21882)
);

AOI322xp5_ASAP7_75t_L g21883 ( 
.A1(n_21821),
.A2(n_9363),
.A3(n_9357),
.B1(n_9371),
.B2(n_9375),
.C1(n_9360),
.C2(n_9352),
.Y(n_21883)
);

OAI211xp5_ASAP7_75t_SL g21884 ( 
.A1(n_21829),
.A2(n_9352),
.B(n_9363),
.C(n_9360),
.Y(n_21884)
);

NAND4xp75_ASAP7_75t_L g21885 ( 
.A(n_21824),
.B(n_11482),
.C(n_11500),
.D(n_11434),
.Y(n_21885)
);

OAI221xp5_ASAP7_75t_L g21886 ( 
.A1(n_21815),
.A2(n_9516),
.B1(n_9527),
.B2(n_9500),
.C(n_9480),
.Y(n_21886)
);

OAI211xp5_ASAP7_75t_L g21887 ( 
.A1(n_21828),
.A2(n_9375),
.B(n_9383),
.C(n_9371),
.Y(n_21887)
);

INVx1_ASAP7_75t_L g21888 ( 
.A(n_21816),
.Y(n_21888)
);

INVx1_ASAP7_75t_L g21889 ( 
.A(n_21818),
.Y(n_21889)
);

OAI22xp33_ASAP7_75t_SL g21890 ( 
.A1(n_21825),
.A2(n_8878),
.B1(n_8675),
.B2(n_9371),
.Y(n_21890)
);

AOI22x1_ASAP7_75t_L g21891 ( 
.A1(n_21831),
.A2(n_9166),
.B1(n_9170),
.B2(n_9160),
.Y(n_21891)
);

AOI322xp5_ASAP7_75t_L g21892 ( 
.A1(n_21834),
.A2(n_9410),
.A3(n_9383),
.B1(n_9420),
.B2(n_9421),
.C1(n_9405),
.C2(n_9375),
.Y(n_21892)
);

XNOR2xp5_ASAP7_75t_L g21893 ( 
.A(n_21823),
.B(n_8860),
.Y(n_21893)
);

INVx2_ASAP7_75t_L g21894 ( 
.A(n_21835),
.Y(n_21894)
);

OAI211xp5_ASAP7_75t_SL g21895 ( 
.A1(n_21860),
.A2(n_9383),
.B(n_9410),
.C(n_9405),
.Y(n_21895)
);

OAI211xp5_ASAP7_75t_SL g21896 ( 
.A1(n_21853),
.A2(n_9405),
.B(n_9420),
.C(n_9410),
.Y(n_21896)
);

INVx1_ASAP7_75t_L g21897 ( 
.A(n_21858),
.Y(n_21897)
);

AOI221xp5_ASAP7_75t_L g21898 ( 
.A1(n_21864),
.A2(n_9429),
.B1(n_9430),
.B2(n_9420),
.C(n_9405),
.Y(n_21898)
);

AOI322xp5_ASAP7_75t_L g21899 ( 
.A1(n_21845),
.A2(n_9430),
.A3(n_9421),
.B1(n_9436),
.B2(n_9438),
.C1(n_9429),
.C2(n_9420),
.Y(n_21899)
);

AOI322xp5_ASAP7_75t_L g21900 ( 
.A1(n_21865),
.A2(n_9436),
.A3(n_9429),
.B1(n_9438),
.B2(n_9450),
.C1(n_9430),
.C2(n_9421),
.Y(n_21900)
);

OAI221xp5_ASAP7_75t_SL g21901 ( 
.A1(n_21859),
.A2(n_21866),
.B1(n_21867),
.B2(n_21850),
.C(n_21848),
.Y(n_21901)
);

OAI322xp33_ASAP7_75t_L g21902 ( 
.A1(n_21851),
.A2(n_9436),
.A3(n_9429),
.B1(n_9438),
.B2(n_9450),
.C1(n_9430),
.C2(n_9421),
.Y(n_21902)
);

OAI322xp33_ASAP7_75t_L g21903 ( 
.A1(n_21847),
.A2(n_21856),
.A3(n_21832),
.B1(n_21863),
.B2(n_21846),
.C1(n_21869),
.C2(n_21843),
.Y(n_21903)
);

AOI322xp5_ASAP7_75t_L g21904 ( 
.A1(n_21826),
.A2(n_9463),
.A3(n_9438),
.B1(n_9465),
.B2(n_9479),
.C1(n_9450),
.C2(n_9436),
.Y(n_21904)
);

AOI322xp5_ASAP7_75t_L g21905 ( 
.A1(n_21838),
.A2(n_9479),
.A3(n_9463),
.B1(n_9480),
.B2(n_9481),
.C1(n_9465),
.C2(n_9450),
.Y(n_21905)
);

AOI322xp5_ASAP7_75t_L g21906 ( 
.A1(n_21873),
.A2(n_9480),
.A3(n_9465),
.B1(n_9481),
.B2(n_9483),
.C1(n_9479),
.C2(n_9463),
.Y(n_21906)
);

AOI322xp5_ASAP7_75t_L g21907 ( 
.A1(n_21857),
.A2(n_9483),
.A3(n_9479),
.B1(n_9491),
.B2(n_9494),
.C1(n_9481),
.C2(n_9465),
.Y(n_21907)
);

AOI32xp33_ASAP7_75t_L g21908 ( 
.A1(n_21862),
.A2(n_11551),
.A3(n_11552),
.B1(n_11542),
.B2(n_11531),
.Y(n_21908)
);

OAI221xp5_ASAP7_75t_L g21909 ( 
.A1(n_21870),
.A2(n_9527),
.B1(n_9516),
.B2(n_9500),
.C(n_9491),
.Y(n_21909)
);

AOI22xp5_ASAP7_75t_L g21910 ( 
.A1(n_21830),
.A2(n_9265),
.B1(n_9312),
.B2(n_9311),
.Y(n_21910)
);

AOI32xp33_ASAP7_75t_L g21911 ( 
.A1(n_21852),
.A2(n_11552),
.A3(n_11553),
.B1(n_11551),
.B2(n_11542),
.Y(n_21911)
);

INVx1_ASAP7_75t_L g21912 ( 
.A(n_21861),
.Y(n_21912)
);

NOR2x1p5_ASAP7_75t_L g21913 ( 
.A(n_21839),
.B(n_21868),
.Y(n_21913)
);

AOI322xp5_ASAP7_75t_L g21914 ( 
.A1(n_21833),
.A2(n_9494),
.A3(n_9483),
.B1(n_9500),
.B2(n_9516),
.C1(n_9491),
.C2(n_9481),
.Y(n_21914)
);

NOR3xp33_ASAP7_75t_L g21915 ( 
.A(n_21841),
.B(n_21844),
.C(n_21854),
.Y(n_21915)
);

INVx4_ASAP7_75t_L g21916 ( 
.A(n_21894),
.Y(n_21916)
);

INVx1_ASAP7_75t_L g21917 ( 
.A(n_21882),
.Y(n_21917)
);

HB1xp67_ASAP7_75t_L g21918 ( 
.A(n_21888),
.Y(n_21918)
);

XNOR2x1_ASAP7_75t_L g21919 ( 
.A(n_21889),
.B(n_21872),
.Y(n_21919)
);

XNOR2x1_ASAP7_75t_L g21920 ( 
.A(n_21913),
.B(n_21897),
.Y(n_21920)
);

XOR2xp5_ASAP7_75t_L g21921 ( 
.A(n_21893),
.B(n_21837),
.Y(n_21921)
);

XOR2xp5_ASAP7_75t_L g21922 ( 
.A(n_21874),
.B(n_21855),
.Y(n_21922)
);

XNOR2xp5_ASAP7_75t_L g21923 ( 
.A(n_21877),
.B(n_21849),
.Y(n_21923)
);

AND2x4_ASAP7_75t_L g21924 ( 
.A(n_21915),
.B(n_9466),
.Y(n_21924)
);

O2A1O1Ixp33_ASAP7_75t_SL g21925 ( 
.A1(n_21912),
.A2(n_9491),
.B(n_9494),
.C(n_9483),
.Y(n_21925)
);

AOI22xp33_ASAP7_75t_SL g21926 ( 
.A1(n_21878),
.A2(n_11542),
.B1(n_11552),
.B2(n_11551),
.Y(n_21926)
);

AOI22x1_ASAP7_75t_L g21927 ( 
.A1(n_21901),
.A2(n_9166),
.B1(n_9170),
.B2(n_9160),
.Y(n_21927)
);

NAND2xp5_ASAP7_75t_L g21928 ( 
.A(n_21876),
.B(n_9251),
.Y(n_21928)
);

NOR2x1p5_ASAP7_75t_L g21929 ( 
.A(n_21903),
.B(n_8039),
.Y(n_21929)
);

OAI22xp5_ASAP7_75t_SL g21930 ( 
.A1(n_21875),
.A2(n_8878),
.B1(n_8675),
.B2(n_9123),
.Y(n_21930)
);

NOR3xp33_ASAP7_75t_L g21931 ( 
.A(n_21909),
.B(n_8983),
.C(n_11095),
.Y(n_21931)
);

INVx2_ASAP7_75t_SL g21932 ( 
.A(n_21881),
.Y(n_21932)
);

INVx1_ASAP7_75t_L g21933 ( 
.A(n_21885),
.Y(n_21933)
);

OAI22xp5_ASAP7_75t_L g21934 ( 
.A1(n_21887),
.A2(n_21910),
.B1(n_21886),
.B2(n_21911),
.Y(n_21934)
);

INVx2_ASAP7_75t_L g21935 ( 
.A(n_21891),
.Y(n_21935)
);

OAI21xp5_ASAP7_75t_L g21936 ( 
.A1(n_21884),
.A2(n_21895),
.B(n_21896),
.Y(n_21936)
);

NAND2xp5_ASAP7_75t_L g21937 ( 
.A(n_21900),
.B(n_9251),
.Y(n_21937)
);

AOI22xp5_ASAP7_75t_L g21938 ( 
.A1(n_21890),
.A2(n_9265),
.B1(n_9312),
.B2(n_9311),
.Y(n_21938)
);

NOR2x1_ASAP7_75t_L g21939 ( 
.A(n_21880),
.B(n_8999),
.Y(n_21939)
);

INVx2_ASAP7_75t_L g21940 ( 
.A(n_21906),
.Y(n_21940)
);

INVx1_ASAP7_75t_L g21941 ( 
.A(n_21879),
.Y(n_21941)
);

OAI22xp5_ASAP7_75t_SL g21942 ( 
.A1(n_21907),
.A2(n_21914),
.B1(n_21904),
.B2(n_21905),
.Y(n_21942)
);

INVx2_ASAP7_75t_L g21943 ( 
.A(n_21916),
.Y(n_21943)
);

OAI22xp33_ASAP7_75t_L g21944 ( 
.A1(n_21917),
.A2(n_21898),
.B1(n_21892),
.B2(n_21902),
.Y(n_21944)
);

INVx3_ASAP7_75t_SL g21945 ( 
.A(n_21919),
.Y(n_21945)
);

INVxp67_ASAP7_75t_L g21946 ( 
.A(n_21918),
.Y(n_21946)
);

INVx2_ASAP7_75t_L g21947 ( 
.A(n_21920),
.Y(n_21947)
);

INVx1_ASAP7_75t_L g21948 ( 
.A(n_21923),
.Y(n_21948)
);

INVx1_ASAP7_75t_L g21949 ( 
.A(n_21929),
.Y(n_21949)
);

INVx2_ASAP7_75t_L g21950 ( 
.A(n_21935),
.Y(n_21950)
);

INVx2_ASAP7_75t_L g21951 ( 
.A(n_21932),
.Y(n_21951)
);

XNOR2xp5_ASAP7_75t_L g21952 ( 
.A(n_21921),
.B(n_21908),
.Y(n_21952)
);

AOI22x1_ASAP7_75t_L g21953 ( 
.A1(n_21922),
.A2(n_21899),
.B1(n_21883),
.B2(n_9170),
.Y(n_21953)
);

OAI22xp5_ASAP7_75t_SL g21954 ( 
.A1(n_21940),
.A2(n_8878),
.B1(n_8675),
.B2(n_8284),
.Y(n_21954)
);

INVx1_ASAP7_75t_L g21955 ( 
.A(n_21933),
.Y(n_21955)
);

AND3x4_ASAP7_75t_L g21956 ( 
.A(n_21924),
.B(n_8744),
.C(n_8740),
.Y(n_21956)
);

XNOR2xp5_ASAP7_75t_L g21957 ( 
.A(n_21928),
.B(n_8744),
.Y(n_21957)
);

NOR2xp67_ASAP7_75t_L g21958 ( 
.A(n_21941),
.B(n_8744),
.Y(n_21958)
);

AO21x1_ASAP7_75t_L g21959 ( 
.A1(n_21934),
.A2(n_11140),
.B(n_11139),
.Y(n_21959)
);

INVx1_ASAP7_75t_L g21960 ( 
.A(n_21942),
.Y(n_21960)
);

XNOR2x1_ASAP7_75t_L g21961 ( 
.A(n_21936),
.B(n_8744),
.Y(n_21961)
);

INVx2_ASAP7_75t_L g21962 ( 
.A(n_21939),
.Y(n_21962)
);

XNOR2x1_ASAP7_75t_L g21963 ( 
.A(n_21937),
.B(n_8744),
.Y(n_21963)
);

INVx1_ASAP7_75t_L g21964 ( 
.A(n_21931),
.Y(n_21964)
);

OAI22xp5_ASAP7_75t_L g21965 ( 
.A1(n_21946),
.A2(n_21960),
.B1(n_21945),
.B2(n_21947),
.Y(n_21965)
);

OAI22xp5_ASAP7_75t_L g21966 ( 
.A1(n_21943),
.A2(n_21927),
.B1(n_21938),
.B2(n_21926),
.Y(n_21966)
);

XNOR2xp5_ASAP7_75t_L g21967 ( 
.A(n_21952),
.B(n_21930),
.Y(n_21967)
);

INVx1_ASAP7_75t_L g21968 ( 
.A(n_21951),
.Y(n_21968)
);

INVx1_ASAP7_75t_L g21969 ( 
.A(n_21950),
.Y(n_21969)
);

OAI22xp5_ASAP7_75t_L g21970 ( 
.A1(n_21948),
.A2(n_21925),
.B1(n_9170),
.B2(n_9270),
.Y(n_21970)
);

AOI22xp5_ASAP7_75t_L g21971 ( 
.A1(n_21955),
.A2(n_9265),
.B1(n_9312),
.B2(n_9311),
.Y(n_21971)
);

NAND2xp5_ASAP7_75t_L g21972 ( 
.A(n_21949),
.B(n_9251),
.Y(n_21972)
);

NAND3xp33_ASAP7_75t_L g21973 ( 
.A(n_21964),
.B(n_9500),
.C(n_9494),
.Y(n_21973)
);

OAI22xp33_ASAP7_75t_L g21974 ( 
.A1(n_21962),
.A2(n_9521),
.B1(n_9525),
.B2(n_9516),
.Y(n_21974)
);

INVx1_ASAP7_75t_L g21975 ( 
.A(n_21944),
.Y(n_21975)
);

AO21x2_ASAP7_75t_L g21976 ( 
.A1(n_21958),
.A2(n_8049),
.B(n_8043),
.Y(n_21976)
);

AOI21xp5_ASAP7_75t_L g21977 ( 
.A1(n_21965),
.A2(n_21961),
.B(n_21957),
.Y(n_21977)
);

OAI21x1_ASAP7_75t_SL g21978 ( 
.A1(n_21967),
.A2(n_21953),
.B(n_21963),
.Y(n_21978)
);

INVx1_ASAP7_75t_L g21979 ( 
.A(n_21968),
.Y(n_21979)
);

NAND2xp5_ASAP7_75t_L g21980 ( 
.A(n_21969),
.B(n_21975),
.Y(n_21980)
);

INVx1_ASAP7_75t_L g21981 ( 
.A(n_21966),
.Y(n_21981)
);

OAI21xp5_ASAP7_75t_L g21982 ( 
.A1(n_21972),
.A2(n_21956),
.B(n_21954),
.Y(n_21982)
);

AOI21xp5_ASAP7_75t_L g21983 ( 
.A1(n_21970),
.A2(n_21959),
.B(n_8049),
.Y(n_21983)
);

INVx1_ASAP7_75t_L g21984 ( 
.A(n_21976),
.Y(n_21984)
);

OA21x2_ASAP7_75t_L g21985 ( 
.A1(n_21973),
.A2(n_11140),
.B(n_11139),
.Y(n_21985)
);

NOR2x1_ASAP7_75t_L g21986 ( 
.A(n_21980),
.B(n_21974),
.Y(n_21986)
);

AOI22xp5_ASAP7_75t_L g21987 ( 
.A1(n_21979),
.A2(n_21971),
.B1(n_9312),
.B2(n_9326),
.Y(n_21987)
);

OAI22xp5_ASAP7_75t_L g21988 ( 
.A1(n_21981),
.A2(n_9170),
.B1(n_9270),
.B2(n_9166),
.Y(n_21988)
);

OAI22xp5_ASAP7_75t_L g21989 ( 
.A1(n_21977),
.A2(n_9170),
.B1(n_9270),
.B2(n_9166),
.Y(n_21989)
);

OAI22xp5_ASAP7_75t_L g21990 ( 
.A1(n_21984),
.A2(n_9270),
.B1(n_9274),
.B2(n_9166),
.Y(n_21990)
);

OAI22xp5_ASAP7_75t_L g21991 ( 
.A1(n_21982),
.A2(n_9274),
.B1(n_9278),
.B2(n_9270),
.Y(n_21991)
);

AOI22xp5_ASAP7_75t_L g21992 ( 
.A1(n_21986),
.A2(n_21983),
.B1(n_21978),
.B2(n_21985),
.Y(n_21992)
);

NAND2xp5_ASAP7_75t_L g21993 ( 
.A(n_21987),
.B(n_9251),
.Y(n_21993)
);

OAI22xp5_ASAP7_75t_L g21994 ( 
.A1(n_21991),
.A2(n_9270),
.B1(n_9278),
.B2(n_9274),
.Y(n_21994)
);

XOR2x2_ASAP7_75t_L g21995 ( 
.A(n_21989),
.B(n_8914),
.Y(n_21995)
);

AOI21xp5_ASAP7_75t_L g21996 ( 
.A1(n_21992),
.A2(n_21988),
.B(n_21990),
.Y(n_21996)
);

OAI21xp5_ASAP7_75t_L g21997 ( 
.A1(n_21993),
.A2(n_11145),
.B(n_11140),
.Y(n_21997)
);

AOI21xp5_ASAP7_75t_L g21998 ( 
.A1(n_21995),
.A2(n_21994),
.B(n_8051),
.Y(n_21998)
);

AOI21xp5_ASAP7_75t_L g21999 ( 
.A1(n_21992),
.A2(n_8051),
.B(n_8043),
.Y(n_21999)
);

AOI21xp5_ASAP7_75t_L g22000 ( 
.A1(n_21992),
.A2(n_9067),
.B(n_9024),
.Y(n_22000)
);

AOI22xp5_ASAP7_75t_L g22001 ( 
.A1(n_21996),
.A2(n_11555),
.B1(n_11561),
.B2(n_11553),
.Y(n_22001)
);

OAI22xp5_ASAP7_75t_L g22002 ( 
.A1(n_21998),
.A2(n_9278),
.B1(n_9299),
.B2(n_9274),
.Y(n_22002)
);

OAI22xp33_ASAP7_75t_L g22003 ( 
.A1(n_21999),
.A2(n_9525),
.B1(n_9527),
.B2(n_9521),
.Y(n_22003)
);

AOI22xp5_ASAP7_75t_L g22004 ( 
.A1(n_21997),
.A2(n_11555),
.B1(n_11561),
.B2(n_11553),
.Y(n_22004)
);

OAI21xp5_ASAP7_75t_L g22005 ( 
.A1(n_22003),
.A2(n_22000),
.B(n_11150),
.Y(n_22005)
);

OR2x6_ASAP7_75t_L g22006 ( 
.A(n_22002),
.B(n_22004),
.Y(n_22006)
);

OR2x6_ASAP7_75t_L g22007 ( 
.A(n_22001),
.B(n_8675),
.Y(n_22007)
);

INVx1_ASAP7_75t_L g22008 ( 
.A(n_22006),
.Y(n_22008)
);

AND2x2_ASAP7_75t_L g22009 ( 
.A(n_22008),
.B(n_22007),
.Y(n_22009)
);

AOI221xp5_ASAP7_75t_L g22010 ( 
.A1(n_22009),
.A2(n_22005),
.B1(n_9527),
.B2(n_9532),
.C(n_9525),
.Y(n_22010)
);

AOI21xp5_ASAP7_75t_L g22011 ( 
.A1(n_22010),
.A2(n_8344),
.B(n_7718),
.Y(n_22011)
);

AOI211xp5_ASAP7_75t_L g22012 ( 
.A1(n_22011),
.A2(n_8710),
.B(n_8738),
.C(n_8701),
.Y(n_22012)
);


endmodule