module real_jpeg_2602_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_1),
.A2(n_37),
.B1(n_39),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_1),
.A2(n_56),
.B1(n_66),
.B2(n_68),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_3),
.A2(n_27),
.B1(n_37),
.B2(n_39),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_3),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_3),
.A2(n_27),
.B1(n_66),
.B2(n_68),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_4),
.A2(n_66),
.B1(n_68),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_4),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_79),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_6),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_6),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_6),
.A2(n_41),
.B1(n_66),
.B2(n_68),
.Y(n_179)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_8),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_8),
.A2(n_37),
.B1(n_39),
.B2(n_70),
.Y(n_126)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_11),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_11),
.A2(n_37),
.B1(n_39),
.B2(n_95),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_95),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_11),
.A2(n_66),
.B1(n_68),
.B2(n_95),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_12),
.B(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_12),
.B(n_42),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_12),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_12),
.A2(n_30),
.B(n_83),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_12),
.B(n_48),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g184 ( 
.A1(n_12),
.A2(n_39),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_12),
.B(n_63),
.C(n_66),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_12),
.B(n_77),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_12),
.B(n_106),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_13),
.A2(n_66),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_13),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_73),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_14),
.A2(n_66),
.B1(n_68),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_37),
.B1(n_39),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_16),
.A2(n_28),
.B1(n_30),
.B2(n_45),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_16),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_16),
.A2(n_45),
.B1(n_66),
.B2(n_68),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_130),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_129),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_108),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_22),
.B(n_108),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.C(n_97),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_23),
.B(n_97),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_57),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_43),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_25),
.B(n_43),
.C(n_57),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_40),
.B2(n_42),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_28),
.A2(n_35),
.A3(n_39),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_33),
.B(n_37),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_36),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_36),
.A2(n_93),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_36),
.A2(n_93),
.B1(n_94),
.B2(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_39),
.B1(n_52),
.B2(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_37),
.B(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_39),
.A2(n_50),
.A3(n_52),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_55),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_47),
.A2(n_90),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_47),
.A2(n_90),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_47),
.A2(n_89),
.B1(n_90),
.B2(n_137),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_47),
.A2(n_90),
.B1(n_136),
.B2(n_184),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

AO22x2_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_49),
.B(n_53),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_50),
.B(n_193),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_52),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_71),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_58),
.B(n_71),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_65),
.B2(n_69),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_59),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_60),
.A2(n_65),
.B1(n_146),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_61),
.A2(n_105),
.B1(n_106),
.B2(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_61),
.A2(n_106),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_61),
.A2(n_106),
.B1(n_147),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_61),
.A2(n_106),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_61),
.A2(n_106),
.B1(n_175),
.B2(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_66),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_66),
.B(n_203),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_76),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_74),
.A2(n_76),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_74),
.A2(n_76),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_77),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_77),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_75),
.A2(n_77),
.B1(n_86),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_75),
.A2(n_77),
.B1(n_155),
.B2(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_75),
.A2(n_77),
.B1(n_151),
.B2(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_75),
.A2(n_77),
.B1(n_205),
.B2(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_80),
.B(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_88),
.C(n_92),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_81),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_82),
.B(n_85),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_88),
.B(n_92),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_107),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_118),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_127),
.B2(n_128),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

AOI31xp33_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_225),
.A3(n_234),
.B(n_238),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_170),
.B(n_224),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_157),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_133),
.B(n_157),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_144),
.C(n_148),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_134),
.B(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_139),
.C(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_144),
.B(n_148),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_159),
.B(n_160),
.C(n_161),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_162),
.B(n_165),
.C(n_169),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_219),
.B(n_223),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_188),
.B(n_218),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_180),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_180),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_178),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_177),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_179),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_183),
.C(n_186),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_199),
.B(n_217),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_197),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_211),
.B(n_216),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_206),
.B(n_210),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_208),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_215),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_222),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_229),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.C(n_233),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);


endmodule