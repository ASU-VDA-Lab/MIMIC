module fake_jpeg_11557_n_582 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_582);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_582;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx8_ASAP7_75t_SL g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_60),
.Y(n_179)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_62),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_66),
.Y(n_149)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_20),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_69),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_20),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_70),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_11),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_76),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_73),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_11),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_77),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_80),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_21),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_82),
.A2(n_23),
.B1(n_52),
.B2(n_50),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_83),
.Y(n_195)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_12),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_86),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_36),
.B(n_12),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_87),
.Y(n_156)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_94),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_101),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_41),
.B(n_12),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_110),
.Y(n_139)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_22),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_106),
.B(n_23),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_38),
.B(n_12),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_121),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_49),
.B(n_17),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_111),
.B(n_118),
.C(n_50),
.Y(n_200)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_56),
.B(n_11),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_20),
.Y(n_119)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_122),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_38),
.B(n_8),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_49),
.A2(n_8),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_1),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_61),
.A2(n_26),
.B1(n_45),
.B2(n_31),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_129),
.A2(n_142),
.B(n_166),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_134),
.B(n_159),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_62),
.A2(n_26),
.B1(n_45),
.B2(n_31),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_103),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_147),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_98),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_155),
.B(n_158),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_83),
.B(n_42),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_83),
.B(n_48),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_87),
.B(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_162),
.B(n_171),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_62),
.A2(n_26),
.B1(n_24),
.B2(n_20),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_87),
.B(n_48),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_172),
.A2(n_198),
.B1(n_13),
.B2(n_14),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_60),
.A2(n_37),
.B1(n_54),
.B2(n_53),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_174),
.B(n_201),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_52),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_193),
.Y(n_235)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_69),
.Y(n_188)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_188),
.Y(n_271)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_70),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_120),
.B(n_68),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_120),
.B(n_113),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_197),
.B(n_199),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_96),
.A2(n_55),
.B1(n_54),
.B2(n_53),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_119),
.B(n_30),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_82),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_74),
.B(n_30),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_105),
.A2(n_55),
.B1(n_54),
.B2(n_53),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_55),
.B1(n_94),
.B2(n_93),
.Y(n_223)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_207),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_204),
.A2(n_79),
.B1(n_115),
.B2(n_101),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_210),
.A2(n_273),
.B1(n_130),
.B2(n_202),
.Y(n_289)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_211),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_213),
.Y(n_302)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_214),
.Y(n_296)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_215),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_136),
.Y(n_217)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_219),
.Y(n_321)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_220),
.Y(n_278)
);

AOI32xp33_ASAP7_75t_L g221 ( 
.A1(n_128),
.A2(n_141),
.A3(n_133),
.B1(n_147),
.B2(n_139),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_221),
.B(n_182),
.Y(n_303)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_223),
.A2(n_225),
.B1(n_231),
.B2(n_251),
.Y(n_285)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_129),
.A2(n_125),
.B1(n_123),
.B2(n_108),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_226),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_227),
.B(n_245),
.Y(n_308)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_142),
.A2(n_107),
.B1(n_102),
.B2(n_99),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_166),
.A2(n_91),
.B1(n_81),
.B2(n_80),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_233),
.A2(n_260),
.B1(n_274),
.B2(n_149),
.Y(n_298)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_153),
.Y(n_237)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_237),
.Y(n_293)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_239),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_240),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_194),
.A2(n_78),
.B1(n_77),
.B2(n_71),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_242),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_194),
.A2(n_63),
.B1(n_43),
.B2(n_6),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_243),
.A2(n_267),
.B1(n_152),
.B2(n_195),
.Y(n_312)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_246),
.B(n_252),
.Y(n_319)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

O2A1O1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_161),
.A2(n_43),
.B(n_5),
.C(n_7),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_249),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_177),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_148),
.A2(n_43),
.B1(n_1),
.B2(n_7),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_132),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_179),
.Y(n_253)
);

INVx4_ASAP7_75t_SL g304 ( 
.A(n_253),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_135),
.B(n_5),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_255),
.B(n_265),
.Y(n_326)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_257),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_177),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_156),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_259),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_178),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_205),
.A2(n_150),
.B1(n_185),
.B2(n_168),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_132),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_169),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_268),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_157),
.B(n_1),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_165),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_195),
.B(n_13),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g267 ( 
.A1(n_144),
.A2(n_43),
.B1(n_14),
.B2(n_15),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_140),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_163),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_269),
.B(n_275),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_151),
.B(n_13),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_270),
.B(n_180),
.Y(n_331)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_178),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_272),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_205),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_165),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_212),
.A2(n_227),
.B1(n_273),
.B2(n_251),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_277),
.A2(n_309),
.B1(n_312),
.B2(n_327),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_218),
.A2(n_140),
.B(n_149),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_288),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_289),
.A2(n_310),
.B1(n_220),
.B2(n_247),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_298),
.Y(n_364)
);

XNOR2x1_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_314),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_144),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_313),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_244),
.A2(n_151),
.B(n_182),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_329),
.C(n_240),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_227),
.A2(n_130),
.B1(n_185),
.B2(n_127),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_236),
.A2(n_138),
.B1(n_181),
.B2(n_127),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_235),
.B(n_181),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_236),
.A2(n_152),
.B(n_15),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_315),
.B(n_318),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_228),
.B(n_137),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_137),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_320),
.B(n_275),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_264),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_208),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_248),
.A2(n_138),
.B1(n_150),
.B2(n_168),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_254),
.B(n_170),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_328),
.B(n_331),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_267),
.A2(n_170),
.B1(n_180),
.B2(n_16),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_332),
.A2(n_333),
.B1(n_345),
.B2(n_346),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_267),
.B1(n_245),
.B2(n_246),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_285),
.A2(n_280),
.B1(n_298),
.B2(n_315),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_334),
.A2(n_338),
.B1(n_357),
.B2(n_358),
.Y(n_377)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_335),
.Y(n_385)
);

AO22x1_ASAP7_75t_L g337 ( 
.A1(n_306),
.A2(n_322),
.B1(n_267),
.B2(n_323),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_337),
.A2(n_341),
.B(n_283),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_285),
.A2(n_250),
.B1(n_209),
.B2(n_219),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_305),
.B(n_213),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_339),
.B(n_347),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_302),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_354),
.Y(n_383)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_291),
.Y(n_342)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_344),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_252),
.B1(n_261),
.B2(n_229),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_308),
.A2(n_217),
.B1(n_214),
.B2(n_206),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_319),
.Y(n_348)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_311),
.Y(n_350)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_350),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_271),
.C(n_224),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_355),
.C(n_371),
.Y(n_391)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_272),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_287),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_360),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_329),
.A2(n_207),
.B1(n_211),
.B2(n_259),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_324),
.A2(n_322),
.B1(n_309),
.B2(n_313),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_359),
.B(n_368),
.Y(n_406)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_325),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_363),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_326),
.B(n_263),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_258),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_318),
.A2(n_215),
.B1(n_234),
.B2(n_257),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_366),
.A2(n_374),
.B1(n_295),
.B2(n_304),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_286),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_370),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_293),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_279),
.B(n_253),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_369),
.Y(n_376)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_230),
.C(n_216),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_340),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_320),
.A2(n_293),
.B1(n_317),
.B2(n_301),
.Y(n_374)
);

OAI32xp33_ASAP7_75t_L g375 ( 
.A1(n_373),
.A2(n_301),
.A3(n_317),
.B1(n_292),
.B2(n_281),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_375),
.B(n_389),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_353),
.A2(n_284),
.B1(n_307),
.B2(n_282),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_388),
.B1(n_399),
.B2(n_332),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_353),
.A2(n_288),
.B(n_299),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_382),
.A2(n_393),
.B(n_395),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_373),
.A2(n_282),
.B(n_307),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_384),
.A2(n_370),
.B(n_350),
.Y(n_436)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_364),
.A2(n_290),
.B1(n_297),
.B2(n_300),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_374),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_283),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_404),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_334),
.A2(n_278),
.B1(n_290),
.B2(n_300),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_394),
.A2(n_402),
.B1(n_408),
.B2(n_366),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_337),
.A2(n_296),
.B(n_316),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_364),
.A2(n_278),
.B1(n_296),
.B2(n_321),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_396),
.A2(n_405),
.B1(n_357),
.B2(n_348),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_358),
.A2(n_297),
.B1(n_321),
.B2(n_316),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_349),
.A2(n_278),
.B1(n_276),
.B2(n_294),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_352),
.B(n_276),
.C(n_294),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_403),
.B(n_409),
.C(n_344),
.Y(n_427)
);

OA22x2_ASAP7_75t_L g404 ( 
.A1(n_333),
.A2(n_295),
.B1(n_284),
.B2(n_304),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_349),
.A2(n_304),
.B1(n_338),
.B2(n_341),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_336),
.Y(n_409)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_393),
.A2(n_337),
.B(n_351),
.C(n_354),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_413),
.B(n_414),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_386),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_371),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_427),
.C(n_391),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_408),
.A2(n_339),
.B1(n_367),
.B2(n_361),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_418),
.A2(n_431),
.B1(n_381),
.B2(n_405),
.Y(n_449)
);

BUFx24_ASAP7_75t_SL g419 ( 
.A(n_401),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_419),
.B(n_437),
.Y(n_466)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_379),
.Y(n_421)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_421),
.Y(n_443)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_378),
.Y(n_422)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_424),
.A2(n_438),
.B1(n_388),
.B2(n_404),
.Y(n_462)
);

FAx1_ASAP7_75t_SL g425 ( 
.A(n_409),
.B(n_355),
.CI(n_356),
.CON(n_425),
.SN(n_425)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_425),
.B(n_428),
.Y(n_460)
);

OAI21xp33_ASAP7_75t_L g426 ( 
.A1(n_376),
.A2(n_362),
.B(n_359),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_426),
.A2(n_403),
.B1(n_391),
.B2(n_406),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_363),
.B(n_335),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_387),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_429),
.B(n_441),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_396),
.B1(n_407),
.B2(n_398),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_377),
.A2(n_345),
.B1(n_346),
.B2(n_372),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_395),
.A2(n_360),
.B(n_342),
.Y(n_432)
);

XOR2x2_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_404),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_387),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_433),
.Y(n_447)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_385),
.Y(n_434)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_434),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_401),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_435),
.Y(n_453)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_R g437 ( 
.A1(n_375),
.A2(n_343),
.B1(n_382),
.B2(n_389),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_400),
.A2(n_407),
.B1(n_398),
.B2(n_397),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_376),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_439),
.B(n_442),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_383),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_440),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_383),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_406),
.B(n_390),
.Y(n_442)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_446),
.Y(n_476)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_449),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_418),
.A2(n_381),
.B1(n_377),
.B2(n_403),
.Y(n_450)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_458),
.C(n_464),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_412),
.A2(n_394),
.B1(n_380),
.B2(n_399),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_455),
.B(n_430),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_456),
.A2(n_425),
.B(n_440),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_415),
.B(n_391),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_457),
.B(n_461),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_415),
.B(n_385),
.C(n_392),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_427),
.B(n_402),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_462),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_463),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_411),
.B(n_392),
.C(n_379),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_410),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_432),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_435),
.A2(n_404),
.B1(n_410),
.B2(n_412),
.Y(n_469)
);

INVxp33_ASAP7_75t_L g475 ( 
.A(n_469),
.Y(n_475)
);

XOR2x2_ASAP7_75t_L g470 ( 
.A(n_411),
.B(n_404),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_463),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_437),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_473),
.B(n_488),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_485),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_471),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_484),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_457),
.B(n_420),
.C(n_441),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_480),
.B(n_483),
.C(n_486),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_420),
.C(n_433),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_444),
.B(n_439),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_467),
.A2(n_428),
.B(n_417),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_414),
.C(n_429),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_487),
.B(n_442),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_423),
.C(n_422),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_490),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_450),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_465),
.Y(n_491)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_491),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_492),
.A2(n_496),
.B1(n_447),
.B2(n_459),
.Y(n_512)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_465),
.Y(n_493)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_493),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_417),
.Y(n_494)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_494),
.Y(n_514)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_448),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_495),
.Y(n_517)
);

CKINVDCx14_ASAP7_75t_R g496 ( 
.A(n_445),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_468),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_501),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_464),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_470),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_510),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_479),
.B(n_466),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_503),
.B(n_509),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_413),
.Y(n_506)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_506),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_494),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_472),
.B(n_445),
.Y(n_510)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_472),
.B(n_449),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_515),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_491),
.Y(n_516)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_516),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_483),
.B(n_467),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_486),
.C(n_488),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_500),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_526),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_514),
.A2(n_475),
.B1(n_482),
.B2(n_497),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_524),
.A2(n_459),
.B1(n_447),
.B2(n_476),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_525),
.B(n_502),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_507),
.C(n_499),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_507),
.B(n_513),
.C(n_498),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_530),
.Y(n_548)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_516),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_508),
.Y(n_531)
);

CKINVDCx14_ASAP7_75t_R g538 ( 
.A(n_531),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_505),
.B(n_453),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_533),
.B(n_534),
.Y(n_536)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_511),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_498),
.B(n_490),
.C(n_505),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_535),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_477),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_546),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_529),
.B(n_510),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_539),
.B(n_547),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_519),
.A2(n_497),
.B1(n_477),
.B2(n_454),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_540),
.A2(n_545),
.B1(n_448),
.B2(n_451),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_542),
.B(n_532),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_543),
.A2(n_549),
.B1(n_481),
.B2(n_504),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_523),
.A2(n_454),
.B1(n_492),
.B2(n_476),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_521),
.B(n_520),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_504),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_525),
.A2(n_481),
.B1(n_485),
.B2(n_478),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_550),
.B(n_556),
.Y(n_562)
);

INVxp33_ASAP7_75t_SL g553 ( 
.A(n_536),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_553),
.B(n_554),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_528),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_520),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_555),
.B(n_557),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_544),
.A2(n_527),
.B(n_535),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_540),
.A2(n_538),
.B(n_542),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_547),
.B(n_532),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_558),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_559),
.B(n_560),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g565 ( 
.A1(n_552),
.A2(n_545),
.B(n_549),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_565),
.A2(n_566),
.B(n_568),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_553),
.A2(n_517),
.B(n_451),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_551),
.A2(n_517),
.B(n_495),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_563),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_571),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_561),
.A2(n_567),
.B1(n_564),
.B2(n_563),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_562),
.B(n_493),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_572),
.A2(n_573),
.B(n_487),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_567),
.A2(n_551),
.B(n_558),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_570),
.B(n_539),
.C(n_515),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_574),
.A2(n_575),
.B1(n_443),
.B2(n_434),
.Y(n_577)
);

MAJx2_ASAP7_75t_L g579 ( 
.A(n_577),
.B(n_578),
.C(n_436),
.Y(n_579)
);

NAND4xp25_ASAP7_75t_SL g578 ( 
.A(n_576),
.B(n_421),
.C(n_443),
.D(n_455),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_413),
.B1(n_424),
.B2(n_425),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_580),
.B(n_425),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_581),
.B(n_416),
.Y(n_582)
);


endmodule