module real_jpeg_28746_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_0),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_1),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_1),
.A2(n_26),
.B1(n_30),
.B2(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_173),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_1),
.A2(n_58),
.B1(n_60),
.B2(n_173),
.Y(n_257)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_3),
.A2(n_26),
.B1(n_30),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_36),
.B1(n_58),
.B2(n_60),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_3),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_4),
.A2(n_24),
.B1(n_52),
.B2(n_53),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_4),
.A2(n_24),
.B1(n_58),
.B2(n_60),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_6),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_6),
.A2(n_26),
.B1(n_30),
.B2(n_138),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_138),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_6),
.A2(n_58),
.B1(n_60),
.B2(n_138),
.Y(n_249)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_9),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_9),
.B(n_25),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_30),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_9),
.A2(n_30),
.B(n_209),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_171),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_9),
.A2(n_55),
.B(n_58),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_9),
.B(n_77),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_9),
.A2(n_116),
.B1(n_117),
.B2(n_257),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_26),
.B1(n_30),
.B2(n_45),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_10),
.A2(n_45),
.B1(n_58),
.B2(n_60),
.Y(n_186)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_12),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_12),
.A2(n_26),
.B1(n_30),
.B2(n_112),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_112),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_12),
.A2(n_58),
.B1(n_60),
.B2(n_112),
.Y(n_244)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_22),
.B1(n_23),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_14),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_14),
.A2(n_47),
.B1(n_58),
.B2(n_60),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_14),
.A2(n_26),
.B1(n_30),
.B2(n_47),
.Y(n_147)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_15),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_84),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_20),
.A2(n_43),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_21),
.A2(n_32),
.B(n_81),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_25),
.B(n_28),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_28),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g170 ( 
.A(n_22),
.B(n_171),
.CON(n_170),
.SN(n_170)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_25),
.A2(n_32),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_26),
.A2(n_30),
.B1(n_66),
.B2(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_26),
.A2(n_33),
.B1(n_170),
.B2(n_184),
.Y(n_183)
);

AOI32xp33_ASAP7_75t_L g207 ( 
.A1(n_26),
.A2(n_52),
.A3(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_207)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_28),
.B(n_30),
.Y(n_184)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_31),
.A2(n_44),
.B(n_48),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_32),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_38),
.B(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_74),
.C(n_79),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_39),
.A2(n_40),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.C(n_63),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_41),
.A2(n_42),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_43),
.A2(n_48),
.B1(n_111),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_43),
.A2(n_48),
.B1(n_137),
.B2(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_49),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_49),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_49),
.A2(n_63),
.B1(n_307),
.B2(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B(n_61),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_57),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_50),
.A2(n_104),
.B(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_50),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_50),
.A2(n_61),
.B(n_120),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_50),
.A2(n_57),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_50),
.A2(n_144),
.B(n_217),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_50),
.A2(n_57),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_50),
.A2(n_57),
.B1(n_216),
.B2(n_234),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_53),
.B(n_72),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_53),
.A2(n_56),
.B(n_171),
.C(n_236),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_103),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_57),
.B(n_171),
.Y(n_255)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_60),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_62),
.B(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_63),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_64),
.A2(n_76),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_65),
.B(n_69),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_65),
.A2(n_70),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_65),
.A2(n_70),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_65),
.A2(n_70),
.B1(n_167),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_65),
.A2(n_70),
.B1(n_195),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_68),
.A2(n_77),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_72),
.Y(n_208)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_76),
.A2(n_78),
.B(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_76),
.A2(n_134),
.B(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_79),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_332),
.B(n_338),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_302),
.A3(n_324),
.B1(n_330),
.B2(n_331),
.C(n_340),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_156),
.B(n_301),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_139),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_88),
.B(n_139),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_113),
.C(n_124),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_89),
.A2(n_90),
.B1(n_113),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_105),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_91),
.B(n_107),
.C(n_109),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_92),
.B(n_102),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_93),
.A2(n_117),
.B(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_94),
.A2(n_101),
.B(n_129),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_94),
.A2(n_99),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_95),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_117),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_98),
.A2(n_116),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_100),
.A2(n_116),
.B1(n_127),
.B2(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_113),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_123),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_114),
.A2(n_115),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_119),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_115),
.A2(n_150),
.B(n_153),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_116),
.A2(n_117),
.B1(n_249),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_119),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_121),
.B(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_124),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.C(n_135),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_125),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_130),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_291),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_133),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_154),
.B2(n_155),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_142),
.B(n_149),
.C(n_155),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_145),
.B(n_148),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_143),
.B(n_145),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_147),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_148),
.B(n_304),
.C(n_314),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_148),
.A2(n_304),
.B1(n_305),
.B2(n_329),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_148),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_295),
.B(n_300),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_199),
.B(n_281),
.C(n_294),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_187),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_159),
.B(n_187),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_174),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_161),
.B(n_162),
.C(n_174),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_169),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_171),
.B(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_172),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_182),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_176),
.B(n_180),
.C(n_182),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_188),
.A2(n_189),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_193),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_198),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_280),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_273),
.B(n_279),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_227),
.B(n_272),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_218),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_203),
.B(n_218),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_211),
.C(n_214),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_204),
.A2(n_205),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_219),
.B(n_225),
.C(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_266),
.B(n_271),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_245),
.B(n_265),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_230),
.B(n_237),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_253),
.B(n_264),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_251),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_258),
.B(n_263),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_256),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_275),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_292),
.B2(n_293),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_289),
.C(n_293),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_316),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_305)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_311),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_313),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_322),
.C(n_323),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_315),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_335),
.Y(n_337)
);


endmodule