module fake_jpeg_11635_n_473 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_473);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_473;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_48),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_92),
.Y(n_102)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx2_ASAP7_75t_SL g127 ( 
.A(n_54),
.Y(n_127)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_56),
.Y(n_150)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_60),
.B(n_81),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_87),
.Y(n_126)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_70),
.Y(n_140)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_78),
.Y(n_158)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_33),
.B(n_1),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_86),
.B(n_90),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_33),
.B(n_1),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_89),
.Y(n_136)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_55),
.B1(n_52),
.B2(n_50),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_17),
.B(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_96),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_100),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_41),
.B1(n_17),
.B2(n_26),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_103),
.A2(n_137),
.B1(n_139),
.B2(n_143),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_47),
.A2(n_30),
.B1(n_18),
.B2(n_26),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_109),
.A2(n_35),
.B1(n_3),
.B2(n_4),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_48),
.A2(n_41),
.B1(n_18),
.B2(n_28),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_109),
.B1(n_131),
.B2(n_24),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_123),
.A2(n_154),
.B1(n_23),
.B2(n_15),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_41),
.B1(n_28),
.B2(n_13),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_156),
.B1(n_14),
.B2(n_43),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_49),
.A2(n_14),
.B1(n_39),
.B2(n_25),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_51),
.A2(n_58),
.B1(n_56),
.B2(n_59),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_67),
.B(n_23),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_142),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_92),
.A2(n_28),
.B1(n_13),
.B2(n_30),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_43),
.C(n_39),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_142),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_54),
.A2(n_82),
.B(n_61),
.C(n_39),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_62),
.A2(n_77),
.B1(n_65),
.B2(n_68),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_96),
.B1(n_90),
.B2(n_86),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_64),
.A2(n_13),
.B1(n_43),
.B2(n_25),
.Y(n_156)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

AOI22x1_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_69),
.B1(n_72),
.B2(n_74),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_161),
.A2(n_169),
.B(n_157),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_61),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_176),
.Y(n_219)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_164),
.A2(n_197),
.B1(n_200),
.B2(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_100),
.B1(n_98),
.B2(n_73),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_180),
.B1(n_184),
.B2(n_192),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_102),
.Y(n_208)
);

AO22x1_ASAP7_75t_SL g174 ( 
.A1(n_104),
.A2(n_14),
.B1(n_15),
.B2(n_22),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_191),
.Y(n_207)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_107),
.B1(n_91),
.B2(n_89),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_107),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_190),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_196),
.Y(n_228)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_126),
.A2(n_24),
.B1(n_22),
.B2(n_15),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_139),
.A2(n_97),
.B1(n_23),
.B2(n_35),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_198),
.B1(n_140),
.B2(n_105),
.Y(n_223)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_120),
.A2(n_35),
.B1(n_3),
.B2(n_4),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_106),
.B(n_2),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_123),
.A2(n_35),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_35),
.B1(n_4),
.B2(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_136),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_147),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx5_ASAP7_75t_SL g235 ( 
.A(n_203),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g260 ( 
.A(n_208),
.B(n_229),
.C(n_219),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_185),
.B1(n_170),
.B2(n_199),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_204),
.B(n_146),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_220),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_237),
.B1(n_154),
.B2(n_140),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_179),
.A2(n_155),
.B1(n_110),
.B2(n_125),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_237),
.A2(n_192),
.B1(n_161),
.B2(n_182),
.Y(n_238)
);

AO21x2_ASAP7_75t_L g275 ( 
.A1(n_238),
.A2(n_258),
.B(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_170),
.B1(n_204),
.B2(n_164),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_240),
.A2(n_205),
.B1(n_220),
.B2(n_224),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_176),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_245),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_191),
.B(n_162),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_260),
.B(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_180),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_249),
.B(n_252),
.Y(n_283)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_206),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_253),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_235),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_185),
.B(n_161),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_234),
.B(n_223),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_165),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_259),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_260),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_185),
.B1(n_198),
.B2(n_174),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_207),
.B(n_208),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_261),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_184),
.B1(n_177),
.B2(n_186),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_263),
.B1(n_216),
.B2(n_232),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_215),
.A2(n_157),
.B1(n_187),
.B2(n_194),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_264),
.Y(n_290)
);

AOI32xp33_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_229),
.A3(n_213),
.B1(n_219),
.B2(n_234),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_265),
.A2(n_268),
.B(n_284),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_285),
.B1(n_287),
.B2(n_240),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_271),
.A2(n_273),
.B(n_291),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_255),
.A2(n_234),
.B(n_224),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_243),
.B1(n_261),
.B2(n_251),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_277),
.A2(n_281),
.B1(n_236),
.B2(n_218),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_256),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_248),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_249),
.A2(n_220),
.B1(n_209),
.B2(n_232),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_238),
.A2(n_125),
.B1(n_150),
.B2(n_101),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_225),
.C(n_235),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_242),
.C(n_258),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_252),
.A2(n_160),
.B1(n_171),
.B2(n_150),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_244),
.A2(n_135),
.B(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_286),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_294),
.Y(n_324)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_267),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_295),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_296),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_270),
.B(n_244),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_297),
.B(n_299),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_246),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_298),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_262),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_313),
.C(n_316),
.Y(n_326)
);

AO22x1_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_258),
.B1(n_174),
.B2(n_239),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_301),
.B(n_302),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_283),
.A2(n_258),
.B1(n_253),
.B2(n_257),
.Y(n_303)
);

XOR2x1_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_314),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g304 ( 
.A1(n_283),
.A2(n_258),
.B(n_263),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_305),
.B1(n_285),
.B2(n_282),
.Y(n_327)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_306),
.B(n_307),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_250),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_233),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_291),
.C(n_265),
.Y(n_319)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_315),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_273),
.B(n_277),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_311),
.A2(n_317),
.B1(n_318),
.B2(n_278),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_236),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_281),
.B(n_272),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_254),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_283),
.B(n_230),
.C(n_227),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_295),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_320),
.B(n_323),
.Y(n_355)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_321),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_271),
.B(n_275),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g369 ( 
.A1(n_322),
.A2(n_339),
.B(n_212),
.Y(n_369)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_287),
.B(n_275),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_327),
.A2(n_333),
.B1(n_345),
.B2(n_321),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_275),
.B(n_282),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_328),
.A2(n_314),
.B(n_311),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_303),
.A2(n_275),
.B1(n_278),
.B2(n_290),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_330),
.A2(n_254),
.B1(n_264),
.B2(n_211),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_304),
.A2(n_275),
.B1(n_290),
.B2(n_288),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_288),
.C(n_218),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_336),
.C(n_338),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_230),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_297),
.B(n_227),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_299),
.A2(n_289),
.B(n_279),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_293),
.B(n_168),
.C(n_210),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_318),
.C(n_306),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_302),
.B(n_298),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_344),
.B(n_201),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_304),
.A2(n_289),
.B1(n_279),
.B2(n_247),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_346),
.B(n_357),
.Y(n_387)
);

NOR3xp33_ASAP7_75t_SL g347 ( 
.A(n_324),
.B(n_294),
.C(n_325),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_370),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_SL g371 ( 
.A1(n_349),
.A2(n_328),
.B(n_331),
.C(n_333),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_307),
.Y(n_350)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_351),
.A2(n_331),
.B1(n_327),
.B2(n_345),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_332),
.A2(n_305),
.B1(n_316),
.B2(n_315),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_352),
.A2(n_359),
.B1(n_360),
.B2(n_362),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_332),
.A2(n_292),
.B1(n_317),
.B2(n_309),
.Y(n_353)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_301),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_368),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_217),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_363),
.C(n_364),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_330),
.A2(n_304),
.B1(n_301),
.B2(n_247),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_335),
.A2(n_322),
.B1(n_342),
.B2(n_339),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_210),
.C(n_226),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_334),
.B(n_337),
.C(n_336),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_342),
.A2(n_264),
.B1(n_217),
.B2(n_171),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_366),
.A2(n_101),
.B1(n_145),
.B2(n_212),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_329),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_226),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_349),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_325),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_359),
.C(n_369),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_341),
.C(n_337),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_381),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_352),
.Y(n_395)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_378),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_338),
.C(n_344),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_384),
.B(n_367),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_385),
.A2(n_152),
.B1(n_112),
.B2(n_114),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_196),
.C(n_195),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_386),
.B(n_390),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_370),
.A2(n_145),
.B1(n_114),
.B2(n_117),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_366),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_163),
.C(n_193),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_172),
.Y(n_391)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_391),
.Y(n_404)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_393),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_355),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_399),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_383),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_405),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_350),
.Y(n_398)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_398),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_358),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_374),
.B(n_362),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_402),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_356),
.C(n_368),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_382),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_360),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_406),
.Y(n_424)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_408),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_388),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_385),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_386),
.C(n_390),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_420),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_417),
.B(n_418),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_400),
.A2(n_371),
.B(n_383),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_409),
.A2(n_376),
.B(n_381),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_423),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_378),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_375),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_425),
.B(n_426),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_375),
.Y(n_426)
);

AO21x1_ASAP7_75t_L g427 ( 
.A1(n_398),
.A2(n_371),
.B(n_384),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_427),
.A2(n_410),
.B1(n_203),
.B2(n_105),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_397),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_434),
.C(n_424),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_419),
.B(n_392),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_430),
.B(n_436),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_403),
.C(n_406),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_432),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_371),
.C(n_396),
.Y(n_432)
);

AOI21x1_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_393),
.B(n_389),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_152),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_413),
.B(n_189),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_134),
.C(n_167),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_439),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_167),
.C(n_175),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_427),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_440),
.B(n_122),
.Y(n_452)
);

AOI21xp33_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_415),
.B(n_418),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_442),
.A2(n_449),
.B(n_141),
.Y(n_459)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_433),
.B(n_412),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_446),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_431),
.B(n_424),
.C(n_425),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_448),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_183),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_128),
.Y(n_449)
);

OAI21x1_ASAP7_75t_SL g457 ( 
.A1(n_452),
.A2(n_122),
.B(n_113),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_446),
.B(n_437),
.C(n_432),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_456),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_443),
.A2(n_438),
.B(n_439),
.Y(n_456)
);

O2A1O1Ixp33_ASAP7_75t_SL g463 ( 
.A1(n_457),
.A2(n_141),
.B(n_128),
.C(n_8),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_450),
.A2(n_451),
.B(n_437),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_458),
.Y(n_462)
);

NAND4xp25_ASAP7_75t_L g464 ( 
.A(n_459),
.B(n_6),
.C(n_7),
.D(n_9),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_454),
.A2(n_447),
.B(n_127),
.Y(n_461)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_461),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_463),
.B(n_464),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_462),
.A2(n_465),
.B(n_455),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_467),
.A2(n_11),
.B(n_9),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_466),
.A2(n_453),
.B1(n_460),
.B2(n_11),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_469),
.A2(n_470),
.B1(n_10),
.B2(n_11),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_471),
.A2(n_468),
.B(n_10),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_472),
.B(n_11),
.Y(n_473)
);


endmodule