module fake_jpeg_11690_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_7),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_48),
.B(n_64),
.Y(n_94)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_62),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_7),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_71),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_72),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_18),
.B(n_8),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_8),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_29),
.B1(n_37),
.B2(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_75),
.B1(n_103),
.B2(n_106),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_32),
.B1(n_25),
.B2(n_23),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_40),
.A2(n_17),
.B1(n_25),
.B2(n_23),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_78),
.A2(n_17),
.B1(n_20),
.B2(n_22),
.Y(n_148)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_87),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_38),
.A2(n_35),
.B1(n_18),
.B2(n_31),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_93),
.A2(n_106),
.B1(n_53),
.B2(n_44),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_60),
.B1(n_67),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_32),
.B1(n_25),
.B2(n_23),
.Y(n_106)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_112),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_66),
.B1(n_54),
.B2(n_70),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_113),
.A2(n_139),
.B1(n_144),
.B2(n_148),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_116),
.B(n_134),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_28),
.B(n_69),
.C(n_64),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_47),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_127),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_28),
.B1(n_18),
.B2(n_31),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_71),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_143),
.C(n_61),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_62),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_146),
.Y(n_166)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_31),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_133),
.Y(n_165)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_35),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_56),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_28),
.B1(n_35),
.B2(n_27),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_20),
.B1(n_22),
.B2(n_32),
.Y(n_168)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_27),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_149),
.Y(n_183)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_75),
.A2(n_45),
.B1(n_52),
.B2(n_59),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_86),
.B(n_82),
.C(n_58),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_76),
.A2(n_39),
.B1(n_50),
.B2(n_56),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_150),
.B(n_105),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_90),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_27),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_87),
.B(n_17),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_79),
.A2(n_57),
.B1(n_44),
.B2(n_53),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_151),
.A2(n_104),
.B1(n_83),
.B2(n_55),
.Y(n_154)
);

CKINVDCx6p67_ASAP7_75t_R g207 ( 
.A(n_152),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_124),
.A2(n_55),
.B1(n_83),
.B2(n_79),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_160),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_104),
.B1(n_82),
.B2(n_86),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_89),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_179),
.C(n_181),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_112),
.B(n_20),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_170),
.B(n_150),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_133),
.B1(n_116),
.B2(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_117),
.B1(n_146),
.B2(n_119),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_22),
.B(n_95),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_56),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_175),
.B(n_184),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_141),
.B1(n_139),
.B2(n_148),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_142),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_90),
.C(n_32),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_0),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_131),
.B(n_8),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_161),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_188),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_183),
.B(n_137),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_190),
.B(n_206),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_191),
.A2(n_210),
.B1(n_176),
.B2(n_171),
.Y(n_244)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_169),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_117),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_197),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_123),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_198),
.B(n_200),
.Y(n_250)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_123),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_118),
.B(n_130),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_170),
.B(n_152),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_143),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_202),
.B(n_209),
.C(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_129),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_143),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_160),
.A2(n_141),
.B1(n_132),
.B2(n_136),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_180),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_211),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_121),
.B1(n_147),
.B2(n_140),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_174),
.B(n_169),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_156),
.B1(n_165),
.B2(n_182),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_218),
.B1(n_219),
.B2(n_189),
.Y(n_247)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_145),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_221),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_186),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_172),
.A2(n_141),
.B1(n_138),
.B2(n_0),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_159),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_187),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_0),
.C(n_1),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_185),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_223),
.Y(n_251)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_224),
.B(n_1),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_232),
.B(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_166),
.B1(n_177),
.B2(n_153),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_235),
.B1(n_244),
.B2(n_245),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_194),
.A2(n_181),
.B(n_177),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_177),
.B1(n_181),
.B2(n_167),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_207),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_207),
.A2(n_177),
.B(n_174),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_239),
.A2(n_243),
.B(n_246),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_252),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_187),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_185),
.B1(n_171),
.B2(n_176),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_201),
.A2(n_8),
.B(n_2),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_247),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_211),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_9),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_206),
.A2(n_190),
.B1(n_218),
.B2(n_205),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_189),
.B1(n_204),
.B2(n_219),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_1),
.C(n_3),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_257),
.C(n_222),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_209),
.B(n_15),
.C(n_4),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_259),
.B(n_240),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_193),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_269),
.C(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_247),
.A2(n_207),
.B1(n_188),
.B2(n_197),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_291)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_225),
.Y(n_266)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_274),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_271),
.B1(n_237),
.B2(n_251),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_199),
.C(n_192),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_217),
.B1(n_208),
.B2(n_214),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_204),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_276),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_223),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_278),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_224),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_238),
.A2(n_212),
.B1(n_215),
.B2(n_220),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_238),
.A2(n_220),
.B1(n_4),
.B2(n_5),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_3),
.C(n_5),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_229),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_236),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_230),
.B(n_3),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_255),
.C(n_227),
.Y(n_298)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_288),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_234),
.B(n_5),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_278),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_312),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_235),
.B1(n_231),
.B2(n_253),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_295),
.A2(n_268),
.B1(n_265),
.B2(n_271),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_263),
.A2(n_232),
.B1(n_249),
.B2(n_243),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_296),
.A2(n_311),
.B1(n_245),
.B2(n_251),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_304),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_250),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_300),
.C(n_302),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_252),
.C(n_250),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_272),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_261),
.A2(n_243),
.B(n_258),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_305),
.A2(n_265),
.B(n_287),
.Y(n_327)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_240),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_313),
.C(n_290),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_263),
.A2(n_232),
.B1(n_228),
.B2(n_239),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_288),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_257),
.Y(n_313)
);

XNOR2x1_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_264),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_315),
.B(n_320),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_261),
.B(n_287),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_326),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_319),
.A2(n_312),
.B1(n_314),
.B2(n_291),
.Y(n_343)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_321),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_277),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_323),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_302),
.C(n_300),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_324),
.B(n_335),
.C(n_298),
.Y(n_341)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_297),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_337),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_328),
.A2(n_336),
.B1(n_309),
.B2(n_306),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_295),
.A2(n_233),
.B(n_246),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_331),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_267),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_330),
.A2(n_334),
.B1(n_314),
.B2(n_309),
.Y(n_348)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_299),
.B(n_282),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_333),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_285),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_259),
.C(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

NOR3xp33_ASAP7_75t_SL g340 ( 
.A(n_322),
.B(n_307),
.C(n_301),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_342),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_320),
.C(n_315),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_324),
.B(n_296),
.C(n_289),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_334),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_286),
.C(n_303),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_352),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_306),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_319),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_303),
.C(n_292),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_325),
.B(n_292),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_355),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_322),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_338),
.A2(n_318),
.B(n_327),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_356),
.A2(n_365),
.B(n_337),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_358),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_338),
.A2(n_344),
.B(n_339),
.Y(n_360)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_332),
.C(n_316),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_363),
.B(n_368),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_342),
.A2(n_316),
.B(n_330),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_366),
.B(n_347),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g367 ( 
.A(n_351),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_367),
.B(n_341),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_343),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_329),
.C(n_328),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_370),
.B(n_347),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_372),
.B(n_376),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_359),
.C(n_356),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_382),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_362),
.A2(n_364),
.B1(n_354),
.B2(n_346),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_377),
.A2(n_380),
.B1(n_270),
.B2(n_266),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_366),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_379),
.A2(n_283),
.B(n_262),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_360),
.A2(n_321),
.B1(n_340),
.B2(n_273),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_369),
.B(n_323),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_381),
.B(n_248),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_370),
.A2(n_363),
.B1(n_357),
.B2(n_358),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_387),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_375),
.B(n_349),
.C(n_333),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_384),
.B(n_257),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_242),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_391),
.C(n_392),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_349),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_6),
.Y(n_394)
);

AOI21x1_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_377),
.B(n_371),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_242),
.Y(n_391)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_393),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_394),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_396),
.C(n_397),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_390),
.A2(n_385),
.B(n_384),
.Y(n_398)
);

O2A1O1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_398),
.A2(n_400),
.B(n_12),
.C(n_13),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_387),
.A2(n_6),
.B(n_10),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_12),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_383),
.A2(n_6),
.B(n_10),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_402),
.A2(n_404),
.B(n_405),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_403),
.B(n_13),
.C(n_14),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_407),
.Y(n_408)
);

OAI321xp33_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_406),
.A3(n_401),
.B1(n_402),
.B2(n_15),
.C(n_14),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_14),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_15),
.Y(n_411)
);


endmodule