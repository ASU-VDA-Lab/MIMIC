module fake_jpeg_31241_n_530 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_530);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_12),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_53),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_54),
.Y(n_149)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_60),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_61),
.B(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_13),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_65),
.B(n_66),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_12),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_69),
.B(n_101),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_70),
.Y(n_128)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_36),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_87),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_80),
.Y(n_117)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_0),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_93),
.Y(n_125)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_32),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_97),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_100),
.Y(n_131)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_44),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_0),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_31),
.B(n_1),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_18),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_105),
.B(n_31),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_30),
.B1(n_48),
.B2(n_45),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_116),
.A2(n_92),
.B1(n_96),
.B2(n_102),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_119),
.B(n_127),
.Y(n_190)
);

BUFx2_ASAP7_75t_R g120 ( 
.A(n_66),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_120),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_35),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_124),
.B(n_154),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_63),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_53),
.B(n_37),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_156),
.Y(n_178)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_58),
.B(n_35),
.Y(n_154)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_90),
.Y(n_155)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_50),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_162),
.Y(n_180)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_81),
.B(n_37),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_33),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_93),
.B(n_50),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_74),
.B(n_52),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_74),
.B(n_52),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_113),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_168),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_25),
.B1(n_40),
.B2(n_46),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_169),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_170),
.B(n_177),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_171),
.Y(n_259)
);

OA22x2_ASAP7_75t_L g224 ( 
.A1(n_173),
.A2(n_182),
.B1(n_108),
.B2(n_141),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_108),
.A2(n_56),
.B1(n_67),
.B2(n_73),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_175),
.B1(n_202),
.B2(n_210),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_138),
.A2(n_75),
.B1(n_86),
.B2(n_77),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_132),
.A2(n_25),
.B1(n_29),
.B2(n_46),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_176),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_111),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_25),
.B1(n_29),
.B2(n_46),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_179),
.A2(n_128),
.B1(n_117),
.B2(n_54),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_130),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_181),
.B(n_209),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g182 ( 
.A1(n_105),
.A2(n_76),
.B1(n_91),
.B2(n_89),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_129),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_185),
.B(n_188),
.Y(n_244)
);

CKINVDCx12_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_80),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_191),
.B(n_194),
.Y(n_260)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_80),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_135),
.Y(n_195)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_137),
.B(n_33),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_203),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_140),
.B(n_60),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_217),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_142),
.A2(n_30),
.B1(n_48),
.B2(n_45),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_27),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_144),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_27),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_208),
.Y(n_223)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_28),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_55),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_146),
.A2(n_30),
.B1(n_48),
.B2(n_49),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_125),
.B(n_43),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_43),
.Y(n_236)
);

CKINVDCx9p33_ASAP7_75t_R g213 ( 
.A(n_107),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_216),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_115),
.B(n_31),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_218),
.B(n_24),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_153),
.B(n_114),
.Y(n_219)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_224),
.B(n_245),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_236),
.B(n_183),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_211),
.A2(n_128),
.B1(n_109),
.B2(n_114),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_201),
.A2(n_109),
.B1(n_159),
.B2(n_112),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_240),
.A2(n_213),
.B1(n_117),
.B2(n_214),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_170),
.A2(n_134),
.B(n_121),
.Y(n_243)
);

NAND2x1_ASAP7_75t_SL g292 ( 
.A(n_243),
.B(n_172),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_217),
.A2(n_106),
.B(n_118),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_230),
.B(n_235),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_141),
.B1(n_126),
.B2(n_145),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_173),
.B1(n_143),
.B2(n_99),
.Y(n_273)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_167),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_257),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_106),
.C(n_72),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_218),
.Y(n_290)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_208),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_206),
.Y(n_263)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_187),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_279),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_264),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_190),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_212),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_269),
.A2(n_292),
.B(n_246),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_178),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_270),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_223),
.B(n_220),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_271),
.B(n_273),
.Y(n_312)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_231),
.B(n_180),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_276),
.B(n_289),
.Y(n_317)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_235),
.A2(n_215),
.B1(n_172),
.B2(n_216),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_278),
.A2(n_239),
.B1(n_259),
.B2(n_242),
.Y(n_302)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_280),
.Y(n_303)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_227),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_282),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_224),
.A2(n_182),
.B(n_189),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_283),
.Y(n_332)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_182),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_288),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_221),
.B(n_186),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_244),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_230),
.B(n_218),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g293 ( 
.A1(n_252),
.A2(n_143),
.B1(n_196),
.B2(n_148),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_293),
.A2(n_297),
.B1(n_233),
.B2(n_254),
.Y(n_318)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_298),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_224),
.A2(n_222),
.B1(n_252),
.B2(n_223),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_221),
.B(n_197),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_299),
.B(n_247),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_302),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_286),
.A2(n_222),
.B1(n_224),
.B2(n_249),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_307),
.A2(n_318),
.B1(n_321),
.B2(n_327),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_291),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_269),
.A2(n_256),
.B(n_243),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_309),
.A2(n_319),
.B(n_305),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_287),
.A2(n_236),
.B(n_245),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_283),
.A2(n_145),
.B1(n_150),
.B2(n_148),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_322),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_234),
.C(n_225),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_334),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_283),
.A2(n_150),
.B1(n_133),
.B2(n_126),
.Y(n_327)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_229),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_282),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_283),
.A2(n_233),
.B1(n_168),
.B2(n_166),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_331),
.A2(n_297),
.B1(n_273),
.B2(n_275),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_251),
.C(n_207),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_336),
.B(n_340),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_317),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_337),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_308),
.A2(n_292),
.B(n_267),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_339),
.A2(n_349),
.B(n_314),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_332),
.A2(n_287),
.B1(n_298),
.B2(n_270),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_341),
.A2(n_351),
.B1(n_352),
.B2(n_363),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_292),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_360),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_343),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_271),
.Y(n_345)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_345),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_301),
.B(n_291),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_359),
.C(n_309),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_317),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_347),
.Y(n_373)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_313),
.Y(n_348)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_263),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_355),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_312),
.A2(n_270),
.B1(n_279),
.B2(n_289),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_272),
.B1(n_277),
.B2(n_284),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_310),
.B(n_272),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_353),
.B(n_357),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_331),
.A2(n_264),
.B1(n_296),
.B2(n_295),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_321),
.Y(n_386)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_255),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_301),
.B(n_299),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_315),
.B(n_255),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_300),
.B(n_237),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_362),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_322),
.B(n_239),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_333),
.A2(n_242),
.B1(n_264),
.B2(n_171),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

OAI32xp33_ASAP7_75t_L g365 ( 
.A1(n_305),
.A2(n_281),
.A3(n_274),
.B1(n_294),
.B2(n_237),
.Y(n_365)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_300),
.B(n_239),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_187),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_304),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_367),
.A2(n_318),
.B1(n_307),
.B2(n_327),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_344),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_364),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_378),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_337),
.B(n_304),
.Y(n_378)
);

XOR2x2_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_319),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_320),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_381),
.A2(n_386),
.B1(n_251),
.B2(n_204),
.Y(n_424)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_384),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_387),
.A2(n_349),
.B(n_339),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_330),
.Y(n_388)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_388),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_348),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_280),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_391),
.B(n_349),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_314),
.Y(n_392)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_338),
.B(n_326),
.Y(n_393)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_341),
.A2(n_320),
.B1(n_328),
.B2(n_316),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_394),
.A2(n_355),
.B1(n_313),
.B2(n_316),
.Y(n_414)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_395),
.Y(n_423)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_396),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_344),
.B(n_329),
.C(n_328),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_350),
.C(n_325),
.Y(n_415)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_356),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_398),
.Y(n_405)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_401),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_389),
.A2(n_306),
.B1(n_354),
.B2(n_358),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_403),
.A2(n_404),
.B1(n_409),
.B2(n_413),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_389),
.A2(n_396),
.B1(n_377),
.B2(n_387),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_406),
.B(n_410),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_408),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_388),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_399),
.A2(n_358),
.B1(n_335),
.B2(n_340),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_399),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_416),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_395),
.A2(n_335),
.B1(n_359),
.B2(n_342),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_414),
.A2(n_424),
.B1(n_375),
.B2(n_382),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_420),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_380),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_372),
.B(n_325),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_373),
.A2(n_306),
.B1(n_311),
.B2(n_303),
.Y(n_421)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_421),
.Y(n_439)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_425),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_199),
.C(n_192),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_426),
.B(n_375),
.C(n_394),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_370),
.B(n_372),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_392),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_428),
.B(n_431),
.C(n_437),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_429),
.B(n_441),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_400),
.A2(n_391),
.B(n_379),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_430),
.A2(n_198),
.B(n_2),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_374),
.C(n_379),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_433),
.A2(n_443),
.B1(n_450),
.B2(n_192),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_416),
.B(n_369),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_435),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_369),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_436),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_374),
.C(n_398),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_400),
.A2(n_414),
.B1(n_417),
.B2(n_418),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_376),
.Y(n_444)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_444),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_402),
.B(n_376),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_445),
.B(n_280),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_404),
.Y(n_446)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_413),
.A2(n_371),
.B(n_385),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_447),
.A2(n_41),
.B(n_20),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_409),
.A2(n_386),
.B1(n_381),
.B2(n_371),
.Y(n_450)
);

OAI321xp33_ASAP7_75t_L g451 ( 
.A1(n_438),
.A2(n_405),
.A3(n_422),
.B1(n_410),
.B2(n_419),
.C(n_385),
.Y(n_451)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_405),
.Y(n_452)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_450),
.A2(n_426),
.B1(n_420),
.B2(n_427),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_455),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_458),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_41),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_464),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_434),
.A2(n_439),
.B1(n_449),
.B2(n_433),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_463),
.A2(n_428),
.B1(n_429),
.B2(n_440),
.Y(n_481)
);

BUFx12_ASAP7_75t_L g464 ( 
.A(n_436),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_465),
.A2(n_430),
.B(n_2),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_1),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_1),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_446),
.A2(n_122),
.B1(n_118),
.B2(n_59),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_467),
.A2(n_469),
.B1(n_40),
.B2(n_24),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_443),
.A2(n_122),
.B1(n_193),
.B2(n_24),
.Y(n_469)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_470),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_437),
.C(n_431),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_474),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_462),
.B(n_434),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_477),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_452),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_459),
.B(n_461),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_482),
.C(n_24),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_458),
.B(n_441),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_481),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_466),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_432),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_484),
.A2(n_31),
.B(n_3),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_440),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_485),
.Y(n_494)
);

A2O1A1Ixp33_ASAP7_75t_SL g488 ( 
.A1(n_486),
.A2(n_465),
.B(n_469),
.C(n_467),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_476),
.A2(n_464),
.B(n_468),
.Y(n_487)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_487),
.Y(n_507)
);

AO21x1_ASAP7_75t_L g504 ( 
.A1(n_488),
.A2(n_489),
.B(n_493),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_SL g489 ( 
.A1(n_473),
.A2(n_456),
.B(n_463),
.C(n_454),
.Y(n_489)
);

MAJx2_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_454),
.C(n_460),
.Y(n_490)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_490),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_496),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_40),
.C(n_3),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_473),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_499),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_2),
.C(n_3),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_484),
.C(n_485),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_501),
.B(n_483),
.Y(n_503)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_503),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_475),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_505),
.B(n_506),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_478),
.C(n_486),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_478),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_512),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_494),
.A2(n_470),
.B(n_474),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_5),
.C(n_6),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_4),
.C(n_5),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_507),
.A2(n_491),
.B1(n_488),
.B2(n_493),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_514),
.B(n_518),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_511),
.A2(n_4),
.B(n_5),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_516),
.A2(n_508),
.B(n_504),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_7),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_519),
.B(n_515),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_513),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_521),
.B(n_522),
.C(n_523),
.Y(n_524)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g525 ( 
.A1(n_520),
.A2(n_504),
.B(n_517),
.C(n_512),
.D(n_519),
.Y(n_525)
);

AOI31xp33_ASAP7_75t_L g526 ( 
.A1(n_525),
.A2(n_524),
.A3(n_502),
.B(n_10),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_7),
.B(n_9),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_9),
.C(n_10),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_528),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_529),
.B(n_11),
.Y(n_530)
);


endmodule