module fake_aes_1999_n_691 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_691);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_691;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_597;
wire n_349;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_59), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_42), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_30), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_8), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_34), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_36), .Y(n_84) );
INVx3_ASAP7_75t_L g85 ( .A(n_2), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_50), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_31), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_57), .Y(n_88) );
INVx1_ASAP7_75t_SL g89 ( .A(n_63), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_4), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_72), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_20), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_38), .Y(n_93) );
INVxp67_ASAP7_75t_SL g94 ( .A(n_56), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_17), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_19), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_60), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_5), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_78), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_58), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_10), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_29), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_27), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_62), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_15), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_76), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_26), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_37), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_47), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_39), .Y(n_110) );
BUFx2_ASAP7_75t_SL g111 ( .A(n_10), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_51), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_64), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_6), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_21), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_48), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_1), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_16), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_12), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_41), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_3), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_6), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_49), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_11), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_67), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_46), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_117), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_117), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_111), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_99), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
INVx4_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_80), .B(n_33), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_85), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_99), .Y(n_136) );
NAND2xp33_ASAP7_75t_SL g137 ( .A(n_113), .B(n_0), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_125), .B(n_0), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_80), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_105), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_105), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_125), .B(n_1), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_119), .B(n_2), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_90), .Y(n_146) );
XOR2xp5_ASAP7_75t_L g147 ( .A(n_121), .B(n_3), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_88), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_79), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_86), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_90), .Y(n_152) );
INVxp67_ASAP7_75t_L g153 ( .A(n_111), .Y(n_153) );
BUFx8_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_96), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_124), .B(n_4), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_91), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_124), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_97), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_102), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_82), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_104), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_98), .B(n_5), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_106), .B(n_43), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_101), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_114), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_107), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_108), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_157), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_140), .B(n_112), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_157), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_158), .A2(n_122), .B(n_84), .C(n_83), .Y(n_172) );
AOI22x1_ASAP7_75t_L g173 ( .A1(n_140), .A2(n_116), .B1(n_123), .B2(n_120), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_133), .B(n_92), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_141), .B(n_115), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_133), .B(n_91), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_145), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_133), .B(n_92), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_135), .B(n_84), .Y(n_181) );
BUFx6f_ASAP7_75t_SL g182 ( .A(n_138), .Y(n_182) );
BUFx5_ASAP7_75t_L g183 ( .A(n_134), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_141), .B(n_88), .Y(n_185) );
NAND3xp33_ASAP7_75t_L g186 ( .A(n_130), .B(n_88), .C(n_118), .Y(n_186) );
NOR3xp33_ASAP7_75t_L g187 ( .A(n_137), .B(n_100), .C(n_94), .Y(n_187) );
O2A1O1Ixp5_ASAP7_75t_L g188 ( .A1(n_160), .A2(n_95), .B(n_89), .C(n_88), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_160), .B(n_88), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_145), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_128), .B(n_126), .Y(n_192) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_138), .B(n_126), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_149), .Y(n_195) );
INVxp67_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_153), .B(n_110), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_128), .B(n_110), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_149), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_168), .B(n_109), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_138), .B(n_109), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_149), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_168), .B(n_103), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_127), .B(n_103), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_138), .A2(n_81), .B1(n_8), .B2(n_9), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_146), .B(n_81), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_165), .B(n_44), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_129), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_139), .B(n_45), .Y(n_209) );
NAND2x1p5_ASAP7_75t_L g210 ( .A(n_156), .B(n_7), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_129), .B(n_7), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_132), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_139), .B(n_52), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_161), .B(n_9), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_156), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_165), .B(n_11), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_150), .B(n_12), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_150), .B(n_13), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_151), .B(n_13), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_144), .A2(n_14), .B1(n_15), .B2(n_18), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_165), .B(n_14), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_151), .B(n_22), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_166), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_155), .B(n_23), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_166), .B(n_24), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_178), .A2(n_167), .B(n_155), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_217), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_223), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_169), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_225), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_208), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_208), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_179), .B(n_163), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_212), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_183), .B(n_219), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_213), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_201), .A2(n_154), .B1(n_163), .B2(n_134), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_174), .B(n_154), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_176), .B(n_154), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_171), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_210), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_171), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_180), .B(n_166), .Y(n_245) );
BUFx2_ASAP7_75t_L g246 ( .A(n_169), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_181), .B(n_167), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_219), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_183), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_209), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_183), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_196), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_209), .Y(n_254) );
AND2x6_ASAP7_75t_L g255 ( .A(n_201), .B(n_134), .Y(n_255) );
INVx4_ASAP7_75t_L g256 ( .A(n_182), .Y(n_256) );
INVx4_ASAP7_75t_L g257 ( .A(n_182), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_183), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_184), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_183), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_214), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_216), .B(n_162), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_201), .B(n_162), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_189), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_203), .B(n_159), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_191), .B(n_159), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_183), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_182), .B(n_143), .Y(n_269) );
OR2x6_ASAP7_75t_L g270 ( .A(n_200), .B(n_143), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_183), .B(n_136), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_177), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_170), .B(n_134), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_224), .B(n_136), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_187), .B(n_143), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_211), .Y(n_276) );
BUFx2_ASAP7_75t_L g277 ( .A(n_192), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_218), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_170), .B(n_134), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_175), .B(n_134), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_204), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_177), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_188), .A2(n_164), .B(n_134), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_193), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_220), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_175), .B(n_164), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_215), .B(n_164), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_172), .B(n_164), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_193), .B(n_148), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_221), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_198), .B(n_164), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_234), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_239), .A2(n_205), .B1(n_197), .B2(n_200), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_234), .Y(n_294) );
OAI33xp33_ASAP7_75t_L g295 ( .A1(n_263), .A2(n_142), .A3(n_148), .B1(n_206), .B2(n_131), .B3(n_226), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_248), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_233), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_242), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_236), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_253), .B(n_147), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_287), .A2(n_185), .B(n_190), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_289), .B(n_186), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_266), .B(n_173), .Y(n_303) );
NOR2xp67_ASAP7_75t_SL g304 ( .A(n_256), .B(n_164), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_238), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_242), .B(n_147), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_264), .B(n_142), .Y(n_308) );
OR2x6_ASAP7_75t_L g309 ( .A(n_264), .B(n_131), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_267), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_256), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_246), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_243), .B(n_222), .Y(n_313) );
AOI22xp33_ASAP7_75t_SL g314 ( .A1(n_284), .A2(n_227), .B1(n_207), .B2(n_214), .Y(n_314) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_256), .B(n_25), .Y(n_315) );
BUFx4_ASAP7_75t_SL g316 ( .A(n_244), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_266), .B(n_190), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_244), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_229), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_248), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_230), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_252), .B(n_185), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_286), .A2(n_202), .B(n_199), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_248), .B(n_202), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_247), .B(n_28), .Y(n_325) );
CKINVDCx8_ASAP7_75t_R g326 ( .A(n_277), .Y(n_326) );
BUFx2_ASAP7_75t_SL g327 ( .A(n_257), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_273), .A2(n_199), .B(n_195), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_235), .B(n_32), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_257), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_281), .B(n_35), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_279), .A2(n_195), .B(n_194), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_257), .B(n_40), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_260), .B(n_53), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_259), .Y(n_335) );
INVx4_ASAP7_75t_L g336 ( .A(n_255), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_255), .A2(n_289), .B1(n_275), .B2(n_265), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_280), .A2(n_194), .B(n_55), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_270), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_275), .B(n_54), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_231), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_275), .B(n_77), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_299), .Y(n_343) );
AOI211x1_ASAP7_75t_L g344 ( .A1(n_293), .A2(n_228), .B(n_288), .C(n_291), .Y(n_344) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_338), .A2(n_283), .B(n_274), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_312), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_305), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_325), .A2(n_323), .B(n_332), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_328), .A2(n_274), .B(n_261), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_308), .B(n_284), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_336), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_292), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_292), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_335), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_308), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_296), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_326), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_297), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_336), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_340), .A2(n_268), .B(n_251), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_302), .A2(n_265), .B(n_237), .Y(n_362) );
HB1xp67_ASAP7_75t_SL g363 ( .A(n_298), .Y(n_363) );
AOI21xp33_ASAP7_75t_SL g364 ( .A1(n_315), .A2(n_231), .B(n_240), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_297), .Y(n_365) );
AO31x2_ASAP7_75t_L g366 ( .A1(n_303), .A2(n_269), .A3(n_245), .B(n_290), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_296), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_306), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_310), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_296), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_320), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_313), .A2(n_255), .B1(n_270), .B2(n_276), .Y(n_372) );
NAND3xp33_ASAP7_75t_L g373 ( .A(n_314), .B(n_270), .C(n_269), .Y(n_373) );
OA21x2_ASAP7_75t_L g374 ( .A1(n_301), .A2(n_271), .B(n_285), .Y(n_374) );
NOR2x1_ASAP7_75t_SL g375 ( .A(n_350), .B(n_308), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_356), .B(n_309), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_359), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_369), .B(n_315), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_369), .B(n_294), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_359), .B(n_294), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_356), .B(n_365), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_365), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_351), .B(n_333), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_351), .B(n_333), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_352), .B(n_313), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_351), .B(n_311), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_357), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_354), .B(n_337), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_354), .B(n_337), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_354), .B(n_321), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_343), .B(n_319), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_353), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_353), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_343), .B(n_309), .Y(n_400) );
NAND2x1_ASAP7_75t_L g401 ( .A(n_367), .B(n_320), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_347), .Y(n_402) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_377), .A2(n_372), .B1(n_373), .B2(n_241), .C(n_364), .Y(n_403) );
OAI211xp5_ASAP7_75t_SL g404 ( .A1(n_395), .A2(n_307), .B(n_358), .C(n_368), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_379), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_378), .Y(n_406) );
AOI31xp33_ASAP7_75t_L g407 ( .A1(n_380), .A2(n_364), .A3(n_316), .B(n_300), .Y(n_407) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_380), .A2(n_270), .B1(n_368), .B2(n_347), .C(n_355), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_383), .A2(n_350), .B1(n_373), .B2(n_309), .Y(n_409) );
OA21x2_ASAP7_75t_L g410 ( .A1(n_396), .A2(n_348), .B(n_361), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_378), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_383), .B(n_355), .Y(n_412) );
AO21x2_ASAP7_75t_L g413 ( .A1(n_396), .A2(n_398), .B(n_399), .Y(n_413) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_378), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_389), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_379), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_397), .B(n_339), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_389), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_400), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_397), .B(n_302), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_381), .B(n_366), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_400), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_396), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_398), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_366), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_398), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_392), .B(n_357), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_382), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_387), .B(n_331), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_387), .A2(n_393), .B1(n_392), .B2(n_318), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_399), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_394), .B(n_366), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_399), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_384), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_394), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_433), .B(n_402), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_411), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_433), .B(n_402), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_421), .B(n_393), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_405), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g443 ( .A1(n_404), .A2(n_318), .B(n_329), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_436), .B(n_376), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_421), .B(n_391), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_426), .B(n_375), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_405), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_426), .B(n_428), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_429), .B(n_376), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_415), .B(n_366), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_420), .B(n_375), .Y(n_451) );
OAI32xp33_ASAP7_75t_L g452 ( .A1(n_412), .A2(n_391), .A3(n_342), .B1(n_316), .B2(n_367), .Y(n_452) );
AND2x4_ASAP7_75t_SL g453 ( .A(n_425), .B(n_385), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_431), .A2(n_255), .B1(n_385), .B2(n_386), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_416), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_412), .B(n_344), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_415), .B(n_391), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_416), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_435), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_415), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_435), .B(n_344), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_418), .B(n_366), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_414), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_407), .B(n_350), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_403), .B(n_295), .C(n_334), .Y(n_465) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_418), .B(n_385), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_411), .Y(n_467) );
NOR2x1p5_ASAP7_75t_L g468 ( .A(n_417), .B(n_386), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_419), .B(n_366), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_437), .B(n_386), .Y(n_470) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_411), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_425), .B(n_391), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_437), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_422), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_408), .A2(n_295), .B1(n_322), .B2(n_317), .C(n_278), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_406), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_428), .B(n_385), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_431), .B(n_386), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_428), .B(n_388), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_406), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_423), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_430), .B(n_350), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_423), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_424), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_427), .B(n_388), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_438), .B(n_428), .Y(n_487) );
INVx5_ASAP7_75t_L g488 ( .A(n_463), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_439), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_441), .B(n_427), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_447), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_441), .B(n_434), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_443), .B(n_409), .C(n_278), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_445), .B(n_434), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_445), .B(n_434), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_438), .B(n_432), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_463), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_464), .B(n_327), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_440), .B(n_432), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_440), .B(n_432), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_474), .B(n_424), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_442), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_460), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_448), .B(n_424), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_444), .B(n_413), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_448), .B(n_413), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_448), .B(n_413), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_479), .B(n_410), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_479), .B(n_410), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_439), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_453), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_446), .B(n_410), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_449), .B(n_410), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_455), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_450), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_451), .B(n_350), .Y(n_517) );
OR2x6_ASAP7_75t_L g518 ( .A(n_446), .B(n_401), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_446), .B(n_388), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_467), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_458), .B(n_390), .Y(n_521) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_466), .B(n_401), .Y(n_522) );
INVxp67_ASAP7_75t_L g523 ( .A(n_462), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_467), .Y(n_524) );
AOI222xp33_ASAP7_75t_L g525 ( .A1(n_468), .A2(n_255), .B1(n_362), .B2(n_390), .C1(n_341), .C2(n_322), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_450), .B(n_388), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_453), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_481), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_457), .B(n_390), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_473), .B(n_390), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_457), .B(n_388), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_470), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_476), .Y(n_534) );
NOR2xp67_ASAP7_75t_SL g535 ( .A(n_469), .B(n_311), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_456), .B(n_388), .Y(n_536) );
NOR2x1_ASAP7_75t_L g537 ( .A(n_462), .B(n_357), .Y(n_537) );
NAND5xp2_ASAP7_75t_SL g538 ( .A(n_454), .B(n_362), .C(n_65), .D(n_66), .E(n_68), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_482), .B(n_330), .Y(n_539) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_471), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_478), .B(n_330), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_481), .B(n_374), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_465), .B(n_278), .C(n_314), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_483), .B(n_374), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_503), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_492), .B(n_485), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_515), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_526), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_540), .A2(n_452), .B(n_461), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_490), .B(n_469), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_492), .B(n_485), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_491), .Y(n_552) );
AOI31xp33_ASAP7_75t_L g553 ( .A1(n_528), .A2(n_478), .A3(n_477), .B(n_475), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_498), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_512), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_543), .A2(n_452), .B1(n_472), .B2(n_477), .C(n_484), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_509), .B(n_483), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_509), .B(n_472), .Y(n_558) );
OR2x6_ASAP7_75t_L g559 ( .A(n_518), .B(n_480), .Y(n_559) );
NOR2xp67_ASAP7_75t_SL g560 ( .A(n_488), .B(n_370), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_533), .B(n_480), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_505), .B(n_486), .Y(n_562) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_490), .B(n_486), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_501), .B(n_374), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_510), .B(n_348), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_505), .B(n_370), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_501), .B(n_374), .Y(n_567) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_497), .A2(n_370), .B(n_367), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_534), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_488), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_500), .B(n_367), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_510), .B(n_348), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_502), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_500), .B(n_371), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_507), .B(n_361), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_516), .B(n_523), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_493), .A2(n_345), .B1(n_262), .B2(n_254), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_496), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_506), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_507), .B(n_508), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_508), .B(n_361), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_487), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_494), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_494), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_488), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_535), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_513), .B(n_345), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_489), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_495), .B(n_345), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_495), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_521), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_489), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_488), .B(n_353), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_514), .B(n_345), .Y(n_596) );
NAND2xp33_ASAP7_75t_L g597 ( .A(n_512), .B(n_371), .Y(n_597) );
NAND4xp75_ASAP7_75t_L g598 ( .A(n_556), .B(n_563), .C(n_570), .D(n_587), .Y(n_598) );
NAND2xp33_ASAP7_75t_SL g599 ( .A(n_570), .B(n_513), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_584), .B(n_488), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_555), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_597), .A2(n_538), .B(n_537), .Y(n_603) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_581), .A2(n_536), .B(n_541), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_580), .B(n_531), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g606 ( .A(n_549), .B(n_525), .C(n_499), .D(n_517), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_553), .B(n_539), .C(n_519), .Y(n_607) );
NOR4xp25_ASAP7_75t_L g608 ( .A(n_547), .B(n_527), .C(n_544), .D(n_542), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_548), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g610 ( .A(n_588), .B(n_519), .C(n_542), .Y(n_610) );
NOR4xp25_ASAP7_75t_L g611 ( .A(n_574), .B(n_527), .C(n_544), .D(n_520), .Y(n_611) );
NAND4xp25_ASAP7_75t_L g612 ( .A(n_578), .B(n_532), .C(n_529), .D(n_524), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_576), .B(n_518), .C(n_511), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_569), .B(n_518), .C(n_511), .Y(n_614) );
OAI321xp33_ASAP7_75t_L g615 ( .A1(n_559), .A2(n_518), .A3(n_522), .B1(n_530), .B2(n_532), .C(n_529), .Y(n_615) );
AOI222xp33_ASAP7_75t_L g616 ( .A1(n_593), .A2(n_524), .B1(n_520), .B2(n_262), .C1(n_250), .C2(n_254), .Y(n_616) );
NAND4xp25_ASAP7_75t_SL g617 ( .A(n_550), .B(n_530), .C(n_522), .D(n_70), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_573), .B(n_353), .C(n_371), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_554), .Y(n_620) );
OA211x2_ASAP7_75t_L g621 ( .A1(n_568), .A2(n_61), .B(n_69), .C(n_71), .Y(n_621) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_597), .B(n_360), .Y(n_622) );
NOR2x1_ASAP7_75t_L g623 ( .A(n_559), .B(n_360), .Y(n_623) );
NOR2x1p5_ASAP7_75t_L g624 ( .A(n_585), .B(n_360), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_586), .B(n_349), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_582), .B(n_371), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_561), .B(n_351), .C(n_360), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_587), .A2(n_324), .B(n_271), .C(n_237), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_592), .A2(n_262), .B1(n_254), .B2(n_250), .C(n_304), .Y(n_629) );
NAND3xp33_ASAP7_75t_SL g630 ( .A(n_579), .B(n_73), .C(n_74), .Y(n_630) );
NOR2xp67_ASAP7_75t_L g631 ( .A(n_582), .B(n_75), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_563), .A2(n_371), .B1(n_320), .B2(n_349), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_579), .B(n_371), .C(n_262), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_595), .B(n_324), .C(n_349), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_607), .A2(n_565), .B1(n_572), .B2(n_557), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_600), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_608), .B(n_557), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_612), .A2(n_559), .B1(n_571), .B2(n_595), .Y(n_638) );
OAI22xp33_ASAP7_75t_SL g639 ( .A1(n_602), .A2(n_575), .B1(n_567), .B2(n_564), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_598), .B(n_596), .C(n_565), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_609), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_619), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_606), .B(n_558), .Y(n_643) );
NAND4xp25_ASAP7_75t_SL g644 ( .A(n_610), .B(n_558), .C(n_546), .D(n_551), .Y(n_644) );
NAND4xp75_ASAP7_75t_L g645 ( .A(n_631), .B(n_572), .C(n_583), .D(n_577), .Y(n_645) );
INVxp33_ASAP7_75t_SL g646 ( .A(n_611), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_620), .Y(n_647) );
INVx3_ASAP7_75t_L g648 ( .A(n_599), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_604), .A2(n_577), .B1(n_583), .B2(n_546), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_605), .B(n_562), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_601), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_625), .B(n_551), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_613), .A2(n_589), .B(n_566), .Y(n_653) );
AOI21xp33_ASAP7_75t_L g654 ( .A1(n_616), .A2(n_615), .B(n_614), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_627), .B(n_560), .C(n_594), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_624), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_626), .B(n_589), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g658 ( .A1(n_654), .A2(n_603), .B(n_632), .C(n_623), .Y(n_658) );
NOR2x1p5_ASAP7_75t_L g659 ( .A(n_648), .B(n_630), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_643), .B(n_590), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_640), .B(n_629), .C(n_618), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_648), .B(n_622), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_651), .B(n_590), .Y(n_663) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_647), .Y(n_664) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_644), .B(n_617), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_646), .B(n_594), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_637), .A2(n_603), .B(n_633), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_636), .Y(n_668) );
AND4x1_ASAP7_75t_L g669 ( .A(n_635), .B(n_629), .C(n_621), .D(n_634), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g670 ( .A(n_653), .B(n_628), .C(n_591), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_639), .A2(n_254), .B1(n_250), .B2(n_320), .C(n_282), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_665), .A2(n_653), .B1(n_649), .B2(n_645), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_664), .B(n_641), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_666), .A2(n_638), .B1(n_656), .B2(n_650), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_658), .A2(n_655), .B1(n_642), .B2(n_657), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_662), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_668), .Y(n_677) );
AND2x4_ASAP7_75t_L g678 ( .A(n_659), .B(n_652), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g679 ( .A(n_669), .B(n_282), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_677), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_672), .A2(n_667), .B1(n_670), .B2(n_660), .C(n_661), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_673), .Y(n_682) );
NAND5xp2_ASAP7_75t_L g683 ( .A(n_675), .B(n_671), .C(n_661), .D(n_663), .E(n_250), .Y(n_683) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_676), .B(n_258), .C(n_272), .D(n_251), .Y(n_684) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_680), .A2(n_679), .B(n_674), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_681), .B(n_678), .Y(n_686) );
OAI321xp33_ASAP7_75t_L g687 ( .A1(n_682), .A2(n_678), .A3(n_248), .B1(n_272), .B2(n_261), .C(n_268), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_686), .A2(n_683), .B1(n_684), .B2(n_258), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_687), .B(n_249), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_689), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_690), .A2(n_685), .B(n_688), .Y(n_691) );
endmodule