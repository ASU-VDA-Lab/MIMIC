module fake_jpeg_2191_n_98 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_20),
.B1(n_16),
.B2(n_21),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_24),
.A2(n_15),
.B1(n_11),
.B2(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_43),
.B1(n_15),
.B2(n_34),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_14),
.B(n_19),
.C(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_47),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_21),
.B1(n_23),
.B2(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_53),
.B1(n_56),
.B2(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_25),
.B1(n_13),
.B2(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_4),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_28),
.B1(n_27),
.B2(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

OA21x2_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_43),
.B(n_45),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_63),
.B1(n_48),
.B2(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_43),
.B1(n_36),
.B2(n_44),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_50),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_52),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.C(n_62),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_57),
.C(n_59),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_58),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_63),
.B1(n_48),
.B2(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_67),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_72),
.C(n_77),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_88),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_61),
.C(n_65),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_85),
.A2(n_83),
.B(n_81),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_90),
.B(n_65),
.Y(n_92)
);

NOR2xp67_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_83),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_92),
.A2(n_93),
.B(n_7),
.C(n_9),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_5),
.C(n_6),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.C(n_7),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_92),
.A2(n_76),
.B(n_9),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_10),
.B(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_76),
.Y(n_98)
);


endmodule