module fake_jpeg_30834_n_531 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_531);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_4),
.B(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_8),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_55),
.B(n_70),
.Y(n_120)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_62),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_67),
.B(n_96),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_14),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_39),
.B(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_82),
.Y(n_129)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_38),
.B(n_15),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_88),
.B(n_95),
.Y(n_148)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_92),
.Y(n_161)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_33),
.B(n_13),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_34),
.B(n_12),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_51),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_34),
.B(n_13),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_102),
.B(n_17),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_16),
.B1(n_40),
.B2(n_53),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_109),
.A2(n_125),
.B1(n_133),
.B2(n_162),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_116),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_70),
.B(n_51),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_58),
.A2(n_16),
.B1(n_40),
.B2(n_35),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_16),
.B1(n_40),
.B2(n_35),
.Y(n_133)
);

BUFx6f_ASAP7_75t_SL g134 ( 
.A(n_97),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_61),
.A2(n_23),
.B1(n_35),
.B2(n_42),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_74),
.B(n_17),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_82),
.B(n_25),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_63),
.A2(n_23),
.B1(n_35),
.B2(n_42),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_101),
.B1(n_83),
.B2(n_85),
.Y(n_184)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_138),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_177),
.B(n_204),
.Y(n_245)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_179),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_184),
.A2(n_151),
.B1(n_152),
.B2(n_146),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_163),
.A2(n_103),
.B1(n_99),
.B2(n_56),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_185),
.A2(n_198),
.B1(n_219),
.B2(n_224),
.Y(n_241)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_194),
.Y(n_230)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_190),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_195),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_76),
.C(n_64),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_120),
.B(n_25),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_199),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_65),
.B1(n_88),
.B2(n_71),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_62),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_120),
.B(n_20),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_200),
.B(n_202),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

BUFx16f_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_169),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

NOR2x1_ASAP7_75t_R g204 ( 
.A(n_129),
.B(n_42),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_150),
.A2(n_129),
.B(n_131),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_128),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

AO22x2_ASAP7_75t_L g207 ( 
.A1(n_133),
.A2(n_78),
.B1(n_68),
.B2(n_23),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_207),
.A2(n_213),
.B1(n_109),
.B2(n_171),
.Y(n_247)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_123),
.A2(n_27),
.B1(n_52),
.B2(n_31),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_209),
.A2(n_50),
.B1(n_43),
.B2(n_22),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

BUFx2_ASAP7_75t_SL g244 ( 
.A(n_210),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_146),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_216),
.Y(n_233)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_137),
.A2(n_20),
.B1(n_48),
.B2(n_18),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_223),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_148),
.B(n_121),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_161),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_124),
.B(n_19),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_225),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_141),
.A2(n_52),
.B1(n_27),
.B2(n_31),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_113),
.A2(n_88),
.B1(n_52),
.B2(n_31),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_125),
.A2(n_27),
.B(n_19),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_227),
.B(n_230),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_228),
.A2(n_247),
.B1(n_48),
.B2(n_18),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_174),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_235),
.B(n_251),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_237),
.A2(n_240),
.B1(n_257),
.B2(n_198),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_176),
.A2(n_166),
.B1(n_135),
.B2(n_154),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_174),
.B(n_204),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_207),
.A2(n_119),
.B1(n_166),
.B2(n_156),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_252),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_207),
.A2(n_119),
.B1(n_165),
.B2(n_153),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_254),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_207),
.A2(n_153),
.B1(n_167),
.B2(n_161),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_285),
.Y(n_315)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_269),
.Y(n_316)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_270),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_272),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_188),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_183),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_273),
.B(n_287),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_258),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_274),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_183),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_276),
.Y(n_319)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_196),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_295),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_223),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_236),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_281),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_282),
.A2(n_285),
.B1(n_265),
.B2(n_284),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_288),
.B1(n_246),
.B2(n_220),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_227),
.B(n_181),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_178),
.C(n_175),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_231),
.C(n_226),
.Y(n_326)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_241),
.A2(n_162),
.B1(n_224),
.B2(n_185),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_239),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_294),
.B1(n_259),
.B2(n_229),
.Y(n_303)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_292),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_255),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_238),
.B(n_189),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_293),
.A2(n_297),
.B(n_235),
.Y(n_300)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g295 ( 
.A(n_251),
.B(n_217),
.CI(n_117),
.CON(n_295),
.SN(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_245),
.B(n_182),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_296),
.B(n_255),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_230),
.B(n_249),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_249),
.B(n_263),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_298),
.A2(n_299),
.B(n_308),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_263),
.B(n_245),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_322),
.Y(n_351)
);

OAI22x1_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_263),
.B1(n_247),
.B2(n_244),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_302),
.A2(n_303),
.B(n_304),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_279),
.A2(n_288),
.B(n_296),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_278),
.A2(n_253),
.B1(n_246),
.B2(n_215),
.Y(n_308)
);

NOR2x1p5_ASAP7_75t_SL g310 ( 
.A(n_277),
.B(n_127),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_173),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_276),
.B1(n_267),
.B2(n_130),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_313),
.A2(n_302),
.B1(n_308),
.B2(n_282),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_320),
.B(n_232),
.Y(n_342)
);

AO21x2_ASAP7_75t_L g321 ( 
.A1(n_283),
.A2(n_255),
.B(n_258),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_321),
.A2(n_294),
.B1(n_274),
.B2(n_289),
.Y(n_348)
);

AOI32xp33_ASAP7_75t_L g322 ( 
.A1(n_295),
.A2(n_248),
.A3(n_226),
.B1(n_203),
.B2(n_208),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_327),
.C(n_320),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_231),
.C(n_248),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_296),
.A2(n_177),
.B(n_195),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_328),
.A2(n_299),
.B(n_298),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_329),
.A2(n_331),
.B1(n_348),
.B2(n_350),
.Y(n_367)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_306),
.Y(n_330)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_313),
.A2(n_284),
.B1(n_295),
.B2(n_275),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_332),
.B(n_336),
.C(n_353),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_290),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_232),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_304),
.A2(n_266),
.B(n_281),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_335),
.A2(n_341),
.B(n_344),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_324),
.C(n_326),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_312),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_310),
.B(n_315),
.Y(n_339)
);

XOR2x1_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_316),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_312),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_340),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_317),
.A2(n_287),
.B(n_292),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_342),
.B(n_320),
.Y(n_373)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_343),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_345),
.A2(n_323),
.B1(n_314),
.B2(n_303),
.Y(n_360)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_309),
.Y(n_346)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_301),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_302),
.A2(n_271),
.B1(n_216),
.B2(n_179),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_319),
.A2(n_270),
.B(n_269),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_355),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_232),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_319),
.A2(n_210),
.B(n_191),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_357),
.Y(n_370)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_321),
.A2(n_260),
.B1(n_187),
.B2(n_193),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_314),
.B1(n_318),
.B2(n_323),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_359),
.B(n_373),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_360),
.A2(n_365),
.B1(n_382),
.B2(n_355),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_351),
.A2(n_321),
.B1(n_315),
.B2(n_322),
.Y(n_365)
);

OAI22x1_ASAP7_75t_SL g366 ( 
.A1(n_354),
.A2(n_321),
.B1(n_311),
.B2(n_300),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_366),
.A2(n_335),
.B1(n_333),
.B2(n_344),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_371),
.A2(n_372),
.B1(n_378),
.B2(n_387),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_329),
.A2(n_321),
.B1(n_301),
.B2(n_307),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_307),
.Y(n_375)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_358),
.A2(n_321),
.B1(n_328),
.B2(n_325),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_347),
.B(n_325),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_380),
.B(n_388),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_384),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_343),
.A2(n_316),
.B1(n_260),
.B2(n_206),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_342),
.C(n_349),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_201),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_250),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_389),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_350),
.A2(n_218),
.B1(n_264),
.B2(n_154),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_352),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_334),
.B(n_250),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_390),
.A2(n_362),
.B1(n_360),
.B2(n_367),
.Y(n_429)
);

AO21x1_ASAP7_75t_L g393 ( 
.A1(n_386),
.A2(n_354),
.B(n_333),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_400),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_346),
.Y(n_394)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_394),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_395),
.B(n_259),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_340),
.Y(n_396)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_396),
.Y(n_425)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_376),
.Y(n_397)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_386),
.A2(n_341),
.B(n_331),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_399),
.A2(n_413),
.B1(n_415),
.B2(n_372),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_338),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_369),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_403),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_339),
.C(n_353),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_410),
.C(n_359),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_370),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_330),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_404),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_374),
.B(n_356),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_405),
.A2(n_408),
.B(n_411),
.Y(n_430)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_345),
.C(n_357),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_264),
.Y(n_411)
);

FAx1_ASAP7_75t_SL g412 ( 
.A(n_373),
.B(n_365),
.CI(n_383),
.CON(n_412),
.SN(n_412)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_414),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_259),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_201),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_379),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_22),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_420),
.A2(n_417),
.B1(n_411),
.B2(n_392),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_389),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_421),
.B(n_424),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_381),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_412),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_367),
.C(n_371),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_432),
.C(n_436),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_429),
.A2(n_415),
.B1(n_413),
.B2(n_423),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_409),
.B(n_387),
.C(n_256),
.Y(n_432)
);

NOR3xp33_ASAP7_75t_SL g433 ( 
.A(n_407),
.B(n_13),
.C(n_12),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_433),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_259),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_438),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_396),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_256),
.C(n_139),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_147),
.C(n_50),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_418),
.C(n_397),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_393),
.B(n_43),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_435),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_SL g442 ( 
.A(n_391),
.B(n_192),
.Y(n_442)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_442),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_443),
.B(n_444),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_416),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_394),
.Y(n_447)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

FAx1_ASAP7_75t_SL g448 ( 
.A(n_439),
.B(n_391),
.CI(n_403),
.CON(n_448),
.SN(n_448)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_448),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_453),
.Y(n_468)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_460),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_433),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_456),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_398),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_399),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_419),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_426),
.B(n_412),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_395),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_459),
.A2(n_454),
.B1(n_441),
.B2(n_451),
.Y(n_474)
);

XNOR2x1_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_404),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_461),
.A2(n_431),
.B1(n_422),
.B2(n_417),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_434),
.C(n_421),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_472),
.C(n_476),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_446),
.A2(n_423),
.B(n_425),
.Y(n_464)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_467),
.A2(n_192),
.B1(n_2),
.B2(n_3),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_460),
.A2(n_411),
.B1(n_438),
.B2(n_419),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_470),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_450),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_440),
.C(n_436),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_474),
.A2(n_448),
.B1(n_451),
.B2(n_450),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_400),
.C(n_408),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_461),
.A2(n_437),
.B(n_46),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_477),
.A2(n_453),
.B(n_11),
.Y(n_483)
);

FAx1_ASAP7_75t_SL g478 ( 
.A(n_449),
.B(n_11),
.CI(n_12),
.CON(n_478),
.SN(n_478)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_478),
.B(n_9),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_458),
.B(n_46),
.C(n_45),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_45),
.C(n_29),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_473),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_480),
.B(n_483),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_445),
.Y(n_481)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_481),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_485),
.C(n_492),
.Y(n_507)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_486),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_462),
.B(n_46),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_493),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_468),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_491),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_463),
.B(n_45),
.C(n_29),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_29),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_495),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_468),
.B(n_26),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_490),
.A2(n_475),
.B(n_472),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_500),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_466),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_499),
.A2(n_502),
.B(n_491),
.Y(n_513)
);

XOR2x1_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_470),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_488),
.A2(n_469),
.B(n_479),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_501),
.A2(n_17),
.B(n_2),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_SL g502 ( 
.A1(n_483),
.A2(n_478),
.B1(n_466),
.B2(n_471),
.Y(n_502)
);

OAI321xp33_ASAP7_75t_L g503 ( 
.A1(n_493),
.A2(n_26),
.A3(n_17),
.B1(n_3),
.B2(n_4),
.C(n_0),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_503),
.B(n_494),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_498),
.B(n_492),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_510),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_507),
.B(n_482),
.C(n_485),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_511),
.A2(n_497),
.B1(n_504),
.B2(n_505),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_484),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_0),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_513),
.A2(n_515),
.B(n_504),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_514),
.B(n_0),
.C(n_3),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_506),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_519),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_518),
.A2(n_521),
.B(n_515),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_523),
.A2(n_5),
.B(n_6),
.Y(n_526)
);

NOR2xp67_ASAP7_75t_SL g524 ( 
.A(n_520),
.B(n_516),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_0),
.B(n_3),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_525),
.B(n_526),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_527),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_522),
.C(n_6),
.Y(n_529)
);

MAJx2_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_7),
.C(n_5),
.Y(n_530)
);

AOI221xp5_ASAP7_75t_SL g531 ( 
.A1(n_530),
.A2(n_6),
.B1(n_7),
.B2(n_528),
.C(n_433),
.Y(n_531)
);


endmodule