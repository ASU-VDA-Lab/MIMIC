module fake_jpeg_614_n_439 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_439);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_439;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_61),
.Y(n_98)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_15),
.B(n_14),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_44),
.C(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_32),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_68),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_65),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_77),
.Y(n_132)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_19),
.B(n_13),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_44),
.Y(n_103)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_20),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_21),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_85),
.Y(n_128)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_21),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_25),
.B(n_40),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_90),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_41),
.B1(n_35),
.B2(n_27),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_93),
.A2(n_122),
.B1(n_30),
.B2(n_28),
.Y(n_142)
);

OR2x2_ASAP7_75t_SL g168 ( 
.A(n_102),
.B(n_82),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_103),
.B(n_119),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_54),
.B(n_27),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_75),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_64),
.A2(n_20),
.B1(n_24),
.B2(n_27),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_110),
.A2(n_112),
.B1(n_87),
.B2(n_86),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_20),
.B1(n_40),
.B2(n_23),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_116),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_55),
.A2(n_45),
.B1(n_79),
.B2(n_71),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_23),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_49),
.A2(n_35),
.B1(n_42),
.B2(n_36),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_65),
.A2(n_43),
.B1(n_42),
.B2(n_36),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_131),
.A2(n_75),
.B1(n_65),
.B2(n_26),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_62),
.B(n_34),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_62),
.B(n_34),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_58),
.B(n_26),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_52),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_137),
.B(n_161),
.Y(n_217)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_143),
.Y(n_198)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_72),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_141),
.B(n_150),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_142),
.A2(n_162),
.B1(n_135),
.B2(n_50),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_169),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g149 ( 
.A(n_101),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_149),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_30),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_155),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_158),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_120),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_166),
.Y(n_200)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_160),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_28),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_98),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_179),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_29),
.C(n_35),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_73),
.B(n_16),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_170),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_104),
.A2(n_67),
.B1(n_57),
.B2(n_60),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_171),
.A2(n_172),
.B1(n_3),
.B2(n_6),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_104),
.A2(n_91),
.B1(n_88),
.B2(n_89),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_174),
.Y(n_190)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_177),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_125),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_91),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_97),
.B(n_115),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_181),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_SL g182 ( 
.A(n_112),
.B(n_16),
.C(n_29),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_99),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_178),
.B1(n_142),
.B2(n_141),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_186),
.A2(n_199),
.B1(n_214),
.B2(n_157),
.Y(n_244)
);

AO22x1_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_135),
.B1(n_117),
.B2(n_124),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_205),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_131),
.CI(n_110),
.CON(n_189),
.SN(n_189)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_189),
.B(n_152),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_195),
.A2(n_196),
.B1(n_203),
.B2(n_207),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_105),
.B1(n_124),
.B2(n_117),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_150),
.A2(n_51),
.B1(n_59),
.B2(n_47),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_105),
.B(n_1),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_202),
.A2(n_206),
.B(n_7),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_125),
.B1(n_84),
.B2(n_111),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_123),
.B(n_111),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_147),
.A2(n_123),
.B1(n_92),
.B2(n_99),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_218),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_140),
.A2(n_99),
.B1(n_29),
.B2(n_2),
.Y(n_214)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_153),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_163),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_6),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_164),
.A2(n_29),
.B1(n_5),
.B2(n_6),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_176),
.B1(n_173),
.B2(n_159),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_223),
.A2(n_203),
.B1(n_191),
.B2(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_155),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_225),
.B(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_168),
.C(n_167),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_236),
.C(n_257),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_228),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_184),
.A2(n_170),
.B1(n_154),
.B2(n_158),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_244),
.B1(n_258),
.B2(n_199),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_179),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_233),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_215),
.Y(n_231)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_138),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_146),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_240),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_151),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_149),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_237),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_187),
.B(n_200),
.Y(n_261)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_160),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_144),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_242),
.B(n_249),
.Y(n_288)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_192),
.B(n_174),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_187),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_157),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_254),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_188),
.B(n_6),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_252),
.B(n_7),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_253),
.A2(n_202),
.B(n_206),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_210),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_210),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_215),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_256),
.B(n_191),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_188),
.C(n_204),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_259),
.A2(n_264),
.B(n_292),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_261),
.B(n_250),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_193),
.B(n_200),
.Y(n_264)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_195),
.B1(n_196),
.B2(n_193),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_266),
.A2(n_280),
.B1(n_284),
.B2(n_231),
.Y(n_314)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_277),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_198),
.C(n_200),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_290),
.C(n_243),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_198),
.Y(n_277)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_243),
.A2(n_212),
.B1(n_189),
.B2(n_207),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_218),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_283),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_282),
.A2(n_241),
.B1(n_224),
.B2(n_226),
.Y(n_303)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_189),
.B(n_218),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_233),
.A2(n_222),
.B1(n_221),
.B2(n_185),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_183),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_287),
.B(n_291),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_253),
.A2(n_219),
.B(n_214),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_250),
.B(n_247),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_227),
.B(n_218),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_240),
.A2(n_183),
.B(n_9),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_295),
.A2(n_309),
.B(n_318),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_278),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_298),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_271),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_237),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_301),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_245),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_260),
.B(n_236),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_277),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_319),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_307),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_254),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_312),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_243),
.C(n_248),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_321),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_274),
.A2(n_247),
.B1(n_229),
.B2(n_234),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_271),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_255),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_314),
.A2(n_320),
.B1(n_265),
.B2(n_275),
.Y(n_342)
);

INVx3_ASAP7_75t_SL g315 ( 
.A(n_270),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_315),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_262),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_264),
.A2(n_228),
.B(n_231),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_263),
.B(n_251),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_258),
.B1(n_256),
.B2(n_239),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_185),
.C(n_290),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_305),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_322),
.B(n_345),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_283),
.B1(n_286),
.B2(n_281),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_327),
.A2(n_330),
.B1(n_336),
.B2(n_312),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_331),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_314),
.B1(n_320),
.B2(n_297),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_267),
.Y(n_331)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_286),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_297),
.A2(n_283),
.B1(n_280),
.B2(n_266),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_304),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_339),
.C(n_310),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_267),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_295),
.A2(n_261),
.B(n_259),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_340),
.A2(n_293),
.B(n_318),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_317),
.Y(n_341)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_342),
.A2(n_294),
.B1(n_319),
.B2(n_263),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_262),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_343),
.B(n_306),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_301),
.B(n_313),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_346),
.Y(n_348)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_348),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_352),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_332),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_308),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_358),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_331),
.C(n_328),
.Y(n_375)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_344),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_359),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_325),
.B(n_299),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_324),
.A2(n_309),
.B1(n_306),
.B2(n_310),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_360),
.A2(n_366),
.B1(n_369),
.B2(n_294),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_361),
.A2(n_362),
.B(n_368),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_293),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_329),
.Y(n_377)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_365),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_363),
.B(n_329),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_375),
.Y(n_399)
);

AO221x1_ASAP7_75t_L g372 ( 
.A1(n_366),
.A2(n_330),
.B1(n_336),
.B2(n_311),
.C(n_337),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_374),
.Y(n_389)
);

BUFx12_ASAP7_75t_L g374 ( 
.A(n_367),
.Y(n_374)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_376),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_362),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_355),
.A2(n_350),
.B1(n_323),
.B2(n_351),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_386),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_339),
.C(n_364),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_381),
.C(n_384),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_347),
.C(n_340),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_342),
.C(n_323),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_341),
.C(n_326),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_391),
.Y(n_401)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_373),
.Y(n_390)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_381),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_382),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_395),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_361),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_379),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_354),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_394),
.Y(n_411)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_292),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_383),
.A2(n_348),
.B1(n_284),
.B2(n_315),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_400),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_387),
.A2(n_384),
.B1(n_377),
.B2(n_289),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_403),
.A2(n_405),
.B1(n_409),
.B2(n_394),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_404),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_375),
.B1(n_269),
.B2(n_315),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_370),
.C(n_270),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_407),
.B(n_410),
.Y(n_417)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_408),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_398),
.B(n_273),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_285),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g416 ( 
.A(n_412),
.B(n_399),
.Y(n_416)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_407),
.B(n_391),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_415),
.B(n_418),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_416),
.B(n_419),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_405),
.A2(n_403),
.B(n_406),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_411),
.A2(n_393),
.B(n_388),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_401),
.A2(n_400),
.B(n_374),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_422),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_401),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_409),
.Y(n_423)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_423),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_374),
.C(n_285),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_427),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_185),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_426),
.A2(n_417),
.B(n_415),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_431),
.A2(n_432),
.B(n_425),
.Y(n_434)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_425),
.Y(n_432)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_434),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_429),
.C(n_428),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_435),
.C(n_433),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_282),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_291),
.Y(n_439)
);


endmodule