module fake_jpeg_28512_n_69 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

AND2x2_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_22),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_0),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_1),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_30),
.B1(n_26),
.B2(n_7),
.Y(n_46)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_1),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx24_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_10),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_15),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_54),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_13),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_14),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_39),
.B(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_55),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_57),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_16),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_50),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_62),
.C(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_48),
.Y(n_69)
);


endmodule