module fake_jpeg_8833_n_178 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

HAxp5_ASAP7_75t_SL g27 ( 
.A(n_15),
.B(n_0),
.CON(n_27),
.SN(n_27)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_23),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_1),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_21),
.B1(n_18),
.B2(n_23),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_21),
.B1(n_20),
.B2(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_3),
.C(n_4),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_18),
.B1(n_32),
.B2(n_14),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_58),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_13),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_65),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_34),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_64),
.A2(n_14),
.B(n_26),
.Y(n_93)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_24),
.B1(n_20),
.B2(n_17),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_13),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_72),
.Y(n_82)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_33),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_31),
.C(n_30),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_32),
.C(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_93),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_84),
.C(n_32),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_94),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_30),
.B1(n_18),
.B2(n_17),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_92),
.B1(n_57),
.B2(n_51),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_73),
.B(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_93),
.B(n_25),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_31),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_64),
.B1(n_49),
.B2(n_18),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_97),
.B(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_106),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_19),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_104),
.C(n_113),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AO22x1_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_51),
.B1(n_52),
.B2(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_74),
.A3(n_94),
.B1(n_89),
.B2(n_16),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_75),
.B(n_25),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_11),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_11),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_19),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_3),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_5),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_78),
.C(n_90),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_120),
.B(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

AOI221xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_109),
.B1(n_115),
.B2(n_96),
.C(n_113),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_80),
.B1(n_77),
.B2(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_6),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_116),
.C(n_122),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_104),
.C(n_103),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_141),
.C(n_144),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_147),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_120),
.Y(n_146)
);

XNOR2x1_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_149),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_SL g147 ( 
.A(n_143),
.B(n_123),
.C(n_131),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_123),
.B(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_125),
.B1(n_116),
.B2(n_121),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_122),
.B1(n_132),
.B2(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_152),
.B(n_130),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_159),
.Y(n_162)
);

AO221x1_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_91),
.B1(n_54),
.B2(n_137),
.C(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_138),
.C(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_161),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_150),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_166),
.B1(n_167),
.B2(n_165),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_9),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_154),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_6),
.B1(n_16),
.B2(n_10),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_169),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_156),
.C(n_159),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_154),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_170),
.B(n_16),
.Y(n_175)
);

AOI31xp67_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_176),
.A3(n_12),
.B(n_6),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_9),
.B(n_10),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_172),
.Y(n_178)
);


endmodule