module fake_jpeg_15143_n_237 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_14),
.Y(n_50)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_28),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_41),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_50),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_21),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_37),
.B1(n_36),
.B2(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_14),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_27),
.B1(n_17),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_16),
.B1(n_25),
.B2(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_27),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_27),
.B1(n_17),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_59),
.B1(n_45),
.B2(n_16),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_17),
.B1(n_20),
.B2(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_70),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_54),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_65),
.B(n_68),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_18),
.B1(n_24),
.B2(n_20),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_72),
.B1(n_52),
.B2(n_25),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_74),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_41),
.C(n_40),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_85),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_54),
.B1(n_48),
.B2(n_41),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_84),
.B1(n_90),
.B2(n_59),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_49),
.B1(n_40),
.B2(n_42),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_51),
.A3(n_39),
.B1(n_48),
.B2(n_55),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_69),
.A3(n_58),
.B1(n_71),
.B2(n_65),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_42),
.B1(n_45),
.B2(n_53),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_92),
.B1(n_72),
.B2(n_26),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_16),
.B1(n_22),
.B2(n_19),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_103),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_67),
.B1(n_70),
.B2(n_64),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_107),
.B1(n_110),
.B2(n_56),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_113),
.B(n_78),
.Y(n_126)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_71),
.B1(n_67),
.B2(n_61),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_81),
.B1(n_67),
.B2(n_87),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_76),
.C(n_79),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_123),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_118),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_130),
.B1(n_113),
.B2(n_104),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_89),
.B(n_78),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_100),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_95),
.B(n_64),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_129),
.B(n_125),
.Y(n_144)
);

OR2x4_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_58),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_22),
.B(n_19),
.Y(n_131)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_56),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_143),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_114),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_114),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_141),
.B(n_136),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_152),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_110),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_103),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_43),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_121),
.B1(n_135),
.B2(n_130),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_121),
.B1(n_132),
.B2(n_124),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_133),
.B1(n_124),
.B2(n_119),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_119),
.B1(n_120),
.B2(n_123),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_164),
.B(n_168),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_152),
.B(n_145),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_148),
.A2(n_116),
.B1(n_107),
.B2(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_43),
.B1(n_1),
.B2(n_2),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_55),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_155),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_140),
.A2(n_147),
.B(n_146),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_138),
.B(n_26),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_176),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_137),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_179),
.C(n_35),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_146),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_142),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_163),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_22),
.B1(n_15),
.B2(n_26),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_172),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_185),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_19),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_55),
.C(n_35),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_157),
.C(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_169),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_167),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_55),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_188),
.Y(n_199)
);

FAx1_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_156),
.CI(n_159),
.CON(n_189),
.SN(n_189)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_169),
.B1(n_157),
.B2(n_168),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_195),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_197),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_184),
.B1(n_186),
.B2(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_200),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_30),
.C(n_43),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_188),
.B1(n_175),
.B2(n_177),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_1),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_181),
.B(n_15),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_189),
.B(n_8),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_7),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_7),
.B1(n_12),
.B2(n_3),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_201),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_200),
.C(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_215),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_189),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_209),
.B1(n_202),
.B2(n_207),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_211),
.C(n_206),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_211),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_6),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_219),
.A3(n_214),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_223),
.B1(n_212),
.B2(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_217),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_224),
.A2(n_8),
.B(n_9),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_227),
.B(n_8),
.C(n_10),
.Y(n_232)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_221),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_30),
.B(n_10),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_232),
.C(n_225),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_234),
.B(n_10),
.Y(n_235)
);

O2A1O1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_235),
.A2(n_2),
.B(n_11),
.C(n_219),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_2),
.B1(n_11),
.B2(n_219),
.Y(n_237)
);


endmodule