module fake_jpeg_8_n_184 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_184);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_14),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_59),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_SL g90 ( 
.A(n_73),
.Y(n_90)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_57),
.B(n_56),
.C(n_52),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_101),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_78),
.B1(n_61),
.B2(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_108),
.B1(n_17),
.B2(n_47),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_74),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_109),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_89),
.A2(n_61),
.B1(n_70),
.B2(n_75),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_53),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_48),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_72),
.B1(n_64),
.B2(n_70),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_118),
.B1(n_4),
.B2(n_5),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_85),
.B1(n_76),
.B2(n_48),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_124),
.B1(n_131),
.B2(n_8),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_64),
.B1(n_68),
.B2(n_55),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_99),
.C(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_51),
.B1(n_74),
.B2(n_50),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_128),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_22),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_19),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_5),
.C(n_6),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_74),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_10),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_24),
.C(n_44),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_150),
.C(n_25),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_141),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_6),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_142),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_8),
.B(n_9),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_16),
.B(n_23),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_9),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_10),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_11),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_149),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_12),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_15),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_133),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_26),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_160),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_28),
.C(n_30),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_31),
.A3(n_33),
.B1(n_36),
.B2(n_40),
.C1(n_42),
.C2(n_43),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_161),
.B(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_132),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_169),
.C(n_150),
.Y(n_170)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_153),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_163),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_156),
.C(n_160),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_177),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_171),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_169),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_172),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_155),
.Y(n_181)
);

NAND2x1_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_178),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_159),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_165),
.Y(n_184)
);


endmodule