module fake_jpeg_28348_n_195 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_195);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_33),
.Y(n_47)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_15),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_16),
.B(n_11),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_24),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_32),
.B1(n_18),
.B2(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_24),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_25),
.B1(n_29),
.B2(n_31),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_62),
.B1(n_26),
.B2(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_23),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_25),
.B1(n_26),
.B2(n_19),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_22),
.B1(n_23),
.B2(n_18),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_44),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_42),
.B(n_19),
.C(n_22),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_72),
.B1(n_62),
.B2(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_70),
.Y(n_88)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_71),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_78),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_27),
.B(n_20),
.C(n_19),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_60),
.B(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_58),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_81),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_84),
.Y(n_96)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_44),
.B(n_10),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_89),
.B1(n_95),
.B2(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_63),
.B1(n_51),
.B2(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_97),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_60),
.B(n_52),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_101),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_26),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_106),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_82),
.C(n_79),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_111),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_91),
.CI(n_90),
.CON(n_129),
.SN(n_129)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_66),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_74),
.B1(n_69),
.B2(n_83),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_116),
.B1(n_123),
.B2(n_124),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_75),
.B1(n_47),
.B2(n_31),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_20),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_126),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_9),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_121),
.B(n_86),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_20),
.B1(n_71),
.B2(n_2),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_48),
.B1(n_80),
.B2(n_2),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_103),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_9),
.C(n_1),
.Y(n_126)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_118),
.B(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_132),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_87),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_122),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_144),
.B1(n_132),
.B2(n_131),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_86),
.B1(n_113),
.B2(n_100),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_120),
.B(n_96),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_117),
.C(n_111),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_154),
.C(n_158),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_143),
.B(n_129),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_134),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_142),
.C(n_130),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_100),
.C(n_107),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_166),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_148),
.C(n_153),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_141),
.C(n_133),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_165),
.C(n_167),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_137),
.B1(n_133),
.B2(n_87),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_164),
.A2(n_169),
.B1(n_5),
.B2(n_6),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_137),
.C(n_104),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_0),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_3),
.C(n_4),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_5),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_155),
.B(n_157),
.C(n_150),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_175),
.Y(n_184)
);

XOR2x2_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_157),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_172),
.C(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_6),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_184),
.B(n_171),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_181),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_165),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_8),
.B1(n_171),
.B2(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_182),
.B(n_183),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_175),
.B(n_8),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_179),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_188),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_191),
.C(n_187),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_192),
.Y(n_195)
);


endmodule