module fake_jpeg_27444_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_18),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_20),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_18),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_24),
.B1(n_18),
.B2(n_15),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_14),
.B1(n_15),
.B2(n_12),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_18),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_10),
.Y(n_37)
);

AO21x1_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_38),
.B(n_40),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_15),
.B(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_26),
.B1(n_9),
.B2(n_11),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_39),
.B1(n_36),
.B2(n_9),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_13),
.B(n_11),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_13),
.B(n_24),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_38),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_26),
.B1(n_9),
.B2(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_49),
.B1(n_12),
.B2(n_17),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_26),
.B1(n_9),
.B2(n_12),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_51),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_17),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_47),
.B(n_41),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_45),
.C(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_61),
.Y(n_66)
);

A2O1A1O1Ixp25_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_42),
.B(n_43),
.C(n_46),
.D(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_67),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_54),
.B1(n_52),
.B2(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_59),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_60),
.C(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_65),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_0),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_4),
.Y(n_76)
);

AOI31xp67_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_1),
.A3(n_2),
.B(n_3),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_4),
.C(n_5),
.Y(n_77)
);

XNOR2x2_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_73),
.Y(n_78)
);


endmodule