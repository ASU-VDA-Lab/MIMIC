module fake_jpeg_3793_n_215 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_34),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_42),
.Y(n_70)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_28),
.Y(n_61)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_51),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_61),
.B(n_75),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_31),
.B1(n_18),
.B2(n_15),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_63),
.A2(n_32),
.B1(n_21),
.B2(n_12),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_28),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_79),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_78),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_27),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_35),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_25),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_30),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_58),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_98),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_18),
.B1(n_15),
.B2(n_22),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_102),
.B1(n_114),
.B2(n_62),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_30),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_108),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_10),
.B(n_3),
.C(n_4),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_103),
.B(n_104),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_32),
.B(n_5),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_4),
.C(n_5),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_8),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_6),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_80),
.Y(n_125)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_62),
.B1(n_82),
.B2(n_76),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_59),
.A2(n_6),
.B1(n_7),
.B2(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_119),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_65),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_97),
.B(n_71),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_131),
.Y(n_143)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_95),
.A2(n_81),
.B1(n_68),
.B2(n_78),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_92),
.B1(n_112),
.B2(n_69),
.Y(n_151)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_92),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_135),
.A2(n_110),
.B(n_99),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_145),
.B(n_117),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_89),
.C(n_107),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_117),
.C(n_115),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_89),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_143),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_127),
.B1(n_123),
.B2(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_104),
.B1(n_103),
.B2(n_96),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_131),
.B1(n_123),
.B2(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_72),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_155),
.B1(n_144),
.B2(n_147),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_166),
.B1(n_152),
.B2(n_153),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_164),
.C(n_165),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_150),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_116),
.C(n_64),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_129),
.C(n_56),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_173),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_57),
.B(n_67),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_177),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_141),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_179),
.C(n_171),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_180),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_138),
.C(n_145),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_140),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_192),
.C(n_193),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_185),
.B(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_184),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_191),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_147),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_165),
.C(n_164),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_160),
.C(n_140),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_144),
.B1(n_148),
.B2(n_163),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_179),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_189),
.C(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_193),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_133),
.C(n_66),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_175),
.C(n_177),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_183),
.C(n_148),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_174),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_201),
.B(n_91),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_202),
.A2(n_201),
.B(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_203),
.B(n_204),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_206),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_98),
.B1(n_124),
.B2(n_6),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_198),
.A3(n_55),
.B1(n_72),
.B2(n_124),
.C1(n_100),
.C2(n_66),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_210),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);


endmodule