module fake_netlist_1_9694_n_39 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x4_ASAP7_75t_L g12 ( .A(n_4), .B(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_SL g14 ( .A(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
CKINVDCx16_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_16), .B(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_16), .B(n_0), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_14), .A2(n_10), .B(n_11), .Y(n_20) );
NOR2xp67_ASAP7_75t_L g21 ( .A(n_16), .B(n_1), .Y(n_21) );
OAI21x1_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_15), .B(n_12), .Y(n_22) );
AOI21xp5_ASAP7_75t_L g23 ( .A1(n_18), .A2(n_14), .B(n_12), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_21), .Y(n_24) );
BUFx3_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
OR2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_17), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_27), .B(n_25), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_19), .B1(n_13), .B2(n_12), .Y(n_29) );
INVxp67_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
AOI31xp33_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_13), .A3(n_15), .B(n_1), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_28), .B(n_2), .Y(n_32) );
AND2x4_ASAP7_75t_L g33 ( .A(n_30), .B(n_2), .Y(n_33) );
INVx5_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_32), .B(n_30), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
XNOR2xp5_ASAP7_75t_L g37 ( .A(n_35), .B(n_33), .Y(n_37) );
OAI22xp5_ASAP7_75t_SL g38 ( .A1(n_37), .A2(n_34), .B1(n_33), .B2(n_35), .Y(n_38) );
AOI22x1_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_34), .B1(n_36), .B2(n_37), .Y(n_39) );
endmodule