module fake_jpeg_25082_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_47),
.Y(n_51)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_16),
.Y(n_75)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_27),
.B1(n_22),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_27),
.B1(n_22),
.B2(n_32),
.Y(n_80)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_35),
.B1(n_19),
.B2(n_33),
.Y(n_65)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_35),
.B1(n_62),
.B2(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_67),
.Y(n_101)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_46),
.Y(n_102)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_17),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_82),
.Y(n_116)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_98),
.B1(n_115),
.B2(n_44),
.Y(n_122)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_86),
.Y(n_130)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_24),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_95),
.C(n_46),
.Y(n_118)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_94),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_22),
.B1(n_19),
.B2(n_33),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_90),
.B1(n_25),
.B2(n_26),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_20),
.B1(n_34),
.B2(n_16),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_24),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_96),
.B(n_104),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_17),
.B1(n_21),
.B2(n_18),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_100),
.B1(n_37),
.B2(n_47),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_56),
.B1(n_50),
.B2(n_62),
.Y(n_100)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_18),
.B1(n_21),
.B2(n_25),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_114),
.B1(n_21),
.B2(n_44),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_54),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_56),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_103),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_122),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_24),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_133),
.Y(n_149)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_121),
.B1(n_129),
.B2(n_87),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_59),
.B1(n_26),
.B2(n_25),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_95),
.B1(n_85),
.B2(n_79),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_31),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_142),
.B(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_29),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_78),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_88),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_80),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_31),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_96),
.B1(n_77),
.B2(n_85),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_147),
.A2(n_146),
.B1(n_117),
.B2(n_128),
.Y(n_199)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_15),
.C(n_14),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_150),
.B(n_158),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_156),
.B1(n_161),
.B2(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_154),
.B1(n_146),
.B2(n_117),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_121),
.A2(n_92),
.B1(n_104),
.B2(n_79),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_86),
.C(n_84),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_103),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_113),
.B1(n_111),
.B2(n_100),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_165),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_113),
.B1(n_105),
.B2(n_26),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_116),
.A2(n_23),
.B(n_13),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_167),
.B(n_142),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_23),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_23),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_174),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_29),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_28),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_172),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_28),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_99),
.B1(n_1),
.B2(n_3),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_175),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_127),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_124),
.B1(n_120),
.B2(n_139),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_13),
.C(n_4),
.Y(n_179)
);

OAI21x1_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_5),
.B(n_6),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_0),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_8),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_141),
.B1(n_120),
.B2(n_128),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_201),
.B1(n_204),
.B2(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_182),
.B(n_11),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_142),
.B(n_144),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_184),
.B(n_193),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_202),
.B1(n_207),
.B2(n_209),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_152),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_203),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_163),
.A3(n_155),
.B1(n_149),
.B2(n_157),
.C1(n_175),
.C2(n_167),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_171),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_198),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_200),
.B(n_9),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_125),
.B1(n_140),
.B2(n_138),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_158),
.A2(n_125),
.B1(n_140),
.B2(n_7),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_125),
.B1(n_6),
.B2(n_7),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_168),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_208),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_156),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_155),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_213),
.Y(n_219)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_148),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_230),
.B1(n_188),
.B2(n_202),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_165),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_197),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_169),
.C(n_172),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_225),
.C(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_170),
.Y(n_223)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_227),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_180),
.C(n_148),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_177),
.B1(n_174),
.B2(n_164),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_183),
.A2(n_9),
.B(n_11),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_234),
.B(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_194),
.B(n_9),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_11),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_239),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_187),
.A2(n_12),
.B1(n_203),
.B2(n_188),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_204),
.B1(n_181),
.B2(n_186),
.Y(n_244)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_258),
.B1(n_214),
.B2(n_221),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_246),
.A2(n_253),
.B(n_254),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_229),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_256),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_192),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_260),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_238),
.B1(n_218),
.B2(n_236),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_234),
.A2(n_184),
.B(n_212),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_216),
.A2(n_212),
.B(n_213),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_185),
.Y(n_257)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_232),
.B(n_227),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_217),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_197),
.C(n_191),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_228),
.C(n_224),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_185),
.Y(n_264)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_281),
.C(n_265),
.Y(n_293)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_271),
.Y(n_291)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

XOR2x2_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_241),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_246),
.B(n_259),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_217),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_275),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_223),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_230),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_244),
.B1(n_243),
.B2(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_222),
.B1(n_218),
.B2(n_252),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_248),
.B(n_189),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_233),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_262),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_287),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_292),
.B1(n_298),
.B2(n_274),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_299),
.B(n_235),
.Y(n_312)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_261),
.B1(n_256),
.B2(n_245),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_265),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_263),
.C(n_245),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_296),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_275),
.B1(n_277),
.B2(n_269),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_250),
.C(n_248),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_267),
.A2(n_250),
.B1(n_243),
.B2(n_240),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_266),
.A2(n_189),
.B(n_255),
.Y(n_299)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_282),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_304),
.B(n_306),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_309),
.C(n_310),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_278),
.B1(n_279),
.B2(n_274),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_198),
.B1(n_205),
.B2(n_239),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_226),
.B1(n_187),
.B2(n_231),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_312),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_302),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_301),
.A2(n_291),
.B(n_284),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_318),
.C(n_321),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_285),
.C(n_287),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_285),
.C(n_298),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_300),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_328),
.B(n_319),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_307),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_324),
.Y(n_331)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_308),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_306),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_315),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_317),
.A2(n_309),
.B1(n_310),
.B2(n_226),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_326),
.A2(n_315),
.B(n_292),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_327),
.B(n_325),
.C(n_326),
.D(n_209),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_331),
.B(n_237),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_333),
.B(n_210),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_182),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_12),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_12),
.Y(n_340)
);


endmodule