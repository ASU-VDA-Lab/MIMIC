module fake_jpeg_7896_n_46 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_SL g20 ( 
.A(n_19),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_25),
.B(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_12),
.B1(n_6),
.B2(n_7),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_1),
.C(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_10),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_40),
.B1(n_14),
.B2(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_36),
.B(n_33),
.Y(n_44)
);

AO21x1_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_34),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_17),
.Y(n_46)
);


endmodule