module fake_ariane_1483_n_895 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_895);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_895;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_840;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_795;
wire n_398;
wire n_210;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_677;
wire n_614;
wire n_222;
wire n_703;
wire n_478;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_644;
wire n_536;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_767;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_126),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_108),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_172),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_125),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_137),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_72),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_25),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_53),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_171),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_146),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_32),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_107),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_59),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_90),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_33),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_49),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_165),
.Y(n_228)
);

INVxp33_ASAP7_75t_R g229 ( 
.A(n_135),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_149),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_5),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_113),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_117),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_26),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_26),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_46),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_119),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_36),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_12),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_57),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_111),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_148),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_196),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_116),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_27),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_168),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_42),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_99),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_61),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_70),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_29),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_132),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_161),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_112),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_58),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_15),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_15),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_86),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_124),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_95),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_24),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_8),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_175),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_2),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_50),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_13),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_122),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_9),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_159),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_188),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_177),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_198),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_89),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_179),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_173),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_23),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_7),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_154),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_0),
.Y(n_285)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_211),
.B(n_0),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_1),
.Y(n_288)
);

BUFx8_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_208),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_220),
.B(n_1),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_225),
.B(n_2),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_214),
.B(n_28),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_268),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_208),
.B(n_3),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_204),
.B(n_31),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_262),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_221),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g302 ( 
.A(n_214),
.B(n_34),
.Y(n_302)
);

BUFx8_ASAP7_75t_SL g303 ( 
.A(n_217),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_221),
.B(n_3),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_262),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_237),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g307 ( 
.A(n_268),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_226),
.B(n_4),
.Y(n_308)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_232),
.B(n_5),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_227),
.B(n_6),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_230),
.B(n_239),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_212),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_243),
.B(n_6),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_247),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_235),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g325 ( 
.A(n_236),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_273),
.B(n_7),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_250),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_249),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_251),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_259),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_206),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_266),
.B(n_8),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_269),
.B1(n_275),
.B2(n_241),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_285),
.A2(n_272),
.B1(n_274),
.B2(n_205),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_207),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_323),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_209),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_306),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_210),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_281),
.B1(n_280),
.B2(n_279),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_288),
.A2(n_312),
.B1(n_287),
.B2(n_304),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_R g349 ( 
.A1(n_336),
.A2(n_308),
.B1(n_318),
.B2(n_294),
.Y(n_349)
);

AOI22x1_ASAP7_75t_L g350 ( 
.A1(n_298),
.A2(n_278),
.B1(n_277),
.B2(n_276),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_332),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_307),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g354 ( 
.A1(n_322),
.A2(n_331),
.B1(n_307),
.B2(n_328),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_291),
.B(n_213),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g356 ( 
.A1(n_298),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_298),
.A2(n_271),
.B1(n_270),
.B2(n_265),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_291),
.B(n_215),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g359 ( 
.A1(n_322),
.A2(n_263),
.B1(n_258),
.B2(n_257),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_216),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g362 ( 
.A1(n_331),
.A2(n_256),
.B1(n_255),
.B2(n_254),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g363 ( 
.A1(n_328),
.A2(n_253),
.B1(n_248),
.B2(n_246),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g364 ( 
.A1(n_325),
.A2(n_315),
.B1(n_295),
.B2(n_334),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_325),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_336),
.A2(n_245),
.B1(n_242),
.B2(n_240),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_316),
.A2(n_238),
.B1(n_234),
.B2(n_233),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_294),
.A2(n_231),
.B1(n_228),
.B2(n_224),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_321),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_303),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_308),
.A2(n_223),
.B1(n_222),
.B2(n_219),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_L g377 ( 
.A1(n_330),
.A2(n_218),
.B1(n_11),
.B2(n_12),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_289),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_303),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_318),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_335),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_L g382 ( 
.A1(n_330),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_301),
.B(n_18),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_335),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_L g385 ( 
.A1(n_334),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_290),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_335),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_335),
.A2(n_333),
.B1(n_329),
.B2(n_296),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_378),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_333),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_366),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_339),
.B(n_333),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_374),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_341),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_366),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_379),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_342),
.B(n_329),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_379),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_387),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

BUFx6f_ASAP7_75t_SL g407 ( 
.A(n_352),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_384),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_383),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_337),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_289),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_355),
.B(n_329),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_358),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_347),
.B(n_309),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_345),
.B(n_290),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_361),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_360),
.Y(n_419)
);

OR2x2_ASAP7_75t_SL g420 ( 
.A(n_354),
.B(n_289),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_342),
.B(n_292),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_365),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_309),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_373),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_369),
.B(n_309),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_368),
.B(n_309),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_386),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_381),
.Y(n_431)
);

AOI21x1_ASAP7_75t_L g432 ( 
.A1(n_356),
.A2(n_326),
.B(n_324),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_367),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_389),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_388),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_348),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_350),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_380),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_359),
.B(n_354),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_357),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_375),
.B(n_292),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_363),
.A2(n_302),
.B(n_296),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_382),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_R g449 ( 
.A(n_359),
.B(n_320),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_363),
.B(n_313),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_377),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_362),
.A2(n_302),
.B(n_296),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_339),
.B(n_320),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_344),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_342),
.B(n_296),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g459 ( 
.A1(n_376),
.A2(n_302),
.B(n_296),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_344),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_434),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_406),
.B(n_313),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_405),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_404),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

CKINVDCx6p67_ASAP7_75t_R g466 ( 
.A(n_407),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_22),
.Y(n_467)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_392),
.B(n_313),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_402),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_394),
.B(n_313),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_394),
.B(n_319),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_442),
.B(n_401),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_437),
.B(n_319),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_434),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_402),
.B(n_302),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_396),
.B(n_319),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_319),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_425),
.B(n_302),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_425),
.B(n_427),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_434),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_427),
.B(n_293),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_22),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_401),
.B(n_286),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_418),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_422),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_444),
.B(n_23),
.Y(n_488)
);

AND2x2_ASAP7_75t_SL g489 ( 
.A(n_441),
.B(n_293),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_24),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_435),
.B(n_293),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_457),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_413),
.B(n_293),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_460),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_419),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_434),
.Y(n_498)
);

NAND2x1p5_ASAP7_75t_L g499 ( 
.A(n_443),
.B(n_286),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_398),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_432),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_435),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_454),
.B(n_25),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_424),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_458),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_451),
.B(n_27),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_446),
.A2(n_300),
.B(n_286),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_444),
.B(n_35),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_447),
.B(n_305),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_413),
.B(n_305),
.Y(n_511)
);

NAND2x1p5_ASAP7_75t_L g512 ( 
.A(n_458),
.B(n_286),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_430),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_449),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_391),
.Y(n_515)
);

AND2x2_ASAP7_75t_SL g516 ( 
.A(n_454),
.B(n_305),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_448),
.B(n_305),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_459),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_454),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_456),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_408),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_421),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_450),
.B(n_300),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_445),
.B(n_300),
.Y(n_526)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_438),
.A2(n_37),
.B(n_38),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_417),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_431),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_395),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_450),
.B(n_300),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_436),
.B(n_203),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_439),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_461),
.B(n_440),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_433),
.Y(n_535)
);

AO21x2_ASAP7_75t_L g536 ( 
.A1(n_479),
.A2(n_446),
.B(n_455),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_428),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_428),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_484),
.B(n_429),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_469),
.B(n_415),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_481),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_481),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_484),
.B(n_490),
.Y(n_544)
);

AND2x2_ASAP7_75t_SL g545 ( 
.A(n_489),
.B(n_420),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_490),
.B(n_399),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_469),
.B(n_400),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_520),
.B(n_407),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_520),
.B(n_449),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_529),
.B(n_455),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_469),
.B(n_403),
.Y(n_551)
);

AND2x6_ASAP7_75t_L g552 ( 
.A(n_509),
.B(n_412),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_465),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_461),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_520),
.B(n_39),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_475),
.B(n_40),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_472),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_509),
.B(n_476),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_475),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_L g560 ( 
.A(n_502),
.B(n_41),
.Y(n_560)
);

AND2x2_ASAP7_75t_SL g561 ( 
.A(n_489),
.B(n_516),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_L g562 ( 
.A(n_502),
.B(n_43),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_530),
.B(n_44),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_530),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_493),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_529),
.B(n_45),
.Y(n_567)
);

BUFx4f_ASAP7_75t_L g568 ( 
.A(n_466),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_472),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_488),
.B(n_47),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_488),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_516),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_493),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_525),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_512),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_473),
.B(n_48),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_523),
.B(n_51),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_501),
.Y(n_578)
);

BUFx12f_ASAP7_75t_L g579 ( 
.A(n_488),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_482),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_501),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_464),
.Y(n_582)
);

OR2x6_ASAP7_75t_SL g583 ( 
.A(n_466),
.B(n_52),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_525),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_482),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_498),
.B(n_54),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_498),
.Y(n_589)
);

NAND2x1p5_ASAP7_75t_L g590 ( 
.A(n_506),
.B(n_55),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_512),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_467),
.B(n_56),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_564),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_572),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_564),
.Y(n_595)
);

INVx3_ASAP7_75t_SL g596 ( 
.A(n_551),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_582),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_591),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_591),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_582),
.Y(n_600)
);

INVx6_ASAP7_75t_L g601 ( 
.A(n_566),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_587),
.Y(n_602)
);

BUFx12f_ASAP7_75t_L g603 ( 
.A(n_551),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_537),
.B(n_521),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_568),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_566),
.B(n_509),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_549),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_568),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_587),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_572),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_542),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_558),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_549),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_572),
.Y(n_614)
);

NOR2xp67_ASAP7_75t_SL g615 ( 
.A(n_540),
.B(n_491),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_558),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_547),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_554),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_554),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_579),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_579),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_578),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_535),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_535),
.Y(n_625)
);

BUFx4_ASAP7_75t_SL g626 ( 
.A(n_570),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_570),
.B(n_506),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_544),
.B(n_521),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_558),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_538),
.B(n_507),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_542),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_552),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_578),
.Y(n_634)
);

CKINVDCx16_ASAP7_75t_R g635 ( 
.A(n_546),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_534),
.B(n_492),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_593),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_630),
.A2(n_545),
.B1(n_539),
.B2(n_561),
.Y(n_638)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_594),
.Y(n_639)
);

BUFx8_ASAP7_75t_SL g640 ( 
.A(n_605),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_624),
.A2(n_545),
.B1(n_561),
.B2(n_552),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_635),
.A2(n_558),
.B1(n_504),
.B2(n_584),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_594),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_605),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_593),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_611),
.Y(n_646)
);

BUFx8_ASAP7_75t_SL g647 ( 
.A(n_608),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_627),
.A2(n_570),
.B1(n_571),
.B2(n_569),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_595),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_611),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_625),
.A2(n_552),
.B1(n_558),
.B2(n_534),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_628),
.Y(n_652)
);

INVx6_ASAP7_75t_L g653 ( 
.A(n_594),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_627),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_631),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_L g656 ( 
.A1(n_627),
.A2(n_563),
.B1(n_592),
.B2(n_550),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_608),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_617),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_604),
.A2(n_552),
.B1(n_534),
.B2(n_507),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_635),
.B(n_517),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_618),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_627),
.A2(n_553),
.B1(n_557),
.B2(n_586),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_594),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_631),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_603),
.A2(n_552),
.B1(n_528),
.B2(n_581),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_595),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_632),
.A2(n_572),
.B1(n_576),
.B2(n_541),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_603),
.A2(n_528),
.B1(n_581),
.B2(n_527),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_618),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_632),
.A2(n_576),
.B1(n_541),
.B2(n_555),
.Y(n_670)
);

CKINVDCx11_ASAP7_75t_R g671 ( 
.A(n_596),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_619),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_619),
.Y(n_673)
);

CKINVDCx11_ASAP7_75t_R g674 ( 
.A(n_596),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_620),
.Y(n_675)
);

BUFx4f_ASAP7_75t_SL g676 ( 
.A(n_596),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_597),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_620),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_633),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_677),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_652),
.B(n_633),
.Y(n_681)
);

AOI222xp33_ASAP7_75t_L g682 ( 
.A1(n_638),
.A2(n_523),
.B1(n_494),
.B2(n_496),
.C1(n_636),
.C2(n_622),
.Y(n_682)
);

OAI22xp33_ASAP7_75t_L g683 ( 
.A1(n_642),
.A2(n_583),
.B1(n_626),
.B2(n_612),
.Y(n_683)
);

INVx5_ASAP7_75t_SL g684 ( 
.A(n_643),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_SL g685 ( 
.A1(n_656),
.A2(n_548),
.B(n_555),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_SL g686 ( 
.A1(n_656),
.A2(n_548),
.B(n_590),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_670),
.A2(n_590),
.B(n_588),
.Y(n_687)
);

INVx5_ASAP7_75t_SL g688 ( 
.A(n_643),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_638),
.A2(n_606),
.B1(n_636),
.B2(n_607),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_650),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_676),
.A2(n_606),
.B1(n_612),
.B2(n_574),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_668),
.A2(n_471),
.B(n_470),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_640),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_SL g694 ( 
.A1(n_641),
.A2(n_588),
.B(n_556),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_SL g695 ( 
.A1(n_659),
.A2(n_668),
.B(n_662),
.Y(n_695)
);

OAI222xp33_ASAP7_75t_L g696 ( 
.A1(n_659),
.A2(n_607),
.B1(n_613),
.B2(n_615),
.C1(n_606),
.C2(n_636),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_660),
.A2(n_606),
.B1(n_636),
.B2(n_613),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_679),
.B(n_621),
.Y(n_698)
);

OAI21xp33_ASAP7_75t_L g699 ( 
.A1(n_662),
.A2(n_615),
.B(n_532),
.Y(n_699)
);

OAI222xp33_ASAP7_75t_L g700 ( 
.A1(n_667),
.A2(n_629),
.B1(n_634),
.B2(n_623),
.C1(n_597),
.C2(n_602),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_658),
.B(n_600),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_676),
.A2(n_612),
.B1(n_629),
.B2(n_616),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_664),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_651),
.A2(n_526),
.B1(n_463),
.B2(n_474),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_669),
.B(n_577),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_673),
.B(n_610),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_647),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_648),
.A2(n_616),
.B1(n_533),
.B2(n_556),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_651),
.A2(n_463),
.B1(n_474),
.B2(n_500),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_678),
.B(n_533),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_661),
.B(n_610),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_661),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_665),
.A2(n_500),
.B1(n_565),
.B2(n_573),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_665),
.A2(n_616),
.B1(n_533),
.B2(n_567),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_644),
.A2(n_522),
.B1(n_601),
.B2(n_468),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_643),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_675),
.B(n_562),
.C(n_560),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_646),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_643),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_644),
.A2(n_522),
.B1(n_601),
.B2(n_575),
.Y(n_720)
);

BUFx12f_ASAP7_75t_L g721 ( 
.A(n_671),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_657),
.B(n_600),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_646),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_672),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_655),
.A2(n_543),
.B1(n_565),
.B2(n_573),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_663),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_674),
.B(n_614),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_695),
.A2(n_637),
.B1(n_645),
.B2(n_666),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_682),
.A2(n_683),
.B1(n_699),
.B2(n_689),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_683),
.A2(n_709),
.B1(n_704),
.B2(n_692),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_698),
.B(n_649),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_SL g732 ( 
.A1(n_708),
.A2(n_562),
.B1(n_560),
.B2(n_654),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_697),
.A2(n_543),
.B1(n_497),
.B2(n_513),
.Y(n_733)
);

AOI221xp5_ASAP7_75t_L g734 ( 
.A1(n_685),
.A2(n_497),
.B1(n_505),
.B2(n_513),
.C(n_462),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_SL g735 ( 
.A1(n_724),
.A2(n_594),
.B1(n_599),
.B2(n_598),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_690),
.A2(n_505),
.B1(n_602),
.B2(n_634),
.Y(n_736)
);

AOI221xp5_ASAP7_75t_L g737 ( 
.A1(n_681),
.A2(n_462),
.B1(n_518),
.B2(n_510),
.C(n_515),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_712),
.B(n_655),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_706),
.B(n_663),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_703),
.A2(n_623),
.B1(n_609),
.B2(n_478),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_680),
.A2(n_609),
.B1(n_478),
.B2(n_580),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_705),
.A2(n_580),
.B1(n_585),
.B2(n_589),
.Y(n_742)
);

OAI21xp33_ASAP7_75t_L g743 ( 
.A1(n_686),
.A2(n_483),
.B(n_477),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_713),
.A2(n_585),
.B1(n_589),
.B2(n_580),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_723),
.A2(n_585),
.B1(n_589),
.B2(n_580),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_701),
.A2(n_589),
.B1(n_585),
.B2(n_515),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_694),
.A2(n_601),
.B1(n_653),
.B2(n_639),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_SL g748 ( 
.A1(n_717),
.A2(n_654),
.B1(n_601),
.B2(n_614),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_711),
.B(n_663),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_718),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_687),
.A2(n_710),
.B1(n_691),
.B2(n_702),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_714),
.A2(n_487),
.B1(n_486),
.B2(n_510),
.Y(n_752)
);

OAI222xp33_ASAP7_75t_L g753 ( 
.A1(n_722),
.A2(n_598),
.B1(n_599),
.B2(n_518),
.C1(n_499),
.C2(n_524),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_720),
.A2(n_575),
.B1(n_598),
.B2(n_599),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_725),
.A2(n_486),
.B1(n_487),
.B2(n_470),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_716),
.B(n_719),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_721),
.A2(n_536),
.B1(n_487),
.B2(n_486),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_715),
.A2(n_471),
.B1(n_531),
.B2(n_536),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_727),
.A2(n_499),
.B1(n_485),
.B2(n_476),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_700),
.A2(n_653),
.B1(n_639),
.B2(n_663),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_726),
.B(n_495),
.C(n_511),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_726),
.A2(n_499),
.B1(n_476),
.B2(n_653),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_716),
.A2(n_639),
.B1(n_492),
.B2(n_508),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_719),
.A2(n_684),
.B1(n_688),
.B2(n_707),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_693),
.A2(n_492),
.B1(n_512),
.B2(n_519),
.Y(n_765)
);

OAI221xp5_ASAP7_75t_L g766 ( 
.A1(n_700),
.A2(n_519),
.B1(n_502),
.B2(n_63),
.C(n_64),
.Y(n_766)
);

OAI221xp5_ASAP7_75t_L g767 ( 
.A1(n_729),
.A2(n_696),
.B1(n_502),
.B2(n_684),
.C(n_688),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_738),
.B(n_684),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_749),
.B(n_688),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_739),
.B(n_60),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_756),
.B(n_62),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_750),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_751),
.B(n_65),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_729),
.B(n_66),
.Y(n_774)
);

OAI21xp33_ASAP7_75t_L g775 ( 
.A1(n_766),
.A2(n_502),
.B(n_696),
.Y(n_775)
);

NOR2xp67_ASAP7_75t_L g776 ( 
.A(n_728),
.B(n_67),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_742),
.B(n_68),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_SL g778 ( 
.A1(n_747),
.A2(n_69),
.B(n_71),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_731),
.B(n_742),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_757),
.B(n_202),
.Y(n_780)
);

OAI21xp33_ASAP7_75t_SL g781 ( 
.A1(n_730),
.A2(n_73),
.B(n_74),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_757),
.B(n_75),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_730),
.B(n_200),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_743),
.B(n_76),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_735),
.B(n_199),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_734),
.B(n_77),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_754),
.B(n_195),
.Y(n_787)
);

NAND2x1_ASAP7_75t_L g788 ( 
.A(n_764),
.B(n_78),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_760),
.B(n_194),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_765),
.B(n_748),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_740),
.B(n_79),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_761),
.B(n_80),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_758),
.B(n_81),
.C(n_82),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_779),
.B(n_732),
.Y(n_794)
);

AO21x2_ASAP7_75t_L g795 ( 
.A1(n_780),
.A2(n_753),
.B(n_746),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_768),
.B(n_752),
.Y(n_796)
);

AOI221xp5_ASAP7_75t_L g797 ( 
.A1(n_784),
.A2(n_737),
.B1(n_741),
.B2(n_759),
.C(n_733),
.Y(n_797)
);

AOI211xp5_ASAP7_75t_L g798 ( 
.A1(n_773),
.A2(n_83),
.B(n_84),
.C(n_85),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_772),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_776),
.A2(n_775),
.B1(n_774),
.B2(n_767),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_769),
.B(n_745),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_771),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_790),
.Y(n_803)
);

AOI211xp5_ASAP7_75t_L g804 ( 
.A1(n_781),
.A2(n_778),
.B(n_784),
.C(n_792),
.Y(n_804)
);

AOI221xp5_ASAP7_75t_L g805 ( 
.A1(n_783),
.A2(n_736),
.B1(n_755),
.B2(n_762),
.C(n_763),
.Y(n_805)
);

OAI211xp5_ASAP7_75t_SL g806 ( 
.A1(n_786),
.A2(n_744),
.B(n_88),
.C(n_91),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_785),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_770),
.B(n_87),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_787),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_792),
.B(n_92),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_807),
.B(n_788),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_802),
.B(n_782),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_809),
.B(n_778),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_810),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_799),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_794),
.B(n_777),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_801),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_802),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_801),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_803),
.B(n_791),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_SL g821 ( 
.A(n_806),
.B(n_793),
.C(n_789),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_796),
.B(n_93),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_811),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_819),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_815),
.Y(n_825)
);

INVx8_ASAP7_75t_L g826 ( 
.A(n_822),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_814),
.Y(n_827)
);

CKINVDCx8_ASAP7_75t_R g828 ( 
.A(n_813),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_825),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_823),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_826),
.Y(n_831)
);

OA22x2_ASAP7_75t_L g832 ( 
.A1(n_824),
.A2(n_819),
.B1(n_814),
.B2(n_817),
.Y(n_832)
);

OA22x2_ASAP7_75t_L g833 ( 
.A1(n_827),
.A2(n_816),
.B1(n_820),
.B2(n_818),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_830),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_831),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_829),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_833),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_834),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_837),
.A2(n_828),
.B1(n_832),
.B2(n_813),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_SL g840 ( 
.A1(n_835),
.A2(n_804),
.B1(n_800),
.B2(n_826),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_836),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_838),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_841),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_840),
.Y(n_844)
);

OA22x2_ASAP7_75t_L g845 ( 
.A1(n_839),
.A2(n_818),
.B1(n_810),
.B2(n_815),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_842),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_844),
.A2(n_821),
.B1(n_800),
.B2(n_795),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_845),
.A2(n_821),
.B1(n_812),
.B2(n_798),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_SL g849 ( 
.A1(n_843),
.A2(n_795),
.B1(n_797),
.B2(n_808),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_844),
.A2(n_808),
.B1(n_805),
.B2(n_97),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_842),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_844),
.B(n_94),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_846),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_847),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_851),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_852),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_850),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_848),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_849),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_856),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_858),
.A2(n_109),
.B1(n_110),
.B2(n_114),
.Y(n_861)
);

AND4x1_ASAP7_75t_L g862 ( 
.A(n_853),
.B(n_115),
.C(n_120),
.D(n_121),
.Y(n_862)
);

NOR2x1_ASAP7_75t_L g863 ( 
.A(n_855),
.B(n_123),
.Y(n_863)
);

AND4x1_ASAP7_75t_L g864 ( 
.A(n_854),
.B(n_127),
.C(n_128),
.D(n_129),
.Y(n_864)
);

NAND4xp25_ASAP7_75t_L g865 ( 
.A(n_859),
.B(n_130),
.C(n_131),
.D(n_133),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_857),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_866)
);

NOR4xp75_ASAP7_75t_L g867 ( 
.A(n_858),
.B(n_139),
.C(n_140),
.D(n_141),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_863),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_860),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_867),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_861),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_862),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_865),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_864),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_866),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_863),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_868),
.A2(n_145),
.B1(n_147),
.B2(n_150),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_869),
.A2(n_151),
.B1(n_153),
.B2(n_155),
.Y(n_878)
);

AO22x2_ASAP7_75t_L g879 ( 
.A1(n_872),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_873),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_870),
.A2(n_169),
.B1(n_170),
.B2(n_174),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_873),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_882),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_879),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_880),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_878),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_881),
.Y(n_887)
);

AO22x2_ASAP7_75t_L g888 ( 
.A1(n_884),
.A2(n_874),
.B1(n_871),
.B2(n_875),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_883),
.A2(n_876),
.B1(n_877),
.B2(n_180),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_885),
.A2(n_193),
.B1(n_178),
.B2(n_181),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_888),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_891),
.A2(n_889),
.B1(n_887),
.B2(n_886),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_892),
.Y(n_893)
);

AOI221x1_ASAP7_75t_L g894 ( 
.A1(n_893),
.A2(n_890),
.B1(n_182),
.B2(n_183),
.C(n_184),
.Y(n_894)
);

AOI211xp5_ASAP7_75t_L g895 ( 
.A1(n_894),
.A2(n_176),
.B(n_185),
.C(n_186),
.Y(n_895)
);


endmodule