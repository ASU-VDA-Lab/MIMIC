module real_aes_11875_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_1380;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_1352;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVxp33_ASAP7_75t_L g852 ( .A(n_0), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_0), .A2(n_28), .B1(n_535), .B2(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_2), .A2(n_203), .B1(n_394), .B2(n_536), .Y(n_956) );
INVxp33_ASAP7_75t_L g977 ( .A(n_2), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_3), .A2(n_9), .B1(n_303), .B2(n_304), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_3), .A2(n_9), .B1(n_393), .B2(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g737 ( .A(n_4), .Y(n_737) );
INVx1_ASAP7_75t_L g997 ( .A(n_5), .Y(n_997) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_6), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_6), .B(n_179), .Y(n_268) );
INVx1_ASAP7_75t_L g311 ( .A(n_6), .Y(n_311) );
AND2x2_ASAP7_75t_L g319 ( .A(n_6), .B(n_310), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_7), .A2(n_10), .B1(n_484), .B2(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g942 ( .A(n_7), .Y(n_942) );
INVxp67_ASAP7_75t_L g859 ( .A(n_8), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_8), .A2(n_74), .B1(n_529), .B2(n_535), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_10), .A2(n_112), .B1(n_937), .B2(n_939), .C(n_941), .Y(n_936) );
INVx1_ASAP7_75t_L g1253 ( .A(n_11), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_12), .A2(n_103), .B1(n_552), .B2(n_554), .Y(n_551) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_12), .Y(n_613) );
INVxp33_ASAP7_75t_L g1083 ( .A(n_13), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g1114 ( .A1(n_13), .A2(n_131), .B1(n_748), .B2(n_886), .C(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g561 ( .A(n_14), .Y(n_561) );
AO221x2_ASAP7_75t_L g1162 ( .A1(n_15), .A2(n_56), .B1(n_1139), .B2(n_1161), .C(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1180 ( .A(n_16), .Y(n_1180) );
INVx1_ASAP7_75t_L g1385 ( .A(n_17), .Y(n_1385) );
OR2x2_ASAP7_75t_L g338 ( .A(n_18), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g369 ( .A(n_18), .Y(n_369) );
INVx1_ASAP7_75t_L g1119 ( .A(n_19), .Y(n_1119) );
INVx1_ASAP7_75t_L g1164 ( .A(n_20), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_21), .A2(n_220), .B1(n_483), .B2(n_485), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_21), .A2(n_220), .B1(n_290), .B2(n_505), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_22), .Y(n_1021) );
INVx1_ASAP7_75t_L g556 ( .A(n_23), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_24), .A2(n_129), .B1(n_533), .B2(n_535), .Y(n_532) );
INVxp33_ASAP7_75t_SL g581 ( .A(n_24), .Y(n_581) );
OR2x2_ASAP7_75t_L g267 ( .A(n_25), .B(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g283 ( .A(n_25), .Y(n_283) );
INVx1_ASAP7_75t_L g318 ( .A(n_25), .Y(n_318) );
BUFx2_ASAP7_75t_L g476 ( .A(n_25), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_26), .A2(n_156), .B1(n_584), .B2(n_590), .C(n_593), .Y(n_712) );
OAI22xp33_ASAP7_75t_SL g753 ( .A1(n_26), .A2(n_156), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g1251 ( .A(n_27), .Y(n_1251) );
INVxp33_ASAP7_75t_L g848 ( .A(n_28), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_29), .A2(n_144), .B1(n_293), .B2(n_513), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_29), .A2(n_144), .B1(n_692), .B2(n_693), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_30), .A2(n_113), .B1(n_290), .B2(n_315), .C(n_597), .Y(n_660) );
INVx1_ASAP7_75t_L g687 ( .A(n_30), .Y(n_687) );
INVx1_ASAP7_75t_L g809 ( .A(n_31), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_32), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_33), .A2(n_162), .B1(n_549), .B2(n_761), .C(n_786), .Y(n_785) );
INVxp33_ASAP7_75t_SL g829 ( .A(n_33), .Y(n_829) );
INVxp33_ASAP7_75t_L g416 ( .A(n_34), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_34), .A2(n_38), .B1(n_290), .B2(n_505), .Y(n_514) );
AOI22xp33_ASAP7_75t_SL g305 ( .A1(n_35), .A2(n_72), .B1(n_286), .B2(n_290), .Y(n_305) );
INVx1_ASAP7_75t_L g390 ( .A(n_35), .Y(n_390) );
INVxp33_ASAP7_75t_L g709 ( .A(n_36), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_36), .A2(n_39), .B1(n_744), .B2(n_746), .C(n_748), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_37), .A2(n_112), .B1(n_549), .B2(n_761), .C(n_885), .Y(n_912) );
INVx1_ASAP7_75t_L g943 ( .A(n_37), .Y(n_943) );
INVxp67_ASAP7_75t_L g435 ( .A(n_38), .Y(n_435) );
INVxp33_ASAP7_75t_L g707 ( .A(n_39), .Y(n_707) );
CKINVDCx16_ASAP7_75t_R g894 ( .A(n_40), .Y(n_894) );
INVx1_ASAP7_75t_L g1247 ( .A(n_41), .Y(n_1247) );
OAI221xp5_ASAP7_75t_SL g952 ( .A1(n_42), .A2(n_197), .B1(n_542), .B2(n_754), .C(n_953), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_42), .A2(n_197), .B1(n_590), .B2(n_819), .C(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1096 ( .A(n_43), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_44), .Y(n_948) );
INVxp33_ASAP7_75t_SL g710 ( .A(n_45), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_45), .A2(n_219), .B1(n_492), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g285 ( .A1(n_46), .A2(n_187), .B1(n_286), .B2(n_290), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_46), .A2(n_154), .B1(n_352), .B2(n_359), .Y(n_351) );
INVx1_ASAP7_75t_L g735 ( .A(n_47), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g960 ( .A1(n_48), .A2(n_134), .B1(n_961), .B2(n_963), .C(n_966), .Y(n_960) );
INVxp67_ASAP7_75t_SL g989 ( .A(n_48), .Y(n_989) );
INVx1_ASAP7_75t_L g563 ( .A(n_49), .Y(n_563) );
AOI221xp5_ASAP7_75t_SL g907 ( .A1(n_50), .A2(n_65), .B1(n_531), .B2(n_746), .C(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g924 ( .A(n_50), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_51), .A2(n_175), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
INVx1_ASAP7_75t_L g1058 ( .A(n_51), .Y(n_1058) );
INVx1_ASAP7_75t_L g904 ( .A(n_52), .Y(n_904) );
INVx1_ASAP7_75t_L g784 ( .A(n_53), .Y(n_784) );
INVx1_ASAP7_75t_L g676 ( .A(n_54), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_54), .A2(n_135), .B1(n_692), .B2(n_699), .Y(n_698) );
INVxp33_ASAP7_75t_L g472 ( .A(n_55), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_55), .A2(n_125), .B1(n_391), .B2(n_483), .Y(n_494) );
XNOR2x2_ASAP7_75t_L g259 ( .A(n_56), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g903 ( .A(n_57), .Y(n_903) );
INVx1_ASAP7_75t_L g959 ( .A(n_58), .Y(n_959) );
INVxp67_ASAP7_75t_L g469 ( .A(n_59), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_59), .A2(n_79), .B1(n_496), .B2(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g1189 ( .A(n_60), .Y(n_1189) );
AOI22xp33_ASAP7_75t_SL g292 ( .A1(n_61), .A2(n_154), .B1(n_293), .B2(n_298), .Y(n_292) );
AOI21xp33_ASAP7_75t_L g363 ( .A1(n_61), .A2(n_364), .B(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g427 ( .A(n_62), .Y(n_427) );
CKINVDCx16_ASAP7_75t_R g1194 ( .A(n_63), .Y(n_1194) );
INVxp33_ASAP7_75t_SL g1348 ( .A(n_64), .Y(n_1348) );
AOI221xp5_ASAP7_75t_L g1378 ( .A1(n_64), .A2(n_221), .B1(n_1375), .B2(n_1379), .C(n_1380), .Y(n_1378) );
INVx1_ASAP7_75t_L g922 ( .A(n_65), .Y(n_922) );
INVxp67_ASAP7_75t_L g857 ( .A(n_66), .Y(n_857) );
AOI221xp5_ASAP7_75t_L g884 ( .A1(n_66), .A2(n_159), .B1(n_549), .B2(n_885), .C(n_886), .Y(n_884) );
INVxp33_ASAP7_75t_L g422 ( .A(n_67), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_67), .A2(n_85), .B1(n_507), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g1147 ( .A(n_68), .Y(n_1147) );
INVx1_ASAP7_75t_L g803 ( .A(n_69), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_70), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_71), .A2(n_192), .B1(n_899), .B2(n_900), .C(n_901), .Y(n_898) );
INVx1_ASAP7_75t_L g934 ( .A(n_71), .Y(n_934) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_72), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g331 ( .A(n_73), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_73), .A2(n_123), .B1(n_359), .B2(n_364), .Y(n_373) );
INVxp67_ASAP7_75t_L g862 ( .A(n_74), .Y(n_862) );
XNOR2xp5_ASAP7_75t_L g627 ( .A(n_75), .B(n_628), .Y(n_627) );
INVxp33_ASAP7_75t_L g718 ( .A(n_76), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_76), .A2(n_195), .B1(n_763), .B2(n_765), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g1006 ( .A1(n_77), .A2(n_209), .B1(n_969), .B2(n_1007), .C(n_1009), .Y(n_1006) );
INVx1_ASAP7_75t_L g1048 ( .A(n_77), .Y(n_1048) );
CKINVDCx16_ASAP7_75t_R g1196 ( .A(n_78), .Y(n_1196) );
INVxp33_ASAP7_75t_L g465 ( .A(n_79), .Y(n_465) );
INVx1_ASAP7_75t_L g972 ( .A(n_80), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_81), .A2(n_128), .B1(n_1155), .B2(n_1158), .Y(n_1154) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_82), .A2(n_136), .B1(n_761), .B2(n_805), .C(n_807), .Y(n_804) );
INVxp33_ASAP7_75t_SL g817 ( .A(n_82), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g1397 ( .A1(n_83), .A2(n_1398), .B1(n_1399), .B2(n_1400), .Y(n_1397) );
CKINVDCx5p33_ASAP7_75t_R g1399 ( .A(n_83), .Y(n_1399) );
INVx1_ASAP7_75t_L g339 ( .A(n_84), .Y(n_339) );
INVx1_ASAP7_75t_L g368 ( .A(n_84), .Y(n_368) );
INVxp33_ASAP7_75t_L g431 ( .A(n_85), .Y(n_431) );
INVx1_ASAP7_75t_L g623 ( .A(n_86), .Y(n_623) );
INVx1_ASAP7_75t_L g443 ( .A(n_87), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_87), .A2(n_164), .B1(n_458), .B2(n_460), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_88), .Y(n_635) );
INVx1_ASAP7_75t_L g801 ( .A(n_89), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_90), .A2(n_188), .B1(n_789), .B2(n_791), .Y(n_788) );
INVxp67_ASAP7_75t_L g835 ( .A(n_90), .Y(n_835) );
INVx1_ASAP7_75t_L g313 ( .A(n_91), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_91), .A2(n_375), .B(n_376), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_92), .A2(n_115), .B1(n_584), .B2(n_589), .C(n_854), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_92), .A2(n_115), .B1(n_540), .B2(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g902 ( .A(n_93), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g928 ( .A1(n_93), .A2(n_192), .B1(n_929), .B2(n_931), .C(n_933), .Y(n_928) );
INVxp67_ASAP7_75t_SL g1090 ( .A(n_94), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g1111 ( .A1(n_94), .A2(n_182), .B1(n_491), .B2(n_549), .C(n_761), .Y(n_1111) );
INVxp33_ASAP7_75t_SL g1080 ( .A(n_95), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_95), .A2(n_111), .B1(n_885), .B2(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g636 ( .A(n_96), .Y(n_636) );
OAI221xp5_ASAP7_75t_L g654 ( .A1(n_96), .A2(n_155), .B1(n_655), .B2(n_657), .C(n_658), .Y(n_654) );
INVx1_ASAP7_75t_L g1179 ( .A(n_97), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_98), .A2(n_138), .B1(n_490), .B2(n_492), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_98), .A2(n_138), .B1(n_507), .B2(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g633 ( .A(n_99), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_99), .A2(n_140), .B1(n_298), .B2(n_323), .C(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g797 ( .A(n_100), .Y(n_797) );
OAI221xp5_ASAP7_75t_L g818 ( .A1(n_100), .A2(n_196), .B1(n_584), .B2(n_589), .C(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g916 ( .A(n_101), .Y(n_916) );
AO221x2_ASAP7_75t_L g1132 ( .A1(n_102), .A2(n_165), .B1(n_1133), .B2(n_1139), .C(n_1140), .Y(n_1132) );
INVxp33_ASAP7_75t_L g599 ( .A(n_103), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g1012 ( .A(n_104), .Y(n_1012) );
INVx1_ASAP7_75t_L g538 ( .A(n_105), .Y(n_538) );
OAI22xp33_ASAP7_75t_SL g1036 ( .A1(n_106), .A2(n_184), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
INVx1_ASAP7_75t_L g1062 ( .A(n_106), .Y(n_1062) );
INVx1_ASAP7_75t_L g732 ( .A(n_107), .Y(n_732) );
INVx1_ASAP7_75t_L g1093 ( .A(n_108), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_108), .A2(n_153), .B1(n_535), .B2(n_763), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_109), .A2(n_146), .B1(n_789), .B2(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g992 ( .A(n_109), .Y(n_992) );
INVx1_ASAP7_75t_L g240 ( .A(n_110), .Y(n_240) );
INVxp33_ASAP7_75t_SL g1084 ( .A(n_111), .Y(n_1084) );
INVx1_ASAP7_75t_L g690 ( .A(n_113), .Y(n_690) );
XNOR2x1_ASAP7_75t_L g843 ( .A(n_114), .B(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g1365 ( .A(n_116), .Y(n_1365) );
AOI221xp5_ASAP7_75t_L g1374 ( .A1(n_116), .A2(n_181), .B1(n_1007), .B2(n_1375), .C(n_1376), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_117), .A2(n_141), .B1(n_693), .B2(n_1017), .C(n_1019), .Y(n_1016) );
INVx1_ASAP7_75t_L g1065 ( .A(n_117), .Y(n_1065) );
INVx1_ASAP7_75t_L g865 ( .A(n_118), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_119), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_120), .A2(n_160), .B1(n_1139), .B2(n_1161), .Y(n_1160) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_121), .Y(n_1024) );
INVx1_ASAP7_75t_L g1386 ( .A(n_122), .Y(n_1386) );
INVx1_ASAP7_75t_L g324 ( .A(n_123), .Y(n_324) );
INVx1_ASAP7_75t_L g776 ( .A(n_124), .Y(n_776) );
INVxp67_ASAP7_75t_L g451 ( .A(n_125), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_126), .A2(n_166), .B1(n_540), .B2(n_542), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g583 ( .A1(n_126), .A2(n_166), .B1(n_584), .B2(n_589), .C(n_593), .Y(n_583) );
INVx1_ASAP7_75t_L g1165 ( .A(n_127), .Y(n_1165) );
INVxp33_ASAP7_75t_L g574 ( .A(n_129), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_130), .A2(n_190), .B1(n_315), .B2(n_1372), .Y(n_1371) );
OAI22xp5_ASAP7_75t_L g1388 ( .A1(n_130), .A2(n_206), .B1(n_1034), .B2(n_1389), .Y(n_1388) );
INVxp33_ASAP7_75t_L g1081 ( .A(n_131), .Y(n_1081) );
INVx1_ASAP7_75t_L g872 ( .A(n_132), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_133), .Y(n_269) );
INVx1_ASAP7_75t_L g987 ( .A(n_134), .Y(n_987) );
INVx1_ASAP7_75t_L g674 ( .A(n_135), .Y(n_674) );
INVxp33_ASAP7_75t_SL g815 ( .A(n_136), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_137), .A2(n_152), .B1(n_1155), .B2(n_1158), .Y(n_1168) );
INVx1_ASAP7_75t_L g566 ( .A(n_139), .Y(n_566) );
INVx1_ASAP7_75t_L g640 ( .A(n_140), .Y(n_640) );
INVx1_ASAP7_75t_L g1067 ( .A(n_141), .Y(n_1067) );
OAI221xp5_ASAP7_75t_L g1086 ( .A1(n_142), .A2(n_231), .B1(n_584), .B2(n_590), .C(n_854), .Y(n_1086) );
OAI22xp33_ASAP7_75t_L g1118 ( .A1(n_142), .A2(n_231), .B1(n_754), .B2(n_755), .Y(n_1118) );
INVx1_ASAP7_75t_L g1356 ( .A(n_143), .Y(n_1356) );
INVx1_ASAP7_75t_L g954 ( .A(n_145), .Y(n_954) );
INVx1_ASAP7_75t_L g986 ( .A(n_146), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_147), .Y(n_274) );
XNOR2xp5_ASAP7_75t_L g700 ( .A(n_148), .B(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_148), .A2(n_186), .B1(n_1133), .B2(n_1170), .Y(n_1169) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_149), .Y(n_1029) );
INVx1_ASAP7_75t_L g1075 ( .A(n_150), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_151), .Y(n_242) );
AND3x2_ASAP7_75t_L g1137 ( .A(n_151), .B(n_240), .C(n_1138), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_151), .B(n_240), .Y(n_1144) );
INVxp67_ASAP7_75t_SL g1089 ( .A(n_153), .Y(n_1089) );
INVx1_ASAP7_75t_L g637 ( .A(n_155), .Y(n_637) );
INVx2_ASAP7_75t_L g253 ( .A(n_157), .Y(n_253) );
INVx1_ASAP7_75t_L g905 ( .A(n_158), .Y(n_905) );
INVxp33_ASAP7_75t_L g863 ( .A(n_159), .Y(n_863) );
AOI222xp33_ASAP7_75t_L g1340 ( .A1(n_160), .A2(n_1341), .B1(n_1394), .B2(n_1396), .C1(n_1401), .C2(n_1405), .Y(n_1340) );
XNOR2x2_ASAP7_75t_L g1344 ( .A(n_160), .B(n_1345), .Y(n_1344) );
INVxp67_ASAP7_75t_L g723 ( .A(n_161), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_161), .A2(n_211), .B1(n_549), .B2(n_760), .C(n_761), .Y(n_759) );
INVxp67_ASAP7_75t_L g833 ( .A(n_162), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g1206 ( .A1(n_163), .A2(n_170), .B1(n_1139), .B2(n_1161), .Y(n_1206) );
INVx1_ASAP7_75t_L g438 ( .A(n_164), .Y(n_438) );
INVx1_ASAP7_75t_L g867 ( .A(n_167), .Y(n_867) );
INVx1_ASAP7_75t_L g1138 ( .A(n_168), .Y(n_1138) );
AOI221xp5_ASAP7_75t_L g545 ( .A1(n_169), .A2(n_225), .B1(n_534), .B2(n_546), .C(n_549), .Y(n_545) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_169), .Y(n_607) );
INVx1_ASAP7_75t_L g1362 ( .A(n_171), .Y(n_1362) );
CKINVDCx16_ASAP7_75t_R g1176 ( .A(n_172), .Y(n_1176) );
INVx1_ASAP7_75t_L g1249 ( .A(n_173), .Y(n_1249) );
INVx1_ASAP7_75t_L g1350 ( .A(n_174), .Y(n_1350) );
INVx1_ASAP7_75t_L g1060 ( .A(n_175), .Y(n_1060) );
INVx1_ASAP7_75t_L g334 ( .A(n_176), .Y(n_334) );
OAI211xp5_ASAP7_75t_L g386 ( .A1(n_176), .A2(n_387), .B(n_389), .C(n_397), .Y(n_386) );
INVx1_ASAP7_75t_L g1099 ( .A(n_177), .Y(n_1099) );
CKINVDCx5p33_ASAP7_75t_R g1043 ( .A(n_178), .Y(n_1043) );
INVx1_ASAP7_75t_L g255 ( .A(n_179), .Y(n_255) );
INVx2_ASAP7_75t_L g310 ( .A(n_179), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_180), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_181), .A2(n_185), .B1(n_925), .B2(n_1367), .Y(n_1366) );
INVxp67_ASAP7_75t_SL g1092 ( .A(n_182), .Y(n_1092) );
AOI22xp5_ASAP7_75t_L g1205 ( .A1(n_183), .A2(n_204), .B1(n_1155), .B2(n_1158), .Y(n_1205) );
INVx1_ASAP7_75t_L g1056 ( .A(n_184), .Y(n_1056) );
INVx1_ASAP7_75t_L g1377 ( .A(n_185), .Y(n_1377) );
INVx1_ASAP7_75t_L g347 ( .A(n_187), .Y(n_347) );
INVxp67_ASAP7_75t_L g824 ( .A(n_188), .Y(n_824) );
INVxp33_ASAP7_75t_L g851 ( .A(n_189), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g877 ( .A1(n_189), .A2(n_191), .B1(n_391), .B2(n_531), .C(n_746), .Y(n_877) );
OAI22xp33_ASAP7_75t_L g1390 ( .A1(n_190), .A2(n_212), .B1(n_787), .B2(n_1020), .Y(n_1390) );
INVxp33_ASAP7_75t_L g849 ( .A(n_191), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_193), .A2(n_205), .B1(n_533), .B2(n_554), .Y(n_910) );
OAI221xp5_ASAP7_75t_L g919 ( .A1(n_193), .A2(n_205), .B1(n_728), .B2(n_920), .C(n_921), .Y(n_919) );
INVx1_ASAP7_75t_L g1097 ( .A(n_194), .Y(n_1097) );
INVxp67_ASAP7_75t_L g727 ( .A(n_195), .Y(n_727) );
INVx1_ASAP7_75t_L g798 ( .A(n_196), .Y(n_798) );
INVx1_ASAP7_75t_L g1190 ( .A(n_198), .Y(n_1190) );
INVx1_ASAP7_75t_L g871 ( .A(n_199), .Y(n_871) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_200), .A2(n_233), .B1(n_391), .B2(n_529), .C(n_531), .Y(n_528) );
INVxp33_ASAP7_75t_L g580 ( .A(n_200), .Y(n_580) );
INVx1_ASAP7_75t_L g1136 ( .A(n_201), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_201), .B(n_1146), .Y(n_1149) );
AOI21xp33_ASAP7_75t_L g957 ( .A1(n_202), .A2(n_531), .B(n_790), .Y(n_957) );
INVxp33_ASAP7_75t_L g979 ( .A(n_202), .Y(n_979) );
INVxp33_ASAP7_75t_L g980 ( .A(n_203), .Y(n_980) );
INVxp67_ASAP7_75t_SL g1370 ( .A(n_206), .Y(n_1370) );
INVx1_ASAP7_75t_L g795 ( .A(n_207), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_208), .Y(n_874) );
INVx1_ASAP7_75t_L g1053 ( .A(n_209), .Y(n_1053) );
INVx1_ASAP7_75t_L g768 ( .A(n_210), .Y(n_768) );
INVxp33_ASAP7_75t_L g719 ( .A(n_211), .Y(n_719) );
INVxp67_ASAP7_75t_SL g1369 ( .A(n_212), .Y(n_1369) );
INVx1_ASAP7_75t_L g639 ( .A(n_213), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_213), .A2(n_286), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g738 ( .A(n_214), .Y(n_738) );
INVx2_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_216), .Y(n_632) );
INVx1_ASAP7_75t_L g794 ( .A(n_217), .Y(n_794) );
XNOR2x2_ASAP7_75t_L g1003 ( .A(n_218), .B(n_1004), .Y(n_1003) );
INVxp33_ASAP7_75t_L g705 ( .A(n_219), .Y(n_705) );
INVxp33_ASAP7_75t_SL g1352 ( .A(n_221), .Y(n_1352) );
OAI22x1_ASAP7_75t_SL g410 ( .A1(n_222), .A2(n_411), .B1(n_518), .B2(n_519), .Y(n_410) );
INVx1_ASAP7_75t_L g518 ( .A(n_222), .Y(n_518) );
INVx1_ASAP7_75t_L g971 ( .A(n_223), .Y(n_971) );
INVx1_ASAP7_75t_L g1354 ( .A(n_224), .Y(n_1354) );
INVxp33_ASAP7_75t_SL g602 ( .A(n_225), .Y(n_602) );
INVx1_ASAP7_75t_L g1101 ( .A(n_226), .Y(n_1101) );
INVx1_ASAP7_75t_L g342 ( .A(n_227), .Y(n_342) );
BUFx3_ASAP7_75t_L g356 ( .A(n_227), .Y(n_356) );
INVx1_ASAP7_75t_L g344 ( .A(n_228), .Y(n_344) );
BUFx3_ASAP7_75t_L g358 ( .A(n_228), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g1013 ( .A(n_229), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_230), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_232), .Y(n_327) );
INVxp33_ASAP7_75t_L g578 ( .A(n_233), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_256), .B(n_1124), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_243), .Y(n_237) );
AND2x4_ASAP7_75t_L g1395 ( .A(n_238), .B(n_244), .Y(n_1395) );
NOR2xp33_ASAP7_75t_SL g238 ( .A(n_239), .B(n_241), .Y(n_238) );
INVx1_ASAP7_75t_SL g1404 ( .A(n_239), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_239), .B(n_241), .Y(n_1410) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_241), .B(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g475 ( .A(n_246), .B(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g284 ( .A(n_247), .B(n_255), .Y(n_284) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g597 ( .A(n_248), .B(n_464), .Y(n_597) );
INVx8_ASAP7_75t_L g471 ( .A(n_249), .Y(n_471) );
OR2x6_ASAP7_75t_L g249 ( .A(n_250), .B(n_254), .Y(n_249) );
OR2x2_ASAP7_75t_L g333 ( .A(n_250), .B(n_267), .Y(n_333) );
OR2x6_ASAP7_75t_L g474 ( .A(n_250), .B(n_463), .Y(n_474) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_250), .Y(n_601) );
INVx1_ASAP7_75t_L g823 ( .A(n_250), .Y(n_823) );
INVx2_ASAP7_75t_SL g840 ( .A(n_250), .Y(n_840) );
INVx2_ASAP7_75t_SL g870 ( .A(n_250), .Y(n_870) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g273 ( .A(n_252), .Y(n_273) );
INVx1_ASAP7_75t_L g278 ( .A(n_252), .Y(n_278) );
AND2x2_ASAP7_75t_L g289 ( .A(n_252), .B(n_253), .Y(n_289) );
INVx2_ASAP7_75t_L g295 ( .A(n_252), .Y(n_295) );
AND2x4_ASAP7_75t_L g301 ( .A(n_252), .B(n_279), .Y(n_301) );
INVx1_ASAP7_75t_L g265 ( .A(n_253), .Y(n_265) );
INVx2_ASAP7_75t_L g279 ( .A(n_253), .Y(n_279) );
INVx1_ASAP7_75t_L g297 ( .A(n_253), .Y(n_297) );
INVx1_ASAP7_75t_L g605 ( .A(n_253), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_253), .B(n_295), .Y(n_612) );
AND2x4_ASAP7_75t_L g459 ( .A(n_254), .B(n_265), .Y(n_459) );
INVx2_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g460 ( .A(n_255), .B(n_272), .Y(n_460) );
XNOR2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_771), .Y(n_256) );
XNOR2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_407), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND3xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_320), .C(n_335), .Y(n_260) );
AND3x1_ASAP7_75t_L g261 ( .A(n_262), .B(n_280), .C(n_312), .Y(n_261) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_269), .B1(n_270), .B2(n_274), .C(n_275), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_263), .A2(n_270), .B1(n_275), .B2(n_904), .C(n_905), .Y(n_944) );
INVx1_ASAP7_75t_L g1072 ( .A(n_263), .Y(n_1072) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g588 ( .A(n_265), .Y(n_588) );
AND2x4_ASAP7_75t_L g270 ( .A(n_266), .B(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g275 ( .A(n_266), .B(n_276), .Y(n_275) );
NAND2x1_ASAP7_75t_SL g586 ( .A(n_266), .B(n_587), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_266), .B(n_591), .Y(n_590) );
NAND2x1p5_ASAP7_75t_L g594 ( .A(n_266), .B(n_326), .Y(n_594) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g647 ( .A(n_268), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_269), .A2(n_274), .B1(n_398), .B2(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g1070 ( .A(n_270), .Y(n_1070) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g604 ( .A(n_273), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_273), .B(n_605), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_275), .A2(n_1042), .B1(n_1043), .B2(n_1069), .C(n_1071), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1393 ( .A1(n_275), .A2(n_1069), .B1(n_1071), .B2(n_1385), .C(n_1386), .Y(n_1393) );
INVx1_ASAP7_75t_L g453 ( .A(n_276), .Y(n_453) );
BUFx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g291 ( .A(n_277), .Y(n_291) );
BUFx3_ASAP7_75t_L g326 ( .A(n_277), .Y(n_326) );
AND2x4_ASAP7_75t_L g454 ( .A(n_277), .B(n_455), .Y(n_454) );
BUFx3_ASAP7_75t_L g670 ( .A(n_277), .Y(n_670) );
BUFx6f_ASAP7_75t_L g927 ( .A(n_277), .Y(n_927) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI33xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_285), .A3(n_292), .B1(n_302), .B2(n_305), .B3(n_306), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_281), .A2(n_332), .B1(n_916), .B2(n_936), .Y(n_935) );
AND2x4_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
AND2x2_ASAP7_75t_L g306 ( .A(n_282), .B(n_307), .Y(n_306) );
OR2x6_ASAP7_75t_L g480 ( .A(n_282), .B(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g503 ( .A(n_282), .B(n_284), .Y(n_503) );
INVx2_ASAP7_75t_L g781 ( .A(n_282), .Y(n_781) );
BUFx2_ASAP7_75t_L g1392 ( .A(n_282), .Y(n_1392) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g406 ( .A(n_283), .Y(n_406) );
OR2x6_ASAP7_75t_L g596 ( .A(n_283), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g1367 ( .A(n_287), .Y(n_1367) );
INVx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g505 ( .A(n_288), .Y(n_505) );
AND2x4_ASAP7_75t_L g672 ( .A(n_288), .B(n_319), .Y(n_672) );
BUFx6f_ASAP7_75t_L g923 ( .A(n_288), .Y(n_923) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_294), .Y(n_303) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
AND2x4_ASAP7_75t_L g462 ( .A(n_294), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g675 ( .A(n_294), .B(n_319), .Y(n_675) );
INVx1_ASAP7_75t_L g930 ( .A(n_294), .Y(n_930) );
INVx1_ASAP7_75t_L g938 ( .A(n_294), .Y(n_938) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g592 ( .A(n_295), .Y(n_592) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx3_ASAP7_75t_L g513 ( .A(n_299), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_299), .A2(n_1013), .B1(n_1051), .B2(n_1053), .Y(n_1050) );
INVx2_ASAP7_75t_L g1364 ( .A(n_299), .Y(n_1364) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g330 ( .A(n_300), .Y(n_330) );
INVx3_ASAP7_75t_L g577 ( .A(n_300), .Y(n_577) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_301), .Y(n_304) );
INVx1_ASAP7_75t_L g468 ( .A(n_301), .Y(n_468) );
INVx1_ASAP7_75t_L g679 ( .A(n_301), .Y(n_679) );
BUFx3_ASAP7_75t_L g507 ( .A(n_303), .Y(n_507) );
INVx2_ASAP7_75t_SL g614 ( .A(n_304), .Y(n_614) );
INVx2_ASAP7_75t_SL g728 ( .A(n_304), .Y(n_728) );
INVx4_ASAP7_75t_L g860 ( .A(n_304), .Y(n_860) );
INVx2_ASAP7_75t_SL g940 ( .A(n_304), .Y(n_940) );
BUFx3_ASAP7_75t_L g991 ( .A(n_304), .Y(n_991) );
INVx2_ASAP7_75t_SL g653 ( .A(n_307), .Y(n_653) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x6_ASAP7_75t_L g516 ( .A(n_308), .B(n_517), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g456 ( .A(n_309), .Y(n_456) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g464 ( .A(n_310), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_314), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_314), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_314), .A2(n_582), .B1(n_801), .B2(n_817), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_314), .A2(n_711), .B1(n_851), .B2(n_852), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_314), .A2(n_582), .B1(n_979), .B2(n_980), .Y(n_978) );
BUFx2_ASAP7_75t_L g1045 ( .A(n_314), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_314), .A2(n_1083), .B1(n_1084), .B2(n_1085), .Y(n_1082) );
AOI21xp5_ASAP7_75t_L g1355 ( .A1(n_314), .A2(n_1356), .B(n_1357), .Y(n_1355) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_SL g665 ( .A(n_316), .Y(n_665) );
AND2x2_ASAP7_75t_L g322 ( .A(n_317), .B(n_323), .Y(n_322) );
AND2x6_ASAP7_75t_L g325 ( .A(n_317), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g329 ( .A(n_317), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g576 ( .A(n_317), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g582 ( .A(n_317), .B(n_323), .Y(n_582) );
AND2x2_ASAP7_75t_L g711 ( .A(n_317), .B(n_323), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_317), .A2(n_515), .B1(n_919), .B2(n_928), .Y(n_918) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_317), .B(n_323), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_317), .B(n_323), .Y(n_1353) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g517 ( .A(n_318), .Y(n_517) );
INVx2_ASAP7_75t_L g669 ( .A(n_319), .Y(n_669) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_328), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B1(n_325), .B2(n_327), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_325), .A2(n_574), .B1(n_575), .B2(n_578), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_325), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_325), .A2(n_803), .B1(n_814), .B2(n_815), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_325), .A2(n_576), .B1(n_848), .B2(n_849), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_325), .A2(n_706), .B1(n_954), .B2(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_325), .A2(n_576), .B1(n_1021), .B2(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_325), .A2(n_575), .B1(n_1080), .B2(n_1081), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_325), .A2(n_1348), .B1(n_1349), .B2(n_1350), .Y(n_1347) );
OAI211xp5_ASAP7_75t_L g370 ( .A1(n_327), .A2(n_371), .B(n_373), .C(n_374), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B1(n_332), .B2(n_334), .Y(n_328) );
INVx2_ASAP7_75t_L g734 ( .A(n_330), .Y(n_734) );
INVx2_ASAP7_75t_L g866 ( .A(n_330), .Y(n_866) );
INVx1_ASAP7_75t_L g932 ( .A(n_330), .Y(n_932) );
AOI22xp33_ASAP7_75t_SL g1066 ( .A1(n_332), .A2(n_582), .B1(n_1029), .B2(n_1067), .Y(n_1066) );
AOI22xp33_ASAP7_75t_SL g1351 ( .A1(n_332), .A2(n_1352), .B1(n_1353), .B2(n_1354), .Y(n_1351) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g568 ( .A(n_333), .B(n_569), .Y(n_568) );
OAI31xp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_345), .A3(n_386), .B(n_405), .Y(n_335) );
INVx6_ASAP7_75t_L g562 ( .A(n_337), .Y(n_562) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx2_ASAP7_75t_L g396 ( .A(n_338), .Y(n_396) );
OR2x2_ASAP7_75t_L g565 ( .A(n_338), .B(n_361), .Y(n_565) );
INVx1_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
INVx2_ASAP7_75t_L g686 ( .A(n_340), .Y(n_686) );
INVx1_ASAP7_75t_L g1023 ( .A(n_340), .Y(n_1023) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
AND2x2_ASAP7_75t_L g350 ( .A(n_341), .B(n_343), .Y(n_350) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g362 ( .A(n_342), .B(n_358), .Y(n_362) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g365 ( .A(n_344), .B(n_356), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_370), .C(n_379), .Y(n_345) );
OAI211xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B(n_351), .C(n_363), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g955 ( .A(n_349), .Y(n_955) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_349), .Y(n_1020) );
BUFx4f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_350), .Y(n_1011) );
INVx1_ASAP7_75t_L g764 ( .A(n_352), .Y(n_764) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g375 ( .A(n_353), .Y(n_375) );
INVx2_ASAP7_75t_L g421 ( .A(n_353), .Y(n_421) );
INVx1_ASAP7_75t_L g484 ( .A(n_353), .Y(n_484) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_353), .Y(n_530) );
INVx2_ASAP7_75t_L g747 ( .A(n_353), .Y(n_747) );
INVx2_ASAP7_75t_L g790 ( .A(n_353), .Y(n_790) );
INVx6_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g388 ( .A(n_354), .B(n_382), .Y(n_388) );
AND2x4_ASAP7_75t_L g428 ( .A(n_354), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g553 ( .A(n_354), .Y(n_553) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_354), .Y(n_1115) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g404 ( .A(n_355), .Y(n_404) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g385 ( .A(n_356), .B(n_358), .Y(n_385) );
INVx1_ASAP7_75t_L g401 ( .A(n_357), .Y(n_401) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g900 ( .A(n_359), .Y(n_900) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g395 ( .A(n_360), .Y(n_395) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g1117 ( .A(n_361), .Y(n_1117) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_362), .Y(n_433) );
INVx1_ASAP7_75t_L g493 ( .A(n_362), .Y(n_493) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_362), .Y(n_536) );
BUFx3_ASAP7_75t_L g692 ( .A(n_364), .Y(n_692) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_365), .Y(n_394) );
AND2x6_ASAP7_75t_L g423 ( .A(n_365), .B(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_365), .Y(n_491) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_365), .Y(n_496) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_365), .Y(n_534) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_365), .Y(n_752) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_365), .Y(n_760) );
BUFx2_ASAP7_75t_L g885 ( .A(n_365), .Y(n_885) );
INVx2_ASAP7_75t_SL g1018 ( .A(n_365), .Y(n_1018) );
INVx1_ASAP7_75t_L g967 ( .A(n_366), .Y(n_967) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g481 ( .A(n_367), .Y(n_481) );
BUFx3_ASAP7_75t_L g550 ( .A(n_367), .Y(n_550) );
INVx1_ASAP7_75t_L g1015 ( .A(n_367), .Y(n_1015) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
AND2x4_ASAP7_75t_L g377 ( .A(n_368), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g413 ( .A(n_368), .Y(n_413) );
INVx2_ASAP7_75t_L g378 ( .A(n_369), .Y(n_378) );
INVx1_ASAP7_75t_L g420 ( .A(n_369), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_369), .Y(n_425) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_369), .Y(n_430) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g689 ( .A(n_372), .Y(n_689) );
INVx1_ASAP7_75t_L g1008 ( .A(n_375), .Y(n_1008) );
INVx1_ASAP7_75t_L g1025 ( .A(n_376), .Y(n_1025) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g500 ( .A(n_377), .B(n_476), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_377), .Y(n_531) );
INVx1_ASAP7_75t_L g748 ( .A(n_377), .Y(n_748) );
INVx2_ASAP7_75t_L g807 ( .A(n_377), .Y(n_807) );
HB1xp67_ASAP7_75t_L g1381 ( .A(n_377), .Y(n_1381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_378), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .Y(n_380) );
BUFx3_ASAP7_75t_L g1031 ( .A(n_381), .Y(n_1031) );
BUFx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g398 ( .A(n_382), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g402 ( .A(n_382), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g541 ( .A(n_382), .B(n_399), .Y(n_541) );
AND2x2_ASAP7_75t_L g543 ( .A(n_382), .B(n_403), .Y(n_543) );
INVx1_ASAP7_75t_L g559 ( .A(n_382), .Y(n_559) );
BUFx4f_ASAP7_75t_L g391 ( .A(n_384), .Y(n_391) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
AND2x4_ASAP7_75t_L g555 ( .A(n_384), .B(n_396), .Y(n_555) );
INVx1_ASAP7_75t_L g745 ( .A(n_384), .Y(n_745) );
BUFx3_ASAP7_75t_L g761 ( .A(n_384), .Y(n_761) );
INVx2_ASAP7_75t_SL g909 ( .A(n_384), .Y(n_909) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_385), .Y(n_448) );
INVx2_ASAP7_75t_L g915 ( .A(n_387), .Y(n_915) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g570 ( .A(n_388), .B(n_476), .Y(n_570) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_392), .C(n_396), .Y(n_389) );
INVx1_ASAP7_75t_L g1379 ( .A(n_393), .Y(n_1379) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g787 ( .A(n_394), .Y(n_787) );
INVx1_ASAP7_75t_L g699 ( .A(n_395), .Y(n_699) );
AND2x4_ASAP7_75t_L g537 ( .A(n_396), .B(n_534), .Y(n_537) );
AOI222xp33_ASAP7_75t_L g897 ( .A1(n_396), .A2(n_541), .B1(n_543), .B2(n_898), .C1(n_904), .C2(n_905), .Y(n_897) );
OAI21xp33_ASAP7_75t_L g1032 ( .A1(n_396), .A2(n_1033), .B(n_1036), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_396), .B(n_491), .Y(n_1107) );
OAI21xp5_ASAP7_75t_L g1387 ( .A1(n_396), .A2(n_1388), .B(n_1390), .Y(n_1387) );
INVx2_ASAP7_75t_L g754 ( .A(n_398), .Y(n_754) );
INVx4_ASAP7_75t_L g1041 ( .A(n_398), .Y(n_1041) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g442 ( .A(n_401), .Y(n_442) );
INVx2_ASAP7_75t_L g755 ( .A(n_402), .Y(n_755) );
INVx2_ASAP7_75t_SL g882 ( .A(n_402), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_402), .A2(n_1040), .B1(n_1042), .B2(n_1043), .Y(n_1039) );
BUFx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x6_ASAP7_75t_L g444 ( .A(n_404), .B(n_425), .Y(n_444) );
INVx2_ASAP7_75t_L g973 ( .A(n_405), .Y(n_973) );
OAI31xp33_ASAP7_75t_SL g1005 ( .A1(n_405), .A2(n_1006), .A3(n_1016), .B(n_1026), .Y(n_1005) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g412 ( .A(n_406), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g525 ( .A(n_406), .Y(n_525) );
XOR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_625), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_520), .B2(n_624), .Y(n_408) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g519 ( .A(n_411), .Y(n_519) );
AO211x2_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B(n_449), .C(n_477), .Y(n_411) );
AOI221x1_ASAP7_75t_SL g628 ( .A1(n_412), .A2(n_629), .B1(n_641), .B2(n_680), .C(n_681), .Y(n_628) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_415), .B(n_426), .C(n_434), .D(n_445), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B1(n_422), .B2(n_423), .Y(n_415) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_418), .A2(n_423), .B1(n_639), .B2(n_640), .Y(n_638) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
AND2x6_ASAP7_75t_L g432 ( .A(n_419), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g447 ( .A(n_424), .Y(n_447) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_431), .B2(n_432), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_427), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_428), .A2(n_432), .B1(n_632), .B2(n_633), .Y(n_631) );
AND2x4_ASAP7_75t_L g440 ( .A(n_429), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g498 ( .A(n_433), .Y(n_498) );
INVx2_ASAP7_75t_L g766 ( .A(n_433), .Y(n_766) );
BUFx6f_ASAP7_75t_L g969 ( .A(n_433), .Y(n_969) );
BUFx6f_ASAP7_75t_L g1375 ( .A(n_433), .Y(n_1375) );
AOI222xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_438), .B2(n_439), .C1(n_443), .C2(n_444), .Y(n_434) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_439), .A2(n_444), .B1(n_485), .B2(n_635), .C1(n_636), .C2(n_637), .Y(n_634) );
BUFx4f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g630 ( .A(n_445), .Y(n_630) );
INVx5_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx2_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_448), .Y(n_548) );
INVx1_ASAP7_75t_L g965 ( .A(n_448), .Y(n_965) );
AOI31xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_461), .A3(n_470), .B(n_475), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_454), .C(n_457), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_465), .B1(n_466), .B2(n_469), .Y(n_461) );
AND2x4_ASAP7_75t_L g466 ( .A(n_463), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_468), .Y(n_511) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_501), .Y(n_477) );
AOI33xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_482), .A3(n_489), .B1(n_494), .B2(n_495), .B3(n_499), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g683 ( .A(n_480), .Y(n_683) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g901 ( .A1(n_491), .A2(n_548), .B1(n_902), .B2(n_903), .Y(n_901) );
INVx1_ASAP7_75t_L g962 ( .A(n_491), .Y(n_962) );
INVx1_ASAP7_75t_L g1037 ( .A(n_491), .Y(n_1037) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g554 ( .A(n_493), .Y(n_554) );
INVx1_ASAP7_75t_L g914 ( .A(n_493), .Y(n_914) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx4f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx4_ASAP7_75t_L g694 ( .A(n_500), .Y(n_694) );
AOI33xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_504), .A3(n_506), .B1(n_512), .B2(n_514), .B3(n_515), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g834 ( .A(n_513), .Y(n_834) );
INVx1_ASAP7_75t_L g1057 ( .A(n_513), .Y(n_1057) );
INVx2_ASAP7_75t_L g842 ( .A(n_515), .Y(n_842) );
INVx6_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx5_ASAP7_75t_L g622 ( .A(n_516), .Y(n_622) );
BUFx2_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g624 ( .A(n_521), .Y(n_624) );
XOR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_623), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_571), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_526), .B1(n_566), .B2(n_567), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx8_ASAP7_75t_SL g680 ( .A(n_525), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_544), .C(n_560), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_532), .B1(n_537), .B2(n_538), .C(n_539), .Y(n_527) );
INVx4_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g1028 ( .A(n_530), .Y(n_1028) );
INVxp67_ASAP7_75t_L g800 ( .A(n_533), .Y(n_800) );
BUFx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g880 ( .A(n_534), .Y(n_880) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g693 ( .A(n_536), .Y(n_693) );
INVx1_ASAP7_75t_L g792 ( .A(n_536), .Y(n_792) );
INVx1_ASAP7_75t_L g1035 ( .A(n_536), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_537), .A2(n_562), .B1(n_732), .B2(n_737), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_537), .B(n_809), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_537), .A2(n_865), .B1(n_877), .B2(n_878), .C(n_881), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_537), .A2(n_951), .B(n_952), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_538), .A2(n_563), .B1(n_608), .B2(n_616), .Y(n_615) );
INVx2_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_541), .A2(n_543), .B1(n_797), .B2(n_798), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_541), .A2(n_543), .B1(n_1385), .B2(n_1386), .Y(n_1384) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_551), .B1(n_555), .B2(n_556), .C(n_557), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g1030 ( .A(n_547), .Y(n_1030) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g557 ( .A(n_548), .B(n_558), .Y(n_557) );
BUFx6f_ASAP7_75t_L g886 ( .A(n_548), .Y(n_886) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g802 ( .A(n_554), .Y(n_802) );
INVx1_ASAP7_75t_L g758 ( .A(n_555), .Y(n_758) );
BUFx6f_ASAP7_75t_L g888 ( .A(n_555), .Y(n_888) );
INVx2_ASAP7_75t_SL g1110 ( .A(n_555), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_556), .A2(n_561), .B1(n_600), .B2(n_619), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_557), .A2(n_738), .B1(n_757), .B2(n_759), .C(n_762), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_557), .A2(n_757), .B1(n_784), .B2(n_785), .C(n_788), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_557), .A2(n_872), .B1(n_884), .B2(n_887), .C(n_888), .Y(n_883) );
AOI21xp33_ASAP7_75t_L g906 ( .A1(n_557), .A2(n_907), .B(n_910), .Y(n_906) );
AOI221xp5_ASAP7_75t_L g958 ( .A1(n_557), .A2(n_888), .B1(n_959), .B2(n_960), .C(n_968), .Y(n_958) );
AOI221xp5_ASAP7_75t_L g1108 ( .A1(n_557), .A2(n_1101), .B1(n_1109), .B2(n_1111), .C(n_1112), .Y(n_1108) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B1(n_563), .B2(n_564), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_562), .A2(n_564), .B1(n_794), .B2(n_795), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_562), .A2(n_564), .B1(n_867), .B2(n_871), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_562), .A2(n_564), .B1(n_971), .B2(n_972), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g1104 ( .A1(n_562), .A2(n_1096), .B1(n_1099), .B2(n_1105), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g742 ( .A1(n_564), .A2(n_735), .B1(n_743), .B2(n_749), .C(n_753), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g1113 ( .A1(n_564), .A2(n_1097), .B1(n_1114), .B2(n_1116), .C(n_1118), .Y(n_1113) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_567), .A2(n_779), .B1(n_782), .B2(n_810), .Y(n_778) );
AOI21xp33_ASAP7_75t_SL g873 ( .A1(n_567), .A2(n_874), .B(n_875), .Y(n_873) );
AOI21xp33_ASAP7_75t_SL g947 ( .A1(n_567), .A2(n_948), .B(n_949), .Y(n_947) );
INVx5_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g769 ( .A(n_568), .Y(n_769) );
INVx1_ASAP7_75t_L g1120 ( .A(n_568), .Y(n_1120) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NOR3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_583), .C(n_595), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_579), .Y(n_572) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g706 ( .A(n_576), .Y(n_706) );
BUFx2_ASAP7_75t_L g814 ( .A(n_576), .Y(n_814) );
BUFx2_ASAP7_75t_L g1349 ( .A(n_576), .Y(n_1349) );
BUFx3_ASAP7_75t_L g617 ( .A(n_577), .Y(n_617) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g982 ( .A(n_585), .Y(n_982) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2x1p5_ASAP7_75t_L g655 ( .A(n_587), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx4f_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x6_ASAP7_75t_L g657 ( .A(n_592), .B(n_646), .Y(n_657) );
BUFx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g819 ( .A(n_594), .Y(n_819) );
BUFx2_ASAP7_75t_L g854 ( .A(n_594), .Y(n_854) );
OAI33xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .A3(n_606), .B1(n_615), .B2(n_618), .B3(n_621), .Y(n_595) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_596), .Y(n_714) );
OAI33xp33_ASAP7_75t_L g820 ( .A1(n_596), .A2(n_821), .A3(n_830), .B1(n_836), .B2(n_837), .B3(n_842), .Y(n_820) );
OAI33xp33_ASAP7_75t_L g855 ( .A1(n_596), .A2(n_621), .A3(n_856), .B1(n_861), .B2(n_864), .B3(n_868), .Y(n_855) );
OAI33xp33_ASAP7_75t_L g983 ( .A1(n_596), .A2(n_621), .A3(n_984), .B1(n_988), .B2(n_993), .B3(n_994), .Y(n_983) );
OAI33xp33_ASAP7_75t_L g1046 ( .A1(n_596), .A2(n_842), .A3(n_1047), .B1(n_1050), .B2(n_1054), .B3(n_1059), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_596), .A2(n_621), .B1(n_1358), .B2(n_1368), .Y(n_1357) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B1(n_602), .B2(n_603), .Y(n_598) );
BUFx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g717 ( .A(n_601), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g933 ( .A1(n_601), .A2(n_721), .B1(n_903), .B2(n_934), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_601), .A2(n_721), .B1(n_942), .B2(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g996 ( .A(n_601), .Y(n_996) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g620 ( .A(n_604), .Y(n_620) );
INVx2_ASAP7_75t_L g645 ( .A(n_604), .Y(n_645) );
INVx3_ASAP7_75t_L g721 ( .A(n_604), .Y(n_721) );
OAI22xp5_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_608), .B1(n_613), .B2(n_614), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g858 ( .A(n_609), .Y(n_858) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g1095 ( .A(n_610), .Y(n_1095) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx3_ASAP7_75t_L g731 ( .A(n_611), .Y(n_731) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g726 ( .A(n_612), .Y(n_726) );
BUFx2_ASAP7_75t_L g1361 ( .A(n_612), .Y(n_1361) );
OAI221xp5_ASAP7_75t_L g1368 ( .A1(n_614), .A2(n_1055), .B1(n_1369), .B2(n_1370), .C(n_1371), .Y(n_1368) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_617), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_619), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_984) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI33xp33_ASAP7_75t_L g713 ( .A1(n_621), .A2(n_714), .A3(n_715), .B1(n_722), .B2(n_729), .B3(n_736), .Y(n_713) );
OAI33xp33_ASAP7_75t_L g1087 ( .A1(n_621), .A2(n_714), .A3(n_1088), .B1(n_1091), .B2(n_1094), .B3(n_1098), .Y(n_1087) );
CKINVDCx8_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
AO22x2_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_700), .B2(n_770), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .C(n_634), .D(n_638), .Y(n_629) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_632), .A2(n_662), .B1(n_666), .B2(n_667), .C1(n_671), .C2(n_672), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g649 ( .A1(n_635), .A2(n_650), .B(n_652), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_661), .C(n_673), .Y(n_641) );
NOR3xp33_ASAP7_75t_SL g642 ( .A(n_643), .B(n_648), .C(n_654), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OR2x6_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g651 ( .A(n_645), .Y(n_651) );
INVx1_ASAP7_75t_L g656 ( .A(n_646), .Y(n_656) );
INVx1_ASAP7_75t_L g664 ( .A(n_646), .Y(n_664) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g1049 ( .A(n_651), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_666), .A2(n_671), .B1(n_688), .B2(n_696), .C(n_698), .Y(n_695) );
AND2x4_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
AND2x4_ASAP7_75t_L g677 ( .A(n_668), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx6f_ASAP7_75t_L g1372 ( .A(n_670), .Y(n_1372) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_673) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx5_ASAP7_75t_L g740 ( .A(n_680), .Y(n_740) );
AOI31xp33_ASAP7_75t_L g875 ( .A1(n_680), .A2(n_876), .A3(n_883), .B(n_889), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_694), .B2(n_695), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B1(n_688), .B2(n_690), .C(n_691), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_686), .Y(n_697) );
INVx2_ASAP7_75t_L g899 ( .A(n_686), .Y(n_899) );
INVx2_ASAP7_75t_L g1034 ( .A(n_686), .Y(n_1034) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g770 ( .A(n_700), .Y(n_770) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_739), .Y(n_701) );
NOR3xp33_ASAP7_75t_SL g702 ( .A(n_703), .B(n_712), .C(n_713), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_708), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_716), .A2(n_720), .B1(n_737), .B2(n_738), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_716), .A2(n_720), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_716), .A2(n_1099), .B1(n_1100), .B2(n_1101), .Y(n_1098) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_720), .A2(n_869), .B1(n_871), .B2(n_872), .Y(n_868) );
OAI22xp33_ASAP7_75t_L g994 ( .A1(n_720), .A2(n_959), .B1(n_971), .B2(n_995), .Y(n_994) );
BUFx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_727), .B2(n_728), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_724), .A2(n_860), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
BUFx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_725), .A2(n_989), .B1(n_990), .B2(n_992), .Y(n_988) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g1052 ( .A(n_726), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_732), .B1(n_733), .B2(n_735), .Y(n_729) );
INVx2_ASAP7_75t_L g832 ( .A(n_730), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_730), .A2(n_733), .B1(n_951), .B2(n_972), .Y(n_993) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g920 ( .A(n_731), .Y(n_920) );
INVx2_ASAP7_75t_SL g1055 ( .A(n_731), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_768), .B2(n_769), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g1102 ( .A1(n_740), .A2(n_1103), .B1(n_1119), .B2(n_1120), .Y(n_1102) );
NAND3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_756), .C(n_767), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g806 ( .A(n_747), .Y(n_806) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI221xp5_ASAP7_75t_L g1009 ( .A1(n_751), .A2(n_1010), .B1(n_1012), .B2(n_1013), .C(n_1014), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g1376 ( .A1(n_751), .A2(n_967), .B1(n_1038), .B2(n_1362), .C(n_1377), .Y(n_1376) );
INVx2_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_1001), .B2(n_1123), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AO22x1_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_890), .B1(n_999), .B2(n_1000), .Y(n_773) );
INVx1_ASAP7_75t_L g1000 ( .A(n_774), .Y(n_1000) );
XOR2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_843), .Y(n_774) );
XNOR2x1_ASAP7_75t_L g775 ( .A(n_776), .B(n_777), .Y(n_775) );
AND2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_811), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AOI31xp33_ASAP7_75t_SL g896 ( .A1(n_780), .A2(n_897), .A3(n_906), .B(n_911), .Y(n_896) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND5xp2_ASAP7_75t_SL g782 ( .A(n_783), .B(n_793), .C(n_796), .D(n_799), .E(n_808), .Y(n_782) );
OAI22xp33_ASAP7_75t_L g837 ( .A1(n_784), .A2(n_794), .B1(n_838), .B2(n_841), .Y(n_837) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
BUFx3_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_795), .A2(n_809), .B1(n_831), .B2(n_834), .Y(n_836) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B1(n_802), .B2(n_803), .C(n_804), .Y(n_799) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NOR3xp33_ASAP7_75t_L g811 ( .A(n_812), .B(n_818), .C(n_820), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_816), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_824), .B1(n_825), .B2(n_829), .Y(n_821) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_822), .A2(n_1012), .B1(n_1048), .B2(n_1049), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1059 ( .A1(n_822), .A2(n_1060), .B1(n_1061), .B2(n_1062), .Y(n_1059) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g985 ( .A(n_823), .Y(n_985) );
OAI22xp33_ASAP7_75t_L g861 ( .A1(n_825), .A2(n_839), .B1(n_862), .B2(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g1061 ( .A(n_826), .Y(n_1061) );
INVx2_ASAP7_75t_L g1100 ( .A(n_826), .Y(n_1100) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
BUFx3_ASAP7_75t_L g841 ( .A(n_827), .Y(n_841) );
BUFx6f_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AND2x2_ASAP7_75t_L g844 ( .A(n_845), .B(n_873), .Y(n_844) );
NOR3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_853), .C(n_855), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_850), .Y(n_846) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_858), .B1(n_859), .B2(n_860), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_858), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_860), .A2(n_1095), .B1(n_1096), .B2(n_1097), .Y(n_1094) );
INVx3_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
A2O1A1Ixp33_ASAP7_75t_L g1383 ( .A1(n_886), .A2(n_1031), .B(n_1115), .C(n_1354), .Y(n_1383) );
INVx1_ASAP7_75t_L g999 ( .A(n_890), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_892), .B1(n_945), .B2(n_998), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
XNOR2x1_ASAP7_75t_L g893 ( .A(n_894), .B(n_895), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g1174 ( .A1(n_894), .A2(n_1175), .B1(n_1176), .B2(n_1177), .Y(n_1174) );
OR2x2_ASAP7_75t_L g895 ( .A(n_896), .B(n_917), .Y(n_895) );
INVx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_913), .B1(n_915), .B2(n_916), .Y(n_911) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_935), .C(n_944), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_923), .B1(n_924), .B2(n_925), .Y(n_921) );
INVx2_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx2_ASAP7_75t_SL g926 ( .A(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVxp67_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_SL g998 ( .A(n_945), .Y(n_998) );
XNOR2x1_ASAP7_75t_L g945 ( .A(n_946), .B(n_997), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_974), .Y(n_946) );
AOI31xp33_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_958), .A3(n_970), .B(n_973), .Y(n_949) );
OAI211xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B(n_956), .C(n_957), .Y(n_953) );
OAI221xp5_ASAP7_75t_L g1380 ( .A1(n_955), .A2(n_1022), .B1(n_1350), .B2(n_1356), .C(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
NOR3xp33_ASAP7_75t_SL g974 ( .A(n_975), .B(n_981), .C(n_983), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_978), .Y(n_975) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1001), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1073), .B1(n_1121), .B2(n_1122), .Y(n_1001) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1002), .Y(n_1121) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
NAND4xp25_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1044), .C(n_1063), .D(n_1068), .Y(n_1004) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx2_ASAP7_75t_SL g1038 ( .A(n_1011), .Y(n_1038) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1017 ( .A(n_1018), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1021), .B1(n_1022), .B2(n_1024), .C(n_1025), .Y(n_1019) );
INVx2_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
AOI21xp5_ASAP7_75t_L g1044 ( .A1(n_1024), .A2(n_1045), .B(n_1046), .Y(n_1044) );
NAND3xp33_ASAP7_75t_SL g1026 ( .A(n_1027), .B(n_1032), .C(n_1039), .Y(n_1026) );
A2O1A1Ixp33_ASAP7_75t_SL g1027 ( .A1(n_1028), .A2(n_1029), .B(n_1030), .C(n_1031), .Y(n_1027) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
BUFx2_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1056), .B1(n_1057), .B2(n_1058), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1066), .Y(n_1063) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1073), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
XNOR2x1_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1076), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1102), .Y(n_1076) );
NOR3xp33_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1086), .C(n_1087), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1082), .Y(n_1078) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1108), .C(n_1113), .Y(n_1103) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1117), .Y(n_1389) );
OAI21xp33_ASAP7_75t_SL g1124 ( .A1(n_1125), .A2(n_1338), .B(n_1340), .Y(n_1124) );
NOR2x1_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1304), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1255), .Y(n_1126) );
NOR4xp25_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1197), .C(n_1217), .D(n_1233), .Y(n_1127) );
AOI21xp33_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1181), .B(n_1185), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1150), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1130), .B(n_1182), .Y(n_1261) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1130), .Y(n_1299) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1131), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1131), .B(n_1263), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1131), .B(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1131), .Y(n_1329) );
HB1xp67_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1132), .B(n_1204), .Y(n_1203) );
INVx2_ASAP7_75t_SL g1216 ( .A(n_1132), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1132), .B(n_1204), .Y(n_1231) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1133), .Y(n_1195) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1133), .Y(n_1248) );
AND2x4_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1137), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1134), .B(n_1137), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1407 ( .A(n_1134), .Y(n_1407) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
AND2x4_ASAP7_75t_L g1139 ( .A(n_1135), .B(n_1137), .Y(n_1139) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1136), .B(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1138), .Y(n_1146) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1139), .Y(n_1171) );
INVx1_ASAP7_75t_SL g1177 ( .A(n_1139), .Y(n_1177) );
OAI22xp33_ASAP7_75t_L g1140 ( .A1(n_1141), .A2(n_1142), .B1(n_1147), .B2(n_1148), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_1142), .A2(n_1148), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
OAI22xp33_ASAP7_75t_L g1188 ( .A1(n_1142), .A2(n_1189), .B1(n_1190), .B2(n_1191), .Y(n_1188) );
BUFx3_ASAP7_75t_L g1252 ( .A(n_1142), .Y(n_1252) );
BUFx6f_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_1143), .A2(n_1148), .B1(n_1164), .B2(n_1165), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1145), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1144), .B(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1144), .Y(n_1157) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1145), .Y(n_1156) );
HB1xp67_ASAP7_75t_L g1409 ( .A(n_1146), .Y(n_1409) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1148), .Y(n_1192) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1149), .Y(n_1159) );
A2O1A1Ixp33_ASAP7_75t_L g1197 ( .A1(n_1150), .A2(n_1198), .B(n_1202), .C(n_1207), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1166), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1151), .B(n_1201), .Y(n_1200) );
OAI21xp5_ASAP7_75t_L g1226 ( .A1(n_1151), .A2(n_1227), .B(n_1228), .Y(n_1226) );
NAND3xp33_ASAP7_75t_L g1281 ( .A(n_1151), .B(n_1239), .C(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1152), .B(n_1167), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1152), .B(n_1173), .Y(n_1309) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1162), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1153), .B(n_1162), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1153), .B(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1153), .Y(n_1221) );
O2A1O1Ixp33_ASAP7_75t_SL g1233 ( .A1(n_1153), .A2(n_1234), .B(n_1237), .C(n_1244), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1153), .B(n_1173), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1160), .Y(n_1153) );
AND2x4_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1157), .Y(n_1155) );
AND2x4_ASAP7_75t_L g1158 ( .A(n_1157), .B(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1161), .Y(n_1175) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1162), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1162), .B(n_1172), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1162), .B(n_1221), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1162), .B(n_1166), .Y(n_1260) );
AOI32xp33_ASAP7_75t_L g1291 ( .A1(n_1162), .A2(n_1223), .A3(n_1275), .B1(n_1292), .B2(n_1293), .Y(n_1291) );
A2O1A1Ixp33_ASAP7_75t_L g1295 ( .A1(n_1162), .A2(n_1167), .B(n_1230), .C(n_1265), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1166), .B(n_1184), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1172), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1167), .B(n_1184), .Y(n_1183) );
NOR2xp33_ASAP7_75t_L g1201 ( .A(n_1167), .B(n_1172), .Y(n_1201) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1167), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1167), .B(n_1187), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1167), .B(n_1236), .Y(n_1235) );
INVx4_ASAP7_75t_L g1273 ( .A(n_1167), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1167), .B(n_1277), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_1167), .B(n_1278), .Y(n_1283) );
OR2x2_ASAP7_75t_L g1332 ( .A(n_1167), .B(n_1309), .Y(n_1332) );
AND2x6_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1169), .Y(n_1167) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_1171), .A2(n_1247), .B1(n_1248), .B2(n_1249), .Y(n_1246) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1171), .Y(n_1339) );
NOR2xp33_ASAP7_75t_L g1182 ( .A(n_1172), .B(n_1183), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1172), .B(n_1209), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1172), .B(n_1210), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1172), .B(n_1243), .Y(n_1301) );
CKINVDCx6p67_ASAP7_75t_R g1172 ( .A(n_1173), .Y(n_1172) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1173), .B(n_1221), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1173), .B(n_1221), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1173), .B(n_1209), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1173), .B(n_1243), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1173), .B(n_1184), .Y(n_1286) );
OAI211xp5_ASAP7_75t_SL g1290 ( .A1(n_1173), .A2(n_1218), .B(n_1291), .C(n_1295), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1173), .B(n_1298), .Y(n_1297) );
OR2x6_ASAP7_75t_SL g1173 ( .A(n_1174), .B(n_1178), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_1177), .A2(n_1194), .B1(n_1195), .B2(n_1196), .Y(n_1193) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1184), .B(n_1273), .Y(n_1298) );
INVx1_ASAP7_75t_SL g1275 ( .A(n_1185), .Y(n_1275) );
INVx3_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1186), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1186), .B(n_1204), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1186), .B(n_1245), .Y(n_1244) );
OAI211xp5_ASAP7_75t_L g1256 ( .A1(n_1186), .A2(n_1257), .B(n_1261), .C(n_1262), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1186), .B(n_1203), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1186), .B(n_1216), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1186), .B(n_1239), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1186), .B(n_1278), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1186), .B(n_1204), .Y(n_1333) );
INVx3_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1187), .B(n_1204), .Y(n_1303) );
OR2x2_ASAP7_75t_L g1336 ( .A(n_1187), .B(n_1231), .Y(n_1336) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1193), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1254 ( .A(n_1191), .Y(n_1254) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
NOR2xp33_ASAP7_75t_L g1328 ( .A(n_1200), .B(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
AOI221xp5_ASAP7_75t_L g1270 ( .A1(n_1203), .A2(n_1271), .B1(n_1274), .B2(n_1279), .C(n_1280), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1203), .B(n_1272), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g1305 ( .A1(n_1203), .A2(n_1306), .B1(n_1312), .B2(n_1315), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1204), .B(n_1216), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1204), .B(n_1216), .Y(n_1236) );
INVx2_ASAP7_75t_L g1239 ( .A(n_1204), .Y(n_1239) );
AND2x4_ASAP7_75t_L g1204 ( .A(n_1205), .B(n_1206), .Y(n_1204) );
OAI21xp5_ASAP7_75t_L g1207 ( .A1(n_1208), .A2(n_1211), .B(n_1214), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1300 ( .A1(n_1208), .A2(n_1264), .B1(n_1273), .B2(n_1301), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1208), .B(n_1273), .Y(n_1326) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1209), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1209), .B(n_1272), .Y(n_1271) );
O2A1O1Ixp33_ASAP7_75t_L g1327 ( .A1(n_1211), .A2(n_1258), .B(n_1319), .C(n_1328), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1213), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1212), .B(n_1224), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1238 ( .A(n_1212), .B(n_1239), .Y(n_1238) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1212), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1214), .B(n_1219), .Y(n_1218) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx2_ASAP7_75t_SL g1278 ( .A(n_1216), .Y(n_1278) );
OAI221xp5_ASAP7_75t_L g1217 ( .A1(n_1218), .A2(n_1220), .B1(n_1222), .B2(n_1225), .C(n_1226), .Y(n_1217) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1220), .Y(n_1224) );
OAI211xp5_ASAP7_75t_SL g1280 ( .A1(n_1220), .A2(n_1225), .B(n_1281), .C(n_1284), .Y(n_1280) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1232), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1230), .B(n_1273), .Y(n_1315) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_1231), .A2(n_1258), .B1(n_1259), .B2(n_1260), .Y(n_1257) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1236), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1240), .Y(n_1237) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1239), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1242), .Y(n_1240) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
CKINVDCx5p33_ASAP7_75t_R g1284 ( .A(n_1245), .Y(n_1284) );
OR2x6_ASAP7_75t_SL g1245 ( .A(n_1246), .B(n_1250), .Y(n_1245) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1252), .B1(n_1253), .B2(n_1254), .Y(n_1250) );
OAI32xp33_ASAP7_75t_L g1255 ( .A1(n_1256), .A2(n_1266), .A3(n_1284), .B1(n_1290), .B2(n_1296), .Y(n_1255) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1258), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1265), .Y(n_1263) );
OAI211xp5_ASAP7_75t_SL g1266 ( .A1(n_1267), .A2(n_1268), .B(n_1270), .C(n_1285), .Y(n_1266) );
OAI21xp33_ASAP7_75t_L g1331 ( .A1(n_1267), .A2(n_1273), .B(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1269), .B(n_1286), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1272), .B(n_1279), .Y(n_1335) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
NOR2xp33_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1276), .Y(n_1274) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1276), .Y(n_1320) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
A2O1A1Ixp33_ASAP7_75t_SL g1304 ( .A1(n_1284), .A2(n_1305), .B(n_1316), .C(n_1330), .Y(n_1304) );
OAI21xp5_ASAP7_75t_L g1285 ( .A1(n_1286), .A2(n_1287), .B(n_1289), .Y(n_1285) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
A2O1A1Ixp33_ASAP7_75t_L g1334 ( .A1(n_1288), .A2(n_1335), .B(n_1336), .C(n_1337), .Y(n_1334) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
O2A1O1Ixp33_ASAP7_75t_SL g1296 ( .A1(n_1297), .A2(n_1299), .B(n_1300), .C(n_1302), .Y(n_1296) );
O2A1O1Ixp33_ASAP7_75t_L g1316 ( .A1(n_1301), .A2(n_1317), .B(n_1320), .C(n_1321), .Y(n_1316) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
NOR2xp33_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1310), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
NOR2xp33_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1314), .Y(n_1312) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
A2O1A1Ixp33_ASAP7_75t_L g1321 ( .A1(n_1322), .A2(n_1323), .B(n_1325), .C(n_1327), .Y(n_1321) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
AOI21xp5_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1333), .B(n_1334), .Y(n_1330) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
HB1xp67_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1345), .Y(n_1398) );
NAND4xp25_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1355), .C(n_1373), .D(n_1393), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1347), .B(n_1351), .Y(n_1346) );
OAI221xp5_ASAP7_75t_L g1358 ( .A1(n_1359), .A2(n_1362), .B1(n_1363), .B2(n_1365), .C(n_1366), .Y(n_1358) );
INVx2_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVx2_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
OAI31xp33_ASAP7_75t_SL g1373 ( .A1(n_1374), .A2(n_1378), .A3(n_1382), .B(n_1391), .Y(n_1373) );
NAND3xp33_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1384), .C(n_1387), .Y(n_1382) );
CKINVDCx8_ASAP7_75t_R g1391 ( .A(n_1392), .Y(n_1391) );
BUFx2_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
INVxp67_ASAP7_75t_SL g1396 ( .A(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1398), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
CKINVDCx5p33_ASAP7_75t_R g1402 ( .A(n_1403), .Y(n_1402) );
A2O1A1Ixp33_ASAP7_75t_L g1405 ( .A1(n_1404), .A2(n_1406), .B(n_1408), .C(n_1410), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
endmodule