module fake_ariane_574_n_4525 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_350, n_291, n_344, n_381, n_426, n_433, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_4525);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_4525;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_4030;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_3619;
wire n_589;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_4013;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_4342;
wire n_691;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_3853;
wire n_2559;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2509;
wire n_4085;
wire n_4382;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2334;
wire n_2135;
wire n_2680;
wire n_4259;
wire n_3264;
wire n_4475;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_4299;
wire n_4283;
wire n_1916;
wire n_2879;
wire n_610;
wire n_4403;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_3745;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_3742;
wire n_2729;
wire n_4302;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_4178;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_3765;
wire n_2006;
wire n_4058;
wire n_952;
wire n_864;
wire n_4090;
wire n_2446;
wire n_1096;
wire n_4116;
wire n_1379;
wire n_2436;
wire n_3517;
wire n_3352;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_3719;
wire n_4363;
wire n_524;
wire n_2731;
wire n_3703;
wire n_634;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_3954;
wire n_3888;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_2238;
wire n_1503;
wire n_2529;
wire n_764;
wire n_2374;
wire n_4103;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_2873;
wire n_2653;
wire n_737;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_3938;
wire n_568;
wire n_2278;
wire n_4028;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_3965;
wire n_1457;
wire n_2482;
wire n_3905;
wire n_4416;
wire n_1682;
wire n_2750;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4439;
wire n_520;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_958;
wire n_945;
wire n_3943;
wire n_3930;
wire n_2554;
wire n_3145;
wire n_3808;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_4321;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_3858;
wire n_4106;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_500;
wire n_754;
wire n_665;
wire n_4260;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_829;
wire n_4148;
wire n_1062;
wire n_738;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_4512;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_3856;
wire n_4132;
wire n_4038;
wire n_2442;
wire n_2735;
wire n_4159;
wire n_953;
wire n_1364;
wire n_4214;
wire n_2390;
wire n_4331;
wire n_1888;
wire n_4500;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_2634;
wire n_3451;
wire n_625;
wire n_557;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_559;
wire n_2233;
wire n_2663;
wire n_495;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_4515;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_3890;
wire n_3830;
wire n_821;
wire n_561;
wire n_770;
wire n_3252;
wire n_1514;
wire n_4143;
wire n_4273;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_3879;
wire n_569;
wire n_4136;
wire n_2078;
wire n_3315;
wire n_3929;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_3999;
wire n_2201;
wire n_4353;
wire n_787;
wire n_4012;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_4176;
wire n_1207;
wire n_4124;
wire n_3606;
wire n_786;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_3859;
wire n_868;
wire n_3474;
wire n_2232;
wire n_4488;
wire n_1847;
wire n_2458;
wire n_4320;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3756;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_4077;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_3870;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_3749;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_620;
wire n_3948;
wire n_1074;
wire n_3230;
wire n_859;
wire n_3793;
wire n_4268;
wire n_1765;
wire n_4031;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_3960;
wire n_4454;
wire n_4147;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_3975;
wire n_4184;
wire n_3828;
wire n_3073;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_1013;
wire n_3883;
wire n_4032;
wire n_4018;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_661;
wire n_4227;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_4117;
wire n_533;
wire n_3049;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3877;
wire n_4284;
wire n_440;
wire n_3913;
wire n_3817;
wire n_3013;
wire n_3612;
wire n_4505;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_3728;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_612;
wire n_3739;
wire n_3962;
wire n_512;
wire n_1597;
wire n_4082;
wire n_4476;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_579;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_3854;
wire n_3861;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_2956;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_4171;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_4119;
wire n_4443;
wire n_1443;
wire n_1021;
wire n_4000;
wire n_3089;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_3458;
wire n_570;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3860;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_490;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3850;
wire n_575;
wire n_546;
wire n_3472;
wire n_503;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_4498;
wire n_772;
wire n_1216;
wire n_4174;
wire n_3126;
wire n_3754;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_4432;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_3958;
wire n_4495;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2326;
wire n_2145;
wire n_1838;
wire n_3485;
wire n_4357;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_4109;
wire n_3777;
wire n_4108;
wire n_4502;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3767;
wire n_3841;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_3280;
wire n_3234;
wire n_3413;
wire n_3692;
wire n_3900;
wire n_2216;
wire n_4115;
wire n_1274;
wire n_3539;
wire n_4394;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_3095;
wire n_947;
wire n_2134;
wire n_3862;
wire n_930;
wire n_1260;
wire n_3698;
wire n_3716;
wire n_4226;
wire n_4513;
wire n_1179;
wire n_468;
wire n_3284;
wire n_3909;
wire n_4311;
wire n_4220;
wire n_2703;
wire n_1442;
wire n_696;
wire n_2926;
wire n_482;
wire n_2620;
wire n_798;
wire n_1833;
wire n_577;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_2791;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_762;
wire n_4378;
wire n_555;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_4180;
wire n_4354;
wire n_4405;
wire n_2970;
wire n_4235;
wire n_3159;
wire n_4459;
wire n_992;
wire n_966;
wire n_955;
wire n_3549;
wire n_3885;
wire n_3914;
wire n_3624;
wire n_4264;
wire n_1182;
wire n_2855;
wire n_794;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_4345;
wire n_3250;
wire n_4223;
wire n_3029;
wire n_2398;
wire n_4233;
wire n_3538;
wire n_3915;
wire n_1376;
wire n_3839;
wire n_513;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_3717;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_3875;
wire n_4029;
wire n_2202;
wire n_2072;
wire n_3852;
wire n_2952;
wire n_3530;
wire n_4206;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_436;
wire n_3000;
wire n_2930;
wire n_2871;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_3937;
wire n_4130;
wire n_2161;
wire n_1418;
wire n_4175;
wire n_746;
wire n_1357;
wire n_1079;
wire n_4170;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_4033;
wire n_615;
wire n_3747;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_4456;
wire n_517;
wire n_1312;
wire n_4508;
wire n_1717;
wire n_3604;
wire n_4045;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_3871;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_3757;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_4272;
wire n_2219;
wire n_3116;
wire n_4141;
wire n_1855;
wire n_3784;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3629;
wire n_3666;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_990;
wire n_3559;
wire n_1903;
wire n_3792;
wire n_867;
wire n_2147;
wire n_4267;
wire n_3479;
wire n_4020;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_3998;
wire n_3724;
wire n_4150;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_3287;
wire n_2167;
wire n_4285;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_4055;
wire n_3980;
wire n_4410;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_632;
wire n_3257;
wire n_477;
wire n_650;
wire n_3741;
wire n_2388;
wire n_4352;
wire n_3730;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_1911;
wire n_3979;
wire n_3912;
wire n_2567;
wire n_3950;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_2695;
wire n_2557;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_3700;
wire n_3727;
wire n_712;
wire n_976;
wire n_3567;
wire n_909;
wire n_4003;
wire n_1392;
wire n_1832;
wire n_767;
wire n_2795;
wire n_2682;
wire n_4307;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_489;
wire n_2294;
wire n_2274;
wire n_4438;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_506;
wire n_3814;
wire n_3812;
wire n_3127;
wire n_3796;
wire n_1731;
wire n_799;
wire n_4433;
wire n_3884;
wire n_1147;
wire n_2829;
wire n_4367;
wire n_4492;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_471;
wire n_965;
wire n_1914;
wire n_4195;
wire n_3760;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_4056;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_3744;
wire n_4015;
wire n_2924;
wire n_1209;
wire n_4022;
wire n_4445;
wire n_1020;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_646;
wire n_4254;
wire n_4462;
wire n_2507;
wire n_4219;
wire n_4484;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_4043;
wire n_4336;
wire n_4451;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_479;
wire n_3936;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_3661;
wire n_2223;
wire n_836;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_2473;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_564;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_3981;
wire n_1247;
wire n_4234;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3867;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_3031;
wire n_2262;
wire n_3179;
wire n_2565;
wire n_3889;
wire n_1237;
wire n_3262;
wire n_4314;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_3699;
wire n_3971;
wire n_4315;
wire n_2120;
wire n_706;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3869;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_4442;
wire n_776;
wire n_2860;
wire n_3816;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_4494;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_1817;
wire n_3711;
wire n_4201;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_3704;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_4296;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_4051;
wire n_2483;
wire n_4242;
wire n_4074;
wire n_3994;
wire n_441;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_637;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_4386;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3917;
wire n_4122;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_4275;
wire n_3774;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_4522;
wire n_2718;
wire n_4263;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_4426;
wire n_3876;
wire n_3615;
wire n_4362;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_3946;
wire n_4243;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_4225;
wire n_3642;
wire n_2237;
wire n_4153;
wire n_2146;
wire n_4274;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_4186;
wire n_1501;
wire n_4089;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3513;
wire n_3498;
wire n_3682;
wire n_2350;
wire n_3881;
wire n_1068;
wire n_1198;
wire n_4096;
wire n_4506;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3759;
wire n_3377;
wire n_487;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_4007;
wire n_1879;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_3961;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_3863;
wire n_2129;
wire n_855;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_3968;
wire n_4133;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_4337;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_4486;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_4359;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_3118;
wire n_4072;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4441;
wire n_1906;
wire n_4323;
wire n_529;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_3922;
wire n_502;
wire n_4447;
wire n_2194;
wire n_2937;
wire n_4293;
wire n_3508;
wire n_1467;
wire n_4039;
wire n_1828;
wire n_4129;
wire n_4458;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_3831;
wire n_1744;
wire n_3335;
wire n_4523;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_3599;
wire n_3618;
wire n_439;
wire n_677;
wire n_604;
wire n_3705;
wire n_3022;
wire n_478;
wire n_703;
wire n_3983;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_681;
wire n_3286;
wire n_4480;
wire n_3734;
wire n_3370;
wire n_874;
wire n_3773;
wire n_3949;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_4247;
wire n_707;
wire n_3974;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_3988;
wire n_3939;
wire n_3788;
wire n_590;
wire n_2075;
wire n_727;
wire n_1726;
wire n_699;
wire n_3263;
wire n_3569;
wire n_2523;
wire n_1945;
wire n_3542;
wire n_3837;
wire n_3835;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1614;
wire n_1162;
wire n_536;
wire n_1377;
wire n_2031;
wire n_545;
wire n_3260;
wire n_3349;
wire n_3761;
wire n_3996;
wire n_4292;
wire n_3819;
wire n_2118;
wire n_3222;
wire n_1740;
wire n_4348;
wire n_1602;
wire n_688;
wire n_3139;
wire n_636;
wire n_2853;
wire n_3350;
wire n_3801;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_3764;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_4374;
wire n_3653;
wire n_3951;
wire n_3868;
wire n_3035;
wire n_3823;
wire n_729;
wire n_887;
wire n_3403;
wire n_4261;
wire n_2218;
wire n_2057;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_4236;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_3942;
wire n_1202;
wire n_4344;
wire n_4084;
wire n_627;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_2618;
wire n_4121;
wire n_3602;
wire n_4216;
wire n_1402;
wire n_957;
wire n_1242;
wire n_3957;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_4393;
wire n_3611;
wire n_3781;
wire n_2217;
wire n_2226;
wire n_3959;
wire n_3984;
wire n_1586;
wire n_4313;
wire n_861;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_1431;
wire n_4389;
wire n_877;
wire n_3995;
wire n_1119;
wire n_4460;
wire n_3713;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_3908;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_2763;
wire n_4297;
wire n_4461;
wire n_4229;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3750;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3492;
wire n_3737;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_3501;
wire n_2516;
wire n_3931;
wire n_4094;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_735;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_527;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_4049;
wire n_4067;
wire n_3896;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_4182;
wire n_4269;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_551;
wire n_3551;
wire n_4521;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_3710;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_3803;
wire n_3766;
wire n_3985;
wire n_1219;
wire n_1711;
wire n_4387;
wire n_1919;
wire n_710;
wire n_2994;
wire n_534;
wire n_2508;
wire n_1791;
wire n_3186;
wire n_4369;
wire n_2124;
wire n_1894;
wire n_2594;
wire n_1239;
wire n_1460;
wire n_3826;
wire n_2266;
wire n_3944;
wire n_3417;
wire n_2449;
wire n_560;
wire n_890;
wire n_4324;
wire n_842;
wire n_3626;
wire n_1898;
wire n_4428;
wire n_451;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_4464;
wire n_4463;
wire n_1793;
wire n_4446;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_3671;
wire n_4396;
wire n_4440;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_4425;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_3696;
wire n_2474;
wire n_4104;
wire n_2623;
wire n_3392;
wire n_982;
wire n_1800;
wire n_915;
wire n_3791;
wire n_1075;
wire n_2008;
wire n_454;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_4034;
wire n_1529;
wire n_4228;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_655;
wire n_2946;
wire n_3166;
wire n_4237;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_4114;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_657;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_3924;
wire n_4081;
wire n_837;
wire n_812;
wire n_2448;
wire n_3997;
wire n_2211;
wire n_4172;
wire n_4040;
wire n_2292;
wire n_4482;
wire n_2480;
wire n_606;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_3795;
wire n_2306;
wire n_509;
wire n_4328;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_3990;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_3953;
wire n_2414;
wire n_4400;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_4069;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_4280;
wire n_456;
wire n_1867;
wire n_3993;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_704;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_4113;
wire n_2696;
wire n_4351;
wire n_4424;
wire n_3340;
wire n_4429;
wire n_4192;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_3977;
wire n_1400;
wire n_4112;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3735;
wire n_3486;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_608;
wire n_2494;
wire n_4524;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_4071;
wire n_1329;
wire n_4436;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_4160;
wire n_4035;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_3964;
wire n_2540;
wire n_4190;
wire n_3836;
wire n_3302;
wire n_1605;
wire n_4137;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_4009;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_811;
wire n_4145;
wire n_3097;
wire n_4395;
wire n_624;
wire n_3507;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_3864;
wire n_4385;
wire n_2939;
wire n_3425;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_3748;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_4050;
wire n_3173;
wire n_480;
wire n_1327;
wire n_3732;
wire n_1475;
wire n_642;
wire n_2106;
wire n_1804;
wire n_1406;
wire n_595;
wire n_4306;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_602;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_4006;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_592;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_4288;
wire n_3452;
wire n_2091;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_4098;
wire n_4312;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_3789;
wire n_805;
wire n_4319;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3811;
wire n_3422;
wire n_4511;
wire n_4358;
wire n_1658;
wire n_4200;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_695;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_2785;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_4289;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_3925;
wire n_2928;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_3746;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_3780;
wire n_1657;
wire n_878;
wire n_2857;
wire n_3694;
wire n_4118;
wire n_1784;
wire n_3110;
wire n_3857;
wire n_771;
wire n_3787;
wire n_4025;
wire n_4239;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_3157;
wire n_3893;
wire n_3753;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_3702;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_4076;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3495;
wire n_3107;
wire n_3843;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_4065;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_3708;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3543;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_686;
wire n_4279;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_4330;
wire n_1130;
wire n_1450;
wire n_4152;
wire n_3718;
wire n_2022;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_3740;
wire n_4343;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_3976;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_515;
wire n_3381;
wire n_807;
wire n_3455;
wire n_3736;
wire n_4466;
wire n_891;
wire n_3313;
wire n_885;
wire n_1659;
wire n_3955;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3907;
wire n_3086;
wire n_4332;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_4281;
wire n_3317;
wire n_3945;
wire n_3726;
wire n_3336;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_4419;
wire n_1151;
wire n_554;
wire n_960;
wire n_4420;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_714;
wire n_3605;
wire n_3560;
wire n_2170;
wire n_3345;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4404;
wire n_725;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3840;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_4372;
wire n_4097;
wire n_4054;
wire n_3809;
wire n_4162;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_4377;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2477;
wire n_2314;
wire n_2279;
wire n_3169;
wire n_594;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_4173;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4301;
wire n_3573;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_3291;
wire n_3654;
wire n_4188;
wire n_2001;
wire n_1047;
wire n_3783;
wire n_2506;
wire n_1472;
wire n_4399;
wire n_2413;
wire n_4008;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_4140;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2796;
wire n_2173;
wire n_3982;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3973;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_3755;
wire n_2947;
wire n_1367;
wire n_3842;
wire n_4202;
wire n_2044;
wire n_928;
wire n_4304;
wire n_3886;
wire n_1153;
wire n_465;
wire n_3769;
wire n_4078;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_4437;
wire n_1192;
wire n_3738;
wire n_894;
wire n_3098;
wire n_1380;
wire n_4503;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_562;
wire n_4070;
wire n_2020;
wire n_748;
wire n_3987;
wire n_2310;
wire n_510;
wire n_4249;
wire n_4418;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_4125;
wire n_2711;
wire n_1023;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_4139;
wire n_914;
wire n_689;
wire n_1116;
wire n_4327;
wire n_3921;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_4011;
wire n_467;
wire n_1511;
wire n_2177;
wire n_3695;
wire n_2713;
wire n_1422;
wire n_3800;
wire n_2766;
wire n_1965;
wire n_644;
wire n_3462;
wire n_4450;
wire n_4196;
wire n_1197;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_497;
wire n_3733;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_3967;
wire n_3731;
wire n_4291;
wire n_538;
wire n_2845;
wire n_4151;
wire n_1517;
wire n_2036;
wire n_4412;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_588;
wire n_3358;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_3920;
wire n_1307;
wire n_4368;
wire n_3444;
wire n_4370;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_4091;
wire n_3851;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3096;
wire n_667;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_4430;
wire n_1398;
wire n_1921;
wire n_4166;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_1370;
wire n_1603;
wire n_728;
wire n_4191;
wire n_4409;
wire n_4478;
wire n_2401;
wire n_2935;
wire n_4246;
wire n_715;
wire n_889;
wire n_3822;
wire n_3255;
wire n_4355;
wire n_1066;
wire n_1549;
wire n_3818;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_3827;
wire n_2478;
wire n_685;
wire n_911;
wire n_4061;
wire n_2658;
wire n_623;
wire n_3587;
wire n_3509;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1948;
wire n_1534;
wire n_3006;
wire n_2767;
wire n_4518;
wire n_4155;
wire n_810;
wire n_3376;
wire n_4278;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_617;
wire n_3770;
wire n_4375;
wire n_2396;
wire n_3243;
wire n_543;
wire n_3368;
wire n_1362;
wire n_4326;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3865;
wire n_3123;
wire n_2692;
wire n_683;
wire n_601;
wire n_565;
wire n_3927;
wire n_628;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_4308;
wire n_743;
wire n_1194;
wire n_2862;
wire n_4060;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_3790;
wire n_907;
wire n_2749;
wire n_2592;
wire n_1454;
wire n_660;
wire n_464;
wire n_3490;
wire n_2459;
wire n_962;
wire n_4413;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_747;
wire n_4241;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_3101;
wire n_918;
wire n_1968;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_3288;
wire n_3251;
wire n_4093;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_4123;
wire n_1038;
wire n_3603;
wire n_3723;
wire n_4135;
wire n_2371;
wire n_1978;
wire n_4257;
wire n_571;
wire n_4282;
wire n_4294;
wire n_3880;
wire n_4341;
wire n_3720;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3904;
wire n_3887;
wire n_593;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_4027;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_3405;
wire n_4309;
wire n_2313;
wire n_609;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_4126;
wire n_4164;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_4333;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_519;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_3978;
wire n_1767;
wire n_1040;
wire n_674;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_4138;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_3409;
wire n_4079;
wire n_3522;
wire n_3583;
wire n_4381;
wire n_4088;
wire n_4316;
wire n_2882;
wire n_2303;
wire n_4469;
wire n_2669;
wire n_3540;
wire n_3911;
wire n_4455;
wire n_3241;
wire n_4384;
wire n_3899;
wire n_4366;
wire n_1157;
wire n_1584;
wire n_3802;
wire n_848;
wire n_1664;
wire n_3481;
wire n_629;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_1814;
wire n_4210;
wire n_532;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_4041;
wire n_2174;
wire n_2688;
wire n_540;
wire n_692;
wire n_2624;
wire n_3442;
wire n_4208;
wire n_3972;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_3926;
wire n_4209;
wire n_984;
wire n_1687;
wire n_4457;
wire n_2073;
wire n_2150;
wire n_4481;
wire n_4004;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_3992;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_4350;
wire n_2189;
wire n_2648;
wire n_621;
wire n_3305;
wire n_1587;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_2340;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_3991;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_3786;
wire n_697;
wire n_2828;
wire n_4212;
wire n_4270;
wire n_622;
wire n_1626;
wire n_3436;
wire n_4509;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3806;
wire n_4204;
wire n_3553;
wire n_4044;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3833;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_3751;
wire n_4388;
wire n_3402;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_4477;
wire n_1621;
wire n_4110;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_4411;
wire n_1221;
wire n_4217;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_4271;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_4317;
wire n_4406;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_580;
wire n_3664;
wire n_1579;
wire n_494;
wire n_2809;
wire n_4218;
wire n_2181;
wire n_3550;
wire n_434;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_3722;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_3969;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_4068;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_3873;
wire n_2270;
wire n_3470;
wire n_4163;
wire n_3785;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_2428;
wire n_994;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3844;
wire n_3259;
wire n_4262;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3714;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3721;
wire n_3677;
wire n_1564;
wire n_2010;
wire n_3676;
wire n_1054;
wire n_508;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3701;
wire n_3109;
wire n_3706;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_3989;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_1057;
wire n_4131;
wire n_2487;
wire n_1834;
wire n_4215;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_4158;
wire n_1411;
wire n_1359;
wire n_4286;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_558;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3558;
wire n_3576;
wire n_3782;
wire n_4231;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_4435;
wire n_783;
wire n_4053;
wire n_2550;
wire n_1127;
wire n_556;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3963;
wire n_4318;
wire n_3658;
wire n_581;
wire n_3091;
wire n_1024;
wire n_830;
wire n_4496;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_4177;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_3521;
wire n_3855;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_4083;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_4105;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_3940;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_679;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_443;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_3897;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_4005;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_4230;
wire n_4181;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_445;
wire n_3360;
wire n_4470;
wire n_4187;
wire n_1930;
wire n_3687;
wire n_765;
wire n_1809;
wire n_2787;
wire n_4092;
wire n_3585;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_4037;
wire n_1268;
wire n_3804;
wire n_2676;
wire n_4255;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_4057;
wire n_2770;
wire n_631;
wire n_3847;
wire n_1170;
wire n_2724;
wire n_4073;
wire n_3575;
wire n_4347;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_3633;
wire n_898;
wire n_857;
wire n_3042;
wire n_968;
wire n_1067;
wire n_4144;
wire n_4335;
wire n_1323;
wire n_1235;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_4001;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_4167;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_633;
wire n_900;
wire n_4142;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_4021;
wire n_1285;
wire n_3379;
wire n_4379;
wire n_3111;
wire n_761;
wire n_733;
wire n_2212;
wire n_3838;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_4059;
wire n_4434;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_668;
wire n_4499;
wire n_2569;
wire n_758;
wire n_4504;
wire n_4019;
wire n_4199;
wire n_3691;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_3743;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_2897;
wire n_4339;
wire n_1322;
wire n_3273;
wire n_4497;
wire n_3829;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_4510;
wire n_835;
wire n_3155;
wire n_4300;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_701;
wire n_1125;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_2358;
wire n_3316;
wire n_4023;
wire n_4472;
wire n_4253;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2580;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_485;
wire n_1792;
wire n_4064;
wire n_504;
wire n_3351;
wire n_2062;
wire n_483;
wire n_4489;
wire n_435;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_3901;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1459;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_4519;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_759;
wire n_567;
wire n_4156;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_3693;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_614;
wire n_3776;
wire n_4066;
wire n_2775;
wire n_3903;
wire n_1212;
wire n_3581;
wire n_3778;
wire n_831;
wire n_3681;
wire n_4310;
wire n_3933;
wire n_3970;
wire n_4371;
wire n_778;
wire n_2351;
wire n_1619;
wire n_4322;
wire n_3303;
wire n_2260;
wire n_550;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_1902;
wire n_2206;
wire n_997;
wire n_2784;
wire n_635;
wire n_3898;
wire n_4414;
wire n_2541;
wire n_694;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_4448;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_3768;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_4295;
wire n_3932;
wire n_2101;
wire n_1934;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_4193;
wire n_4100;
wire n_4507;
wire n_2104;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_1576;
wire n_1533;
wire n_1806;
wire n_671;
wire n_2552;
wire n_1470;
wire n_3445;
wire n_4087;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_4473;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_3729;
wire n_4398;
wire n_3253;
wire n_4471;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_3952;
wire n_4392;
wire n_1275;
wire n_3103;
wire n_488;
wire n_3018;
wire n_4238;
wire n_904;
wire n_505;
wire n_4365;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_498;
wire n_3028;
wire n_1875;
wire n_4349;
wire n_1059;
wire n_3148;
wire n_3775;
wire n_2736;
wire n_2429;
wire n_2108;
wire n_684;
wire n_3966;
wire n_4397;
wire n_4449;
wire n_3285;
wire n_3824;
wire n_3825;
wire n_4198;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_539;
wire n_1150;
wire n_4266;
wire n_977;
wire n_449;
wire n_2339;
wire n_3846;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_4373;
wire n_4407;
wire n_1497;
wire n_4189;
wire n_1866;
wire n_3874;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_4165;
wire n_4154;
wire n_4479;
wire n_2056;
wire n_2852;
wire n_459;
wire n_1136;
wire n_2515;
wire n_4390;
wire n_3845;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_4107;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_711;
wire n_4380;
wire n_4361;
wire n_3941;
wire n_734;
wire n_1915;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4258;
wire n_2846;
wire n_3371;
wire n_1781;
wire n_709;
wire n_2917;
wire n_3137;
wire n_4250;
wire n_2544;
wire n_809;
wire n_3143;
wire n_3194;
wire n_3690;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_3872;
wire n_4415;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_4232;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_2097;
wire n_1982;
wire n_662;
wire n_641;
wire n_3461;
wire n_3366;
wire n_2430;
wire n_2504;
wire n_910;
wire n_4211;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_3094;
wire n_4276;
wire n_3441;
wire n_4203;
wire n_3020;
wire n_4146;
wire n_4002;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_3815;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_4408;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3752;
wire n_4483;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_448;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3820;
wire n_3555;
wire n_3072;
wire n_4128;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_450;
wire n_4036;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3655;
wire n_4487;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_3918;
wire n_716;
wire n_4010;
wire n_4329;
wire n_1571;
wire n_4501;
wire n_1698;
wire n_3902;
wire n_4101;
wire n_3866;
wire n_1337;
wire n_3763;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_3244;
wire n_4383;
wire n_3499;
wire n_4391;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1168;
wire n_1821;
wire n_4095;
wire n_4444;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3794;
wire n_3762;
wire n_3947;
wire n_3910;
wire n_4485;
wire n_656;
wire n_492;
wire n_574;
wire n_4205;
wire n_3593;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_664;
wire n_2995;
wire n_3361;
wire n_3293;
wire n_4287;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_4356;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_3707;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3779;
wire n_3895;
wire n_3149;
wire n_537;
wire n_1063;
wire n_3934;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_991;
wire n_4338;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_4224;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_3834;
wire n_2761;
wire n_2357;
wire n_4303;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_4520;
wire n_1328;
wire n_895;
wire n_4161;
wire n_2875;
wire n_1639;
wire n_583;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_626;
wire n_4042;
wire n_1581;
wire n_4244;
wire n_3849;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_3709;
wire n_4465;
wire n_3398;
wire n_1634;
wire n_4265;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3557;
wire n_3725;
wire n_3592;
wire n_3986;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_4026;
wire n_4245;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3894;
wire n_3202;
wire n_1794;
wire n_4290;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_3772;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_4149;
wire n_4120;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_2361;
wire n_1001;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3075;
wire n_3030;
wire n_3505;
wire n_4277;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_3547;
wire n_4014;
wire n_3771;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_4516;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_4222;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_3821;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_4016;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_548;
wire n_3427;
wire n_2336;
wire n_523;
wire n_1662;
wire n_3162;
wire n_457;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3483;
wire n_3430;
wire n_4046;
wire n_4467;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_3935;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_4047;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_4063;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_4493;
wire n_3798;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_4248;
wire n_1672;
wire n_4376;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_3832;
wire n_893;
wire n_3525;
wire n_3308;
wire n_3712;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_4134;
wire n_2037;
wire n_4305;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_573;
wire n_796;
wire n_2851;
wire n_2823;
wire n_4017;
wire n_531;
wire n_2345;
wire n_4417;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g434 ( 
.A(n_107),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_380),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_126),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_66),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_35),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_145),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_407),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_310),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_432),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_101),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_116),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_433),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_101),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_192),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_88),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_11),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_110),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_41),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_191),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_401),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_236),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_110),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_304),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_280),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_35),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_140),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_347),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_10),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_406),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_290),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_69),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_431),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_411),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_346),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_377),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_42),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_284),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_157),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_341),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_251),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_279),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_131),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_45),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_17),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_113),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_120),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_41),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_373),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_8),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_182),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_317),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_62),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_308),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_88),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_309),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_345),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_202),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_370),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_168),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_173),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_26),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_244),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_224),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_141),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_368),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_141),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_154),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_117),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_12),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_376),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_46),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_196),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_89),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_259),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_23),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_351),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_425),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_104),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_282),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_385),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_189),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_120),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_261),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_172),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_405),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_153),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_423),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_183),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_418),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_49),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_70),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_275),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_188),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_62),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_209),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_77),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_353),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_313),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_358),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_51),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_32),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_400),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_174),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_378),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_391),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_307),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_38),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_138),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_126),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_225),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_382),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_209),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_21),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_323),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_17),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_333),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_235),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_154),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_53),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_233),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_402),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_312),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_179),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_305),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_20),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_338),
.Y(n_560)
);

CKINVDCx14_ASAP7_75t_R g561 ( 
.A(n_403),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_177),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_241),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_180),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_159),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_167),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_127),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_191),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_340),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_11),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_125),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_225),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_426),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_314),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_67),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_266),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_289),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_14),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_393),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_146),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_386),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_265),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_107),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_20),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_53),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_86),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_242),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_116),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_186),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_5),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_422),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_182),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_77),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_409),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_112),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_138),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_361),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_410),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_211),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_252),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_80),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_12),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_84),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_429),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_248),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_360),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g607 ( 
.A(n_246),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_181),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_146),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_63),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_319),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_383),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_68),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_369),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_231),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_281),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_416),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_106),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_232),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_260),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_356),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_106),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_134),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_32),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_30),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_212),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_51),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_277),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_90),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_348),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_99),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_303),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_178),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_269),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_339),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_179),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_8),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_223),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_253),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_417),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_421),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_177),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_390),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_57),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_66),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_10),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_244),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_47),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_34),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_184),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_75),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_85),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_216),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_145),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_171),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_296),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_413),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_93),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_188),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_388),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_371),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_399),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_322),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_350),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_15),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_70),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_135),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_392),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_111),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_52),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_193),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_214),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_23),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_419),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_56),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_184),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_189),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_343),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g679 ( 
.A(n_223),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_253),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_160),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_6),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_424),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_89),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_213),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_427),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_363),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_123),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_408),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_65),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_252),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_237),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_102),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_87),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_132),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_228),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_367),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_140),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_287),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_430),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_334),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_283),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_124),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_206),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_6),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_50),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_365),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_91),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_99),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_153),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_113),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_357),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_68),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_213),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_197),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_14),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_245),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_57),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_109),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_117),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_398),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_387),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_39),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_76),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_344),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_285),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_201),
.Y(n_727)
);

CKINVDCx16_ASAP7_75t_R g728 ( 
.A(n_397),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_24),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_221),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_187),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_58),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_167),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_404),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_112),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_1),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_412),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_3),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_220),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_30),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_169),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_301),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_428),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_420),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_111),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_224),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_239),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_150),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_2),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_9),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_119),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_22),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_375),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_297),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_236),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_415),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_355),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_204),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_208),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_210),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_306),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_249),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_230),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_31),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_530),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_608),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_608),
.Y(n_767)
);

CKINVDCx16_ASAP7_75t_R g768 ( 
.A(n_679),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_439),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_728),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_691),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_691),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_530),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_434),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_434),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_438),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_438),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_453),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_728),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_442),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_448),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_454),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_454),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_459),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_454),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_448),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_679),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_454),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_449),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_581),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_449),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_451),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_451),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_442),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_452),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_452),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_470),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_460),
.Y(n_798)
);

BUFx8_ASAP7_75t_SL g799 ( 
.A(n_480),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_460),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_563),
.B(n_0),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_465),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_465),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_439),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_442),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_476),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_476),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_537),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_481),
.Y(n_809)
);

CKINVDCx14_ASAP7_75t_R g810 ( 
.A(n_446),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_581),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_458),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_537),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_481),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_486),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_486),
.Y(n_816)
);

INVx4_ASAP7_75t_R g817 ( 
.A(n_656),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_581),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_493),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_493),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_537),
.Y(n_821)
);

BUFx4f_ASAP7_75t_SL g822 ( 
.A(n_457),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_458),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_581),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_657),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_657),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_657),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_495),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_495),
.Y(n_829)
);

INVxp67_ASAP7_75t_SL g830 ( 
.A(n_537),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_497),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_497),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_500),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_500),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_657),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_442),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_507),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_474),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_507),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_488),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_607),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_468),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_436),
.B(n_0),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_516),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_539),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_516),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_529),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_634),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_529),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_471),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_491),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_544),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_683),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_544),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_552),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_471),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_L g857 ( 
.A(n_436),
.B(n_1),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_552),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_554),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_554),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_757),
.Y(n_861)
);

CKINVDCx16_ASAP7_75t_R g862 ( 
.A(n_498),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_559),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_559),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_518),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_562),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_561),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_477),
.B(n_2),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_437),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_537),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_562),
.Y(n_871)
);

CKINVDCx16_ASAP7_75t_R g872 ( 
.A(n_498),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_572),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_567),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_440),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_572),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_567),
.Y(n_877)
);

INVxp67_ASAP7_75t_SL g878 ( 
.A(n_572),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_549),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_572),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_575),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_473),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_444),
.Y(n_883)
);

INVxp33_ASAP7_75t_L g884 ( 
.A(n_575),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_584),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_445),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_447),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_584),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_586),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_586),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_603),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_450),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_603),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_610),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_455),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_477),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_509),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_610),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_613),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_613),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_619),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_456),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_572),
.Y(n_903)
);

NOR2xp67_ASAP7_75t_L g904 ( 
.A(n_509),
.B(n_3),
.Y(n_904)
);

NOR2xp67_ASAP7_75t_L g905 ( 
.A(n_525),
.B(n_4),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_442),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_473),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_619),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_678),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_622),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_551),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_462),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_622),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_498),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_472),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_478),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_483),
.Y(n_917)
);

INVxp33_ASAP7_75t_L g918 ( 
.A(n_625),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_625),
.Y(n_919)
);

CKINVDCx16_ASAP7_75t_R g920 ( 
.A(n_498),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_650),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_650),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_677),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_484),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_475),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_677),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_593),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_682),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_593),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_494),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_682),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_525),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_475),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_593),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_496),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_501),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_564),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_502),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_692),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_692),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_693),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_693),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_694),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_694),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_593),
.Y(n_945)
);

BUFx5_ASAP7_75t_L g946 ( 
.A(n_485),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_503),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_695),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_695),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_505),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_703),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_506),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_515),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_520),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_703),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_713),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_522),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_524),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_713),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_717),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_678),
.Y(n_961)
);

INVxp67_ASAP7_75t_SL g962 ( 
.A(n_593),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_678),
.Y(n_963)
);

NOR2xp67_ASAP7_75t_L g964 ( 
.A(n_708),
.B(n_4),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_717),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_730),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_528),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_730),
.Y(n_968)
);

CKINVDCx16_ASAP7_75t_R g969 ( 
.A(n_541),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_708),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_736),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_736),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_747),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_747),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_633),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_749),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_749),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_763),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_763),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_512),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_512),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_583),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_633),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_678),
.Y(n_984)
);

INVxp67_ASAP7_75t_SL g985 ( 
.A(n_633),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_535),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_534),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_658),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_542),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_535),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_570),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_669),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_570),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_596),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_678),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_596),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_618),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_633),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_618),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_629),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_629),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_543),
.Y(n_1002)
);

BUFx5_ASAP7_75t_L g1003 ( 
.A(n_485),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_649),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_649),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_651),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_651),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_667),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_667),
.Y(n_1009)
);

INVxp67_ASAP7_75t_SL g1010 ( 
.A(n_633),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_723),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_546),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_547),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_723),
.Y(n_1014)
);

NOR2xp67_ASAP7_75t_L g1015 ( 
.A(n_735),
.B(n_5),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_735),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_711),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_698),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_729),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_553),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_698),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_698),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_698),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_698),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_565),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_487),
.Y(n_1026)
);

BUFx5_ASAP7_75t_L g1027 ( 
.A(n_487),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_541),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_758),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_489),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_489),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_490),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_541),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_490),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_741),
.B(n_7),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_479),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_526),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_566),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_568),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_541),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_571),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_526),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_531),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_531),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_578),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_536),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_536),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_550),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_580),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_557),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_550),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_585),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_527),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_604),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_587),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_588),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_555),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_555),
.Y(n_1058)
);

CKINVDCx16_ASAP7_75t_R g1059 ( 
.A(n_557),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_589),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_569),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_590),
.Y(n_1062)
);

INVxp67_ASAP7_75t_SL g1063 ( 
.A(n_569),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_592),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_573),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_573),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_582),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_637),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_595),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_599),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_582),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_611),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_611),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_617),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_617),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_600),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_557),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_601),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_620),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_620),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_602),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_632),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_605),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_632),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_640),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_640),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_641),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_557),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_641),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_643),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_643),
.Y(n_1091)
);

BUFx5_ASAP7_75t_L g1092 ( 
.A(n_662),
.Y(n_1092)
);

CKINVDCx16_ASAP7_75t_R g1093 ( 
.A(n_672),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_609),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_662),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_615),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_623),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_663),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_663),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_672),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_672),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_604),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_668),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_668),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_721),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_721),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_722),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_624),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_722),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_626),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_734),
.B(n_7),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_627),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_734),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_742),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_631),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_742),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_636),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_743),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_672),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_642),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_685),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_743),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_754),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_754),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_685),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_761),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_761),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_638),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_1054),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_842),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_842),
.Y(n_1131)
);

INVxp67_ASAP7_75t_SL g1132 ( 
.A(n_830),
.Y(n_1132)
);

INVxp67_ASAP7_75t_L g1133 ( 
.A(n_1036),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_845),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_797),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_873),
.Y(n_1136)
);

NOR2xp67_ASAP7_75t_L g1137 ( 
.A(n_867),
.B(n_656),
.Y(n_1137)
);

INVxp67_ASAP7_75t_L g1138 ( 
.A(n_1068),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_845),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_851),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_797),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_865),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_865),
.Y(n_1143)
);

CKINVDCx20_ASAP7_75t_R g1144 ( 
.A(n_911),
.Y(n_1144)
);

CKINVDCx14_ASAP7_75t_R g1145 ( 
.A(n_810),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_878),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_848),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_848),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_962),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_985),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_853),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_911),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_853),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_1010),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_937),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_823),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_937),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_1054),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_861),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_867),
.B(n_464),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1120),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_R g1162 ( 
.A(n_782),
.B(n_435),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_982),
.Y(n_1163)
);

INVxp67_ASAP7_75t_SL g1164 ( 
.A(n_766),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_861),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_823),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_882),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_822),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_882),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_780),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_799),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_782),
.B(n_697),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_879),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1019),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_982),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_783),
.B(n_538),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1126),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_770),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_770),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_779),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1126),
.Y(n_1181)
);

NOR2xp67_ASAP7_75t_L g1182 ( 
.A(n_783),
.B(n_697),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_774),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_988),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_884),
.B(n_685),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_779),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_775),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_776),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_777),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_781),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_786),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_785),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_785),
.B(n_510),
.Y(n_1193)
);

CKINVDCx16_ASAP7_75t_R g1194 ( 
.A(n_862),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_988),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_789),
.Y(n_1196)
);

NOR2xp67_ASAP7_75t_L g1197 ( 
.A(n_788),
.B(n_441),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_788),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_790),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_791),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_992),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_792),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_992),
.Y(n_1203)
);

INVxp67_ASAP7_75t_SL g1204 ( 
.A(n_769),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_869),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_793),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_869),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_795),
.Y(n_1208)
);

CKINVDCx14_ASAP7_75t_R g1209 ( 
.A(n_790),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_875),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_808),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_L g1212 ( 
.A(n_811),
.B(n_818),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_1017),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_1017),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_811),
.B(n_443),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_1029),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1029),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_796),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_787),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_SL g1220 ( 
.A(n_773),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_798),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_800),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_787),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_875),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_802),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_883),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_883),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_803),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_807),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_768),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_809),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_814),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_840),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_841),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_1045),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_808),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_815),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1033),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1033),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_816),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_838),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_838),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_819),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_886),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_886),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_887),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_887),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_820),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_828),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1040),
.Y(n_1250)
);

BUFx2_ASAP7_75t_SL g1251 ( 
.A(n_1040),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_829),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_818),
.B(n_712),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_831),
.Y(n_1254)
);

INVxp33_ASAP7_75t_SL g1255 ( 
.A(n_824),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_824),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1050),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_825),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1050),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_832),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1077),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_833),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_769),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_892),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_892),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_834),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_L g1267 ( 
.A(n_825),
.B(n_461),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_837),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1054),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1077),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_839),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_844),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1101),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_895),
.Y(n_1274)
);

INVxp67_ASAP7_75t_L g1275 ( 
.A(n_1045),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_846),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_895),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_902),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_847),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_826),
.B(n_579),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_852),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_826),
.Y(n_1282)
);

CKINVDCx16_ASAP7_75t_R g1283 ( 
.A(n_872),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_854),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_855),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1101),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_858),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_859),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1128),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_860),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_864),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_866),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1119),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_871),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_L g1295 ( 
.A(n_827),
.B(n_463),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_874),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_877),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_881),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_902),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1128),
.Y(n_1300)
);

INVxp33_ASAP7_75t_L g1301 ( 
.A(n_950),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_885),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_912),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_888),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_889),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_912),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_890),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_778),
.B(n_715),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_804),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1069),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_778),
.B(n_718),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1119),
.Y(n_1312)
);

INVxp33_ASAP7_75t_SL g1313 ( 
.A(n_827),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_915),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_1121),
.Y(n_1315)
);

INVxp67_ASAP7_75t_L g1316 ( 
.A(n_1078),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_813),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1121),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1054),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_891),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1117),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1125),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_804),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_835),
.B(n_628),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1125),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_914),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_893),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_894),
.Y(n_1328)
);

NOR2xp67_ASAP7_75t_L g1329 ( 
.A(n_835),
.B(n_466),
.Y(n_1329)
);

NOR2xp67_ASAP7_75t_L g1330 ( 
.A(n_1028),
.B(n_467),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_920),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1057),
.B(n_712),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_969),
.Y(n_1333)
);

CKINVDCx16_ASAP7_75t_R g1334 ( 
.A(n_1059),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_915),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_1093),
.Y(n_1336)
);

NOR2xp67_ASAP7_75t_L g1337 ( 
.A(n_1088),
.B(n_469),
.Y(n_1337)
);

CKINVDCx16_ASAP7_75t_R g1338 ( 
.A(n_784),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_916),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_898),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_916),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_917),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_917),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_899),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_924),
.Y(n_1345)
);

NOR2xp67_ASAP7_75t_L g1346 ( 
.A(n_1100),
.B(n_482),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_924),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_900),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_901),
.Y(n_1349)
);

CKINVDCx16_ASAP7_75t_R g1350 ( 
.A(n_784),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_908),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1054),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_930),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_930),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_935),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_935),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_936),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_910),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_913),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_919),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_936),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_938),
.Y(n_1362)
);

INVxp67_ASAP7_75t_SL g1363 ( 
.A(n_812),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_938),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_947),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_921),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_922),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_947),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_923),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_926),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_952),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_928),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1063),
.B(n_492),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_952),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_931),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1102),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_953),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_953),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_954),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_939),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_954),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_940),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_941),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_813),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_942),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_957),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_957),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_943),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_944),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_948),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_949),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_951),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1102),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_955),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_958),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_956),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_959),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_958),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_967),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_967),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_960),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_965),
.Y(n_1402)
);

XNOR2x1_ASAP7_75t_L g1403 ( 
.A(n_801),
.B(n_724),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_987),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_966),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_987),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1053),
.B(n_499),
.Y(n_1407)
);

BUFx2_ASAP7_75t_SL g1408 ( 
.A(n_843),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_968),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_989),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_989),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_812),
.B(n_733),
.Y(n_1412)
);

NOR2xp67_ASAP7_75t_L g1413 ( 
.A(n_1002),
.B(n_504),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1002),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_765),
.B(n_752),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1012),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1012),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_971),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_972),
.Y(n_1419)
);

CKINVDCx16_ASAP7_75t_R g1420 ( 
.A(n_896),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_973),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1013),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1013),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_974),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_976),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_977),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_978),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_1020),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1020),
.Y(n_1429)
);

INVxp33_ASAP7_75t_L g1430 ( 
.A(n_918),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_979),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1025),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1032),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1025),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1204),
.B(n_946),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1129),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1263),
.B(n_850),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1309),
.B(n_1323),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1129),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1132),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1373),
.B(n_1253),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1154),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1430),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1158),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1133),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1363),
.B(n_1412),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1156),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1158),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1193),
.A2(n_1039),
.B1(n_1041),
.B2(n_1038),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1211),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1269),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1185),
.B(n_850),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1219),
.A2(n_1038),
.B1(n_1041),
.B2(n_1039),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1269),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1280),
.B(n_946),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1319),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1166),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1167),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1319),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1352),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1211),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1352),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1138),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1164),
.B(n_1049),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1136),
.B(n_1049),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1376),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1146),
.B(n_1052),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1324),
.B(n_946),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1412),
.B(n_856),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1376),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1169),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1236),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1176),
.B(n_946),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1412),
.B(n_856),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1177),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1181),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1236),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1161),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1230),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1183),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1172),
.B(n_907),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1187),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1170),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1219),
.A2(n_1052),
.B1(n_1056),
.B2(n_1055),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1188),
.Y(n_1485)
);

BUFx8_ASAP7_75t_SL g1486 ( 
.A(n_1171),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1189),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1317),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1170),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1190),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1149),
.B(n_1055),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1191),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1196),
.Y(n_1493)
);

CKINVDCx6p67_ASAP7_75t_R g1494 ( 
.A(n_1194),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1150),
.B(n_946),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1200),
.Y(n_1496)
);

NOR2x1_ASAP7_75t_L g1497 ( 
.A(n_1212),
.B(n_907),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1170),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1408),
.A2(n_1060),
.B1(n_1062),
.B2(n_1056),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1317),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1407),
.B(n_946),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_SL g1502 ( 
.A1(n_1223),
.A2(n_1060),
.B1(n_1064),
.B2(n_1062),
.Y(n_1502)
);

XNOR2xp5_ASAP7_75t_L g1503 ( 
.A(n_1403),
.B(n_1064),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1135),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1202),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1384),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1384),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1170),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1206),
.B(n_925),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1393),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1208),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1218),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1182),
.B(n_925),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1170),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1221),
.B(n_933),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1222),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1393),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1393),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1225),
.B(n_933),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1433),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1228),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1229),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1332),
.B(n_1137),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1231),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1232),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1237),
.B(n_1058),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1168),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1240),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1243),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1248),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1249),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_L g1532 ( 
.A(n_1192),
.B(n_946),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1252),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1197),
.B(n_1215),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1254),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1260),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1209),
.A2(n_801),
.B1(n_1035),
.B2(n_868),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1262),
.A2(n_1030),
.B(n_1026),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1266),
.B(n_1058),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1160),
.A2(n_1076),
.B1(n_1081),
.B2(n_1070),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1268),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1271),
.B(n_1079),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1272),
.A2(n_1034),
.B(n_1031),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1276),
.Y(n_1544)
);

NAND2xp33_ASAP7_75t_L g1545 ( 
.A(n_1192),
.B(n_946),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1279),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1223),
.A2(n_1070),
.B1(n_1081),
.B2(n_1076),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1281),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1239),
.A2(n_1257),
.B1(n_1259),
.B2(n_1250),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1284),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1267),
.B(n_1003),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1295),
.B(n_1003),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1420),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1285),
.Y(n_1554)
);

AOI22x1_ASAP7_75t_SL g1555 ( 
.A1(n_1239),
.A2(n_644),
.B1(n_645),
.B2(n_639),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1287),
.Y(n_1556)
);

INVx6_ASAP7_75t_L g1557 ( 
.A(n_1283),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1288),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1329),
.B(n_1003),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1290),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1291),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1292),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1235),
.A2(n_1094),
.B1(n_1096),
.B2(n_1083),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1294),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1296),
.B(n_1079),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1297),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1298),
.B(n_1087),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1302),
.B(n_1087),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1304),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1305),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1307),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1320),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1327),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1328),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1340),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1330),
.B(n_1003),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1230),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1344),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1348),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1349),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1338),
.Y(n_1581)
);

BUFx8_ASAP7_75t_L g1582 ( 
.A(n_1242),
.Y(n_1582)
);

BUFx8_ASAP7_75t_L g1583 ( 
.A(n_1357),
.Y(n_1583)
);

AND2x6_ASAP7_75t_L g1584 ( 
.A(n_1351),
.B(n_1032),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1337),
.B(n_1003),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1346),
.B(n_1003),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1358),
.B(n_896),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1359),
.B(n_806),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1360),
.B(n_849),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1366),
.B(n_863),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1367),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1140),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1369),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1413),
.B(n_1003),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1370),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1372),
.B(n_1375),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1162),
.B(n_1003),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1350),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1380),
.B(n_857),
.Y(n_1599)
);

AND2x2_ASAP7_75t_SL g1600 ( 
.A(n_1334),
.B(n_1035),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1382),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1383),
.B(n_904),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1385),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1388),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1389),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1390),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1391),
.B(n_1083),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1392),
.B(n_897),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1394),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1250),
.A2(n_1096),
.B1(n_1097),
.B2(n_1094),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1396),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1397),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1401),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1234),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1402),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1405),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1409),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1418),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1257),
.A2(n_1108),
.B1(n_1110),
.B2(n_1097),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1259),
.A2(n_1110),
.B1(n_1112),
.B2(n_1108),
.Y(n_1620)
);

CKINVDCx6p67_ASAP7_75t_R g1621 ( 
.A(n_1336),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1419),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1421),
.B(n_905),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_L g1624 ( 
.A(n_1198),
.B(n_1115),
.C(n_1112),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1424),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1425),
.Y(n_1626)
);

INVx6_ASAP7_75t_L g1627 ( 
.A(n_1415),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1426),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1427),
.Y(n_1629)
);

XNOR2xp5_ASAP7_75t_L g1630 ( 
.A(n_1403),
.B(n_1115),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1431),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1220),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1220),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1134),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1205),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1207),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1220),
.Y(n_1637)
);

INVx5_ASAP7_75t_L g1638 ( 
.A(n_1145),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1139),
.Y(n_1639)
);

INVx5_ASAP7_75t_L g1640 ( 
.A(n_1255),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1275),
.A2(n_1111),
.B1(n_1015),
.B2(n_964),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1277),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1255),
.A2(n_647),
.B1(n_648),
.B2(n_646),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1289),
.A2(n_1300),
.B1(n_1316),
.B2(n_1310),
.Y(n_1644)
);

AND2x6_ASAP7_75t_L g1645 ( 
.A(n_1345),
.B(n_1067),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1321),
.A2(n_932),
.B1(n_970),
.B2(n_897),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1339),
.B(n_932),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1308),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1210),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1313),
.B(n_1027),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1361),
.B(n_970),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1224),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1313),
.B(n_1027),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1311),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1303),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1147),
.Y(n_1656)
);

OA21x2_ASAP7_75t_L g1657 ( 
.A1(n_1198),
.A2(n_1042),
.B(n_1037),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1335),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1374),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1301),
.B(n_1043),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1226),
.Y(n_1661)
);

INVx5_ASAP7_75t_L g1662 ( 
.A(n_1227),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1148),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1422),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1199),
.B(n_1027),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1233),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1244),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1245),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1199),
.B(n_1044),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1246),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1247),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1256),
.B(n_1027),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1256),
.B(n_1046),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1258),
.A2(n_653),
.B1(n_654),
.B2(n_652),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1151),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1264),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1258),
.B(n_1027),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1282),
.B(n_1027),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1265),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1274),
.Y(n_1680)
);

BUFx8_ASAP7_75t_L g1681 ( 
.A(n_1251),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1278),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1299),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1306),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1314),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1343),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1341),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1343),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1342),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1353),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1153),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1282),
.A2(n_659),
.B1(n_665),
.B2(n_655),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1241),
.A2(n_1072),
.B(n_1067),
.Y(n_1693)
);

CKINVDCx6p67_ASAP7_75t_R g1694 ( 
.A(n_1326),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1354),
.Y(n_1695)
);

OA21x2_ASAP7_75t_L g1696 ( 
.A1(n_1398),
.A2(n_1048),
.B(n_1047),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1135),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1355),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1356),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1434),
.B(n_1027),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1398),
.B(n_1051),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1404),
.B(n_1061),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1365),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1368),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1378),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1404),
.B(n_1065),
.Y(n_1706)
);

INVx3_ASAP7_75t_L g1707 ( 
.A(n_1379),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1381),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1406),
.B(n_1072),
.Y(n_1709)
);

INVx6_ASAP7_75t_L g1710 ( 
.A(n_1386),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1387),
.B(n_1027),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1395),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1406),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1410),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1410),
.Y(n_1715)
);

BUFx8_ASAP7_75t_L g1716 ( 
.A(n_1326),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1411),
.B(n_1066),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1411),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1414),
.B(n_1092),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1414),
.B(n_1092),
.Y(n_1720)
);

XNOR2xp5_ASAP7_75t_L g1721 ( 
.A(n_1141),
.B(n_817),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1417),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1525),
.Y(n_1723)
);

CKINVDCx20_ASAP7_75t_R g1724 ( 
.A(n_1504),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1486),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1525),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1443),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1486),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1634),
.Y(n_1729)
);

CKINVDCx20_ASAP7_75t_R g1730 ( 
.A(n_1504),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1634),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1450),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1639),
.Y(n_1733)
);

CKINVDCx20_ASAP7_75t_R g1734 ( 
.A(n_1697),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1639),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_R g1736 ( 
.A(n_1656),
.B(n_1417),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1656),
.Y(n_1737)
);

OAI21x1_ASAP7_75t_L g1738 ( 
.A1(n_1693),
.A2(n_1086),
.B(n_1075),
.Y(n_1738)
);

NAND2xp33_ASAP7_75t_R g1739 ( 
.A(n_1663),
.B(n_1173),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1570),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1445),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1709),
.B(n_1423),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1663),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1570),
.Y(n_1744)
);

CKINVDCx20_ASAP7_75t_R g1745 ( 
.A(n_1697),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1445),
.Y(n_1746)
);

INVxp33_ASAP7_75t_L g1747 ( 
.A(n_1463),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1450),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1675),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1675),
.Y(n_1750)
);

BUFx3_ASAP7_75t_L g1751 ( 
.A(n_1638),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1478),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1503),
.A2(n_1142),
.B1(n_1143),
.B2(n_1141),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1478),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1494),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1494),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1571),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1581),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1581),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1621),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1621),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1571),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1583),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1461),
.Y(n_1764)
);

CKINVDCx20_ASAP7_75t_R g1765 ( 
.A(n_1583),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1439),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1583),
.Y(n_1767)
);

OAI22xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1627),
.A2(n_1537),
.B1(n_1641),
.B2(n_1713),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1591),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1598),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1598),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1716),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1527),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1591),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1553),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1469),
.B(n_1423),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_R g1777 ( 
.A(n_1638),
.B(n_1429),
.Y(n_1777)
);

CKINVDCx20_ASAP7_75t_R g1778 ( 
.A(n_1716),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1448),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1527),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_1652),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1652),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1461),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_1716),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1582),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1638),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1601),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1601),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1638),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1614),
.Y(n_1790)
);

CKINVDCx20_ASAP7_75t_R g1791 ( 
.A(n_1582),
.Y(n_1791)
);

BUFx10_ASAP7_75t_L g1792 ( 
.A(n_1557),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1605),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_1638),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1592),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1605),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1710),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1710),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1710),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1612),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1612),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1694),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1616),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1694),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1709),
.B(n_1429),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1616),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1614),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1582),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1629),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1472),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1681),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_1681),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1627),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1472),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1629),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1447),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1627),
.B(n_1432),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1681),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1441),
.B(n_1432),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1441),
.B(n_1464),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1457),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1660),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1635),
.Y(n_1823)
);

CKINVDCx20_ASAP7_75t_R g1824 ( 
.A(n_1557),
.Y(n_1824)
);

INVxp67_ASAP7_75t_L g1825 ( 
.A(n_1660),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1477),
.Y(n_1826)
);

CKINVDCx5p33_ASAP7_75t_R g1827 ( 
.A(n_1635),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1477),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_R g1829 ( 
.A(n_1661),
.B(n_1165),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1635),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1635),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_R g1832 ( 
.A(n_1661),
.B(n_1347),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1686),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1636),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1488),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_1557),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1636),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_R g1838 ( 
.A(n_1479),
.B(n_1174),
.Y(n_1838)
);

INVx3_ASAP7_75t_L g1839 ( 
.A(n_1448),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1714),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1488),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1714),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1714),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1464),
.B(n_1178),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_R g1845 ( 
.A(n_1661),
.B(n_1347),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1458),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1714),
.Y(n_1847)
);

NOR2xp67_ASAP7_75t_L g1848 ( 
.A(n_1640),
.B(n_1178),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1636),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1469),
.B(n_1179),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1709),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1500),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1636),
.Y(n_1853)
);

CKINVDCx16_ASAP7_75t_R g1854 ( 
.A(n_1549),
.Y(n_1854)
);

NOR2xp67_ASAP7_75t_L g1855 ( 
.A(n_1640),
.B(n_1179),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1471),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1475),
.Y(n_1857)
);

CKINVDCx20_ASAP7_75t_R g1858 ( 
.A(n_1691),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1448),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1649),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1688),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1476),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1649),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1480),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_R g1865 ( 
.A(n_1670),
.B(n_1362),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1640),
.B(n_1180),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1649),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1439),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1649),
.Y(n_1869)
);

CKINVDCx20_ASAP7_75t_R g1870 ( 
.A(n_1453),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1687),
.Y(n_1871)
);

BUFx2_ASAP7_75t_L g1872 ( 
.A(n_1577),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1500),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1687),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1482),
.Y(n_1875)
);

NOR2xp67_ASAP7_75t_L g1876 ( 
.A(n_1640),
.B(n_1180),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1485),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1687),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1487),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_R g1880 ( 
.A(n_1670),
.B(n_1362),
.Y(n_1880)
);

BUFx6f_ASAP7_75t_L g1881 ( 
.A(n_1439),
.Y(n_1881)
);

NOR2xp67_ASAP7_75t_L g1882 ( 
.A(n_1640),
.B(n_1186),
.Y(n_1882)
);

CKINVDCx20_ASAP7_75t_R g1883 ( 
.A(n_1484),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1687),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1689),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1689),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1439),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1490),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1689),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1506),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1444),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1492),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1506),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1507),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1666),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1701),
.Y(n_1896)
);

XOR2xp5_ASAP7_75t_L g1897 ( 
.A(n_1721),
.B(n_1142),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1701),
.Y(n_1898)
);

CKINVDCx16_ASAP7_75t_R g1899 ( 
.A(n_1502),
.Y(n_1899)
);

BUFx3_ASAP7_75t_L g1900 ( 
.A(n_1436),
.Y(n_1900)
);

NAND2xp33_ASAP7_75t_R g1901 ( 
.A(n_1670),
.B(n_1130),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1493),
.Y(n_1902)
);

CKINVDCx20_ASAP7_75t_R g1903 ( 
.A(n_1547),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_1721),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1689),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1610),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1698),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1698),
.Y(n_1908)
);

AND3x2_ASAP7_75t_L g1909 ( 
.A(n_1713),
.B(n_1333),
.C(n_1331),
.Y(n_1909)
);

NOR2xp67_ASAP7_75t_L g1910 ( 
.A(n_1662),
.B(n_1624),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1698),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1444),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_1619),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1496),
.Y(n_1914)
);

AND3x2_ASAP7_75t_L g1915 ( 
.A(n_1715),
.B(n_1333),
.C(n_1331),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1469),
.B(n_1186),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1698),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1507),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1703),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_R g1920 ( 
.A(n_1704),
.B(n_1364),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1703),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_1703),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1620),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1703),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1505),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1511),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1662),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1662),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1512),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1474),
.B(n_1130),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1662),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1662),
.Y(n_1932)
);

CKINVDCx20_ASAP7_75t_R g1933 ( 
.A(n_1503),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1630),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1630),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1516),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1704),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1704),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1521),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1522),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1528),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1707),
.Y(n_1942)
);

CKINVDCx20_ASAP7_75t_R g1943 ( 
.A(n_1563),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1510),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_1707),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1707),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1449),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1499),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1452),
.B(n_1092),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1530),
.Y(n_1950)
);

CKINVDCx20_ASAP7_75t_R g1951 ( 
.A(n_1540),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1600),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1474),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1600),
.Y(n_1954)
);

CKINVDCx20_ASAP7_75t_R g1955 ( 
.A(n_1644),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1555),
.Y(n_1956)
);

OR2x2_ASAP7_75t_SL g1957 ( 
.A(n_1715),
.B(n_1364),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1533),
.Y(n_1958)
);

BUFx10_ASAP7_75t_L g1959 ( 
.A(n_1647),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1452),
.B(n_1092),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1668),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1668),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_1676),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1676),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1679),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_1702),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1679),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1683),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1683),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1685),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1541),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1518),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1685),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1690),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1690),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1444),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1474),
.Y(n_1977)
);

CKINVDCx20_ASAP7_75t_R g1978 ( 
.A(n_1702),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1544),
.Y(n_1979)
);

BUFx3_ASAP7_75t_L g1980 ( 
.A(n_1436),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1706),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1437),
.B(n_1092),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_1706),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_1695),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_1717),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1695),
.Y(n_1986)
);

CKINVDCx5p33_ASAP7_75t_R g1987 ( 
.A(n_1699),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1546),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1444),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1548),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1666),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1550),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1669),
.B(n_1673),
.Y(n_1993)
);

CKINVDCx20_ASAP7_75t_R g1994 ( 
.A(n_1717),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1699),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1712),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1437),
.B(n_1092),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_1712),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1446),
.Y(n_1999)
);

HB1xp67_ASAP7_75t_L g2000 ( 
.A(n_1446),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1510),
.Y(n_2001)
);

CKINVDCx20_ASAP7_75t_R g2002 ( 
.A(n_1667),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1556),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1671),
.Y(n_2004)
);

CKINVDCx9p33_ASAP7_75t_R g2005 ( 
.A(n_1607),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1680),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1446),
.B(n_1131),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_R g2008 ( 
.A(n_1532),
.B(n_1371),
.Y(n_2008)
);

NAND2xp33_ASAP7_75t_SL g2009 ( 
.A(n_1669),
.B(n_1371),
.Y(n_2009)
);

BUFx10_ASAP7_75t_L g2010 ( 
.A(n_1647),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1517),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1682),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1558),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1673),
.B(n_1131),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1999),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1820),
.B(n_1658),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1751),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1732),
.Y(n_2018)
);

INVx3_ASAP7_75t_L g2019 ( 
.A(n_1751),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1898),
.B(n_1648),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2000),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1864),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1739),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1993),
.A2(n_1645),
.B1(n_1696),
.B2(n_1657),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1819),
.B(n_1844),
.Y(n_2025)
);

INVx5_ASAP7_75t_L g2026 ( 
.A(n_1766),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1981),
.A2(n_1645),
.B1(n_1696),
.B2(n_1657),
.Y(n_2027)
);

INVx4_ASAP7_75t_L g2028 ( 
.A(n_1792),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1840),
.B(n_1842),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1732),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1748),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1766),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1748),
.Y(n_2033)
);

BUFx4f_ASAP7_75t_L g2034 ( 
.A(n_1758),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1875),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1985),
.B(n_1648),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1896),
.B(n_1658),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1825),
.B(n_1437),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1764),
.Y(n_2039)
);

INVx4_ASAP7_75t_L g2040 ( 
.A(n_1792),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1817),
.B(n_1523),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1947),
.B(n_1659),
.Y(n_2042)
);

INVx3_ASAP7_75t_L g2043 ( 
.A(n_1766),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1877),
.Y(n_2044)
);

INVx5_ASAP7_75t_L g2045 ( 
.A(n_1766),
.Y(n_2045)
);

INVx6_ASAP7_75t_L g2046 ( 
.A(n_1792),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1879),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_1824),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1822),
.A2(n_1645),
.B1(n_1696),
.B2(n_1657),
.Y(n_2049)
);

HB1xp67_ASAP7_75t_L g2050 ( 
.A(n_1790),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_1951),
.A2(n_1645),
.B1(n_1596),
.B2(n_1529),
.Y(n_2051)
);

INVx5_ASAP7_75t_L g2052 ( 
.A(n_1766),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1888),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1807),
.B(n_1238),
.Y(n_2054)
);

INVx5_ASAP7_75t_L g2055 ( 
.A(n_1868),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1840),
.B(n_1842),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_1795),
.Y(n_2057)
);

INVx2_ASAP7_75t_SL g2058 ( 
.A(n_1752),
.Y(n_2058)
);

INVx5_ASAP7_75t_L g2059 ( 
.A(n_1868),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1752),
.B(n_1318),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1892),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1851),
.B(n_1523),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1977),
.B(n_1523),
.Y(n_2063)
);

INVx4_ASAP7_75t_L g2064 ( 
.A(n_1797),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1764),
.Y(n_2065)
);

INVx2_ASAP7_75t_SL g2066 ( 
.A(n_1754),
.Y(n_2066)
);

AND2x4_ASAP7_75t_L g2067 ( 
.A(n_1977),
.B(n_1633),
.Y(n_2067)
);

NAND3xp33_ASAP7_75t_L g2068 ( 
.A(n_1754),
.B(n_1159),
.C(n_1718),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1783),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1902),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1783),
.Y(n_2071)
);

INVx5_ASAP7_75t_L g2072 ( 
.A(n_1868),
.Y(n_2072)
);

CKINVDCx20_ASAP7_75t_R g2073 ( 
.A(n_1836),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1810),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_1961),
.B(n_1962),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1914),
.Y(n_2076)
);

BUFx6f_ASAP7_75t_L g2077 ( 
.A(n_1868),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1925),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_1816),
.A2(n_1645),
.B1(n_1596),
.B2(n_1529),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1843),
.B(n_1650),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_1736),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_1813),
.B(n_1633),
.Y(n_2082)
);

INVxp33_ASAP7_75t_SL g2083 ( 
.A(n_1798),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1729),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1821),
.A2(n_1645),
.B1(n_1596),
.B2(n_1529),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1868),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1881),
.Y(n_2087)
);

OR2x2_ASAP7_75t_L g2088 ( 
.A(n_1741),
.B(n_1654),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1926),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_1746),
.B(n_1654),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1810),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1729),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1929),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1814),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1799),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1936),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2007),
.B(n_1647),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1939),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1731),
.Y(n_2099)
);

NAND2x1p5_ASAP7_75t_L g2100 ( 
.A(n_1900),
.B(n_1524),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1940),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_1759),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1941),
.B(n_1440),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_1961),
.B(n_1659),
.Y(n_2104)
);

INVx4_ASAP7_75t_L g2105 ( 
.A(n_1823),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2007),
.B(n_1651),
.Y(n_2106)
);

INVx4_ASAP7_75t_L g2107 ( 
.A(n_1827),
.Y(n_2107)
);

NOR2x1p5_ASAP7_75t_L g2108 ( 
.A(n_1731),
.B(n_1159),
.Y(n_2108)
);

AND2x4_ASAP7_75t_L g2109 ( 
.A(n_1953),
.B(n_1526),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1950),
.Y(n_2110)
);

CKINVDCx11_ASAP7_75t_R g2111 ( 
.A(n_1724),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_1770),
.B(n_1651),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1814),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_1846),
.A2(n_1529),
.B1(n_1566),
.B2(n_1536),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1958),
.Y(n_2115)
);

INVx1_ASAP7_75t_SL g2116 ( 
.A(n_1872),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1826),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1930),
.B(n_1651),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_1962),
.B(n_1963),
.Y(n_2119)
);

INVx3_ASAP7_75t_L g2120 ( 
.A(n_1881),
.Y(n_2120)
);

NOR2x1p5_ASAP7_75t_L g2121 ( 
.A(n_1733),
.B(n_1722),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1971),
.B(n_1442),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_1856),
.A2(n_1566),
.B1(n_1569),
.B2(n_1536),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1979),
.B(n_1607),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1843),
.B(n_1653),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1988),
.B(n_1438),
.Y(n_2126)
);

INVx1_ASAP7_75t_SL g2127 ( 
.A(n_1730),
.Y(n_2127)
);

BUFx8_ASAP7_75t_SL g2128 ( 
.A(n_1728),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1847),
.B(n_1719),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1930),
.B(n_1776),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_1963),
.B(n_1465),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1847),
.B(n_1720),
.Y(n_2132)
);

BUFx8_ASAP7_75t_SL g2133 ( 
.A(n_1728),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1990),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1881),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1992),
.Y(n_2136)
);

INVx2_ASAP7_75t_SL g2137 ( 
.A(n_1770),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1857),
.A2(n_1566),
.B1(n_1569),
.B2(n_1536),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1826),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1828),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1881),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2003),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2013),
.B(n_1465),
.Y(n_2143)
);

OAI22xp33_ASAP7_75t_L g2144 ( 
.A1(n_1948),
.A2(n_1535),
.B1(n_1554),
.B2(n_1524),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1881),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1964),
.B(n_1665),
.Y(n_2146)
);

AND2x2_ASAP7_75t_SL g2147 ( 
.A(n_1899),
.B(n_1532),
.Y(n_2147)
);

NOR2xp33_ASAP7_75t_L g2148 ( 
.A(n_1964),
.B(n_1467),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1862),
.B(n_1467),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1965),
.B(n_1491),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1723),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_1952),
.A2(n_1566),
.B1(n_1569),
.B2(n_1536),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1965),
.B(n_1491),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1726),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_1771),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1740),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1744),
.Y(n_2157)
);

INVx1_ASAP7_75t_SL g2158 ( 
.A(n_1734),
.Y(n_2158)
);

OAI22xp33_ASAP7_75t_SL g2159 ( 
.A1(n_1967),
.A2(n_1646),
.B1(n_1684),
.B2(n_1705),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_1967),
.B(n_1672),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1968),
.B(n_1524),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1757),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1828),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1968),
.B(n_1677),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1762),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_1727),
.Y(n_2166)
);

BUFx4f_ASAP7_75t_L g2167 ( 
.A(n_1776),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1835),
.Y(n_2168)
);

NAND2xp33_ASAP7_75t_SL g2169 ( 
.A(n_1777),
.B(n_1708),
.Y(n_2169)
);

INVx3_ASAP7_75t_L g2170 ( 
.A(n_1887),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_1887),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1969),
.B(n_1678),
.Y(n_2172)
);

OAI22xp33_ASAP7_75t_SL g2173 ( 
.A1(n_1969),
.A2(n_1642),
.B1(n_1664),
.B2(n_1655),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_1850),
.B(n_1588),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1835),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_1887),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_SL g2177 ( 
.A(n_1970),
.B(n_1700),
.Y(n_2177)
);

INVxp67_ASAP7_75t_SL g2178 ( 
.A(n_1887),
.Y(n_2178)
);

INVx6_ASAP7_75t_L g2179 ( 
.A(n_1959),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_L g2180 ( 
.A1(n_1952),
.A2(n_1603),
.B1(n_1613),
.B2(n_1569),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_1771),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_1970),
.B(n_1481),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_L g2183 ( 
.A(n_1973),
.B(n_1481),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1887),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_1973),
.A2(n_1513),
.B1(n_1481),
.B2(n_1545),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1841),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1841),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1974),
.B(n_1535),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_1974),
.B(n_1535),
.Y(n_2189)
);

BUFx10_ASAP7_75t_L g2190 ( 
.A(n_1733),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1769),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_SL g2192 ( 
.A(n_1975),
.B(n_1711),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1774),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1975),
.B(n_1554),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1787),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_1984),
.B(n_1513),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1788),
.Y(n_2197)
);

BUFx3_ASAP7_75t_L g2198 ( 
.A(n_1773),
.Y(n_2198)
);

INVx4_ASAP7_75t_L g2199 ( 
.A(n_1830),
.Y(n_2199)
);

AO22x2_ASAP7_75t_L g2200 ( 
.A1(n_1897),
.A2(n_1637),
.B1(n_1632),
.B2(n_1599),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1793),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1984),
.B(n_1554),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1796),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1800),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1801),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_1775),
.B(n_1747),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1803),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1852),
.Y(n_2208)
);

AOI22xp33_ASAP7_75t_SL g2209 ( 
.A1(n_2008),
.A2(n_1270),
.B1(n_1273),
.B2(n_1261),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1806),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_L g2211 ( 
.A1(n_1954),
.A2(n_1613),
.B1(n_1615),
.B2(n_1603),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1809),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1735),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1986),
.B(n_1578),
.Y(n_2214)
);

INVx4_ASAP7_75t_L g2215 ( 
.A(n_1831),
.Y(n_2215)
);

INVx5_ASAP7_75t_L g2216 ( 
.A(n_1891),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1986),
.B(n_1513),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1987),
.B(n_1578),
.Y(n_2218)
);

BUFx2_ASAP7_75t_L g2219 ( 
.A(n_1745),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1987),
.B(n_1578),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1815),
.Y(n_2221)
);

BUFx8_ASAP7_75t_SL g2222 ( 
.A(n_1725),
.Y(n_2222)
);

OR2x6_ASAP7_75t_L g2223 ( 
.A(n_1753),
.B(n_1588),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1895),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_1995),
.B(n_1595),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1995),
.B(n_1455),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1991),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1735),
.Y(n_2228)
);

BUFx4f_ASAP7_75t_L g2229 ( 
.A(n_1850),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_1954),
.A2(n_1613),
.B1(n_1615),
.B2(n_1603),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1996),
.B(n_1595),
.Y(n_2231)
);

OR2x6_ASAP7_75t_L g2232 ( 
.A(n_1916),
.B(n_1588),
.Y(n_2232)
);

NAND2xp33_ASAP7_75t_L g2233 ( 
.A(n_1927),
.B(n_1473),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1852),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1891),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1944),
.Y(n_2236)
);

AND2x6_ASAP7_75t_L g2237 ( 
.A(n_1916),
.B(n_1589),
.Y(n_2237)
);

OR2x6_ASAP7_75t_L g2238 ( 
.A(n_1833),
.B(n_1589),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1944),
.Y(n_2239)
);

INVx4_ASAP7_75t_L g2240 ( 
.A(n_1834),
.Y(n_2240)
);

INVx5_ASAP7_75t_L g2241 ( 
.A(n_1891),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_1737),
.B(n_1589),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_1737),
.B(n_1590),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_1996),
.B(n_1595),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_1891),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_1959),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2001),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_1998),
.B(n_1468),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2001),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1998),
.B(n_1609),
.Y(n_2250)
);

NAND3xp33_ASAP7_75t_L g2251 ( 
.A(n_1743),
.B(n_1692),
.C(n_1545),
.Y(n_2251)
);

INVx2_ASAP7_75t_SL g2252 ( 
.A(n_1959),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2011),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1873),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2011),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1873),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2010),
.B(n_1501),
.Y(n_2257)
);

INVx3_ASAP7_75t_L g2258 ( 
.A(n_1891),
.Y(n_2258)
);

OAI21xp33_ASAP7_75t_SL g2259 ( 
.A1(n_1742),
.A2(n_1693),
.B(n_1611),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1890),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_1743),
.B(n_1590),
.Y(n_2261)
);

INVx3_ASAP7_75t_L g2262 ( 
.A(n_1912),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1937),
.B(n_1609),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_1938),
.B(n_1609),
.Y(n_2264)
);

BUFx2_ASAP7_75t_L g2265 ( 
.A(n_1966),
.Y(n_2265)
);

OR2x6_ASAP7_75t_L g2266 ( 
.A(n_1861),
.B(n_1805),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_2010),
.B(n_2014),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2010),
.B(n_1768),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1749),
.B(n_1590),
.Y(n_2269)
);

OAI22xp33_ASAP7_75t_SL g2270 ( 
.A1(n_1854),
.A2(n_1674),
.B1(n_1643),
.B2(n_1599),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1890),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_2004),
.B(n_1611),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_L g2273 ( 
.A(n_2004),
.B(n_1611),
.Y(n_2273)
);

INVx1_ASAP7_75t_SL g2274 ( 
.A(n_1858),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_1837),
.B(n_1617),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1893),
.Y(n_2276)
);

NAND2x1p5_ASAP7_75t_L g2277 ( 
.A(n_1900),
.B(n_1617),
.Y(n_2277)
);

INVxp67_ASAP7_75t_SL g2278 ( 
.A(n_1912),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_1849),
.B(n_1526),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1942),
.B(n_1617),
.Y(n_2280)
);

OR2x2_ASAP7_75t_L g2281 ( 
.A(n_1749),
.B(n_1587),
.Y(n_2281)
);

INVx1_ASAP7_75t_SL g2282 ( 
.A(n_1781),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1893),
.Y(n_2283)
);

AOI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_1901),
.A2(n_1399),
.B1(n_1400),
.B2(n_1377),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2006),
.A2(n_1399),
.B1(n_1400),
.B2(n_1377),
.Y(n_2285)
);

OR2x6_ASAP7_75t_L g2286 ( 
.A(n_1848),
.B(n_1526),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1912),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1894),
.Y(n_2288)
);

INVx4_ASAP7_75t_L g2289 ( 
.A(n_1853),
.Y(n_2289)
);

NAND2xp33_ASAP7_75t_L g2290 ( 
.A(n_1928),
.B(n_1534),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_SL g2291 ( 
.A(n_1761),
.Y(n_2291)
);

AND2x6_ASAP7_75t_L g2292 ( 
.A(n_1779),
.B(n_1623),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1894),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1945),
.B(n_1509),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_1860),
.B(n_1594),
.Y(n_2295)
);

INVx6_ASAP7_75t_L g2296 ( 
.A(n_1980),
.Y(n_2296)
);

INVx1_ASAP7_75t_SL g2297 ( 
.A(n_1782),
.Y(n_2297)
);

BUFx2_ASAP7_75t_L g2298 ( 
.A(n_1978),
.Y(n_2298)
);

INVx3_ASAP7_75t_L g2299 ( 
.A(n_1912),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1918),
.Y(n_2300)
);

NAND2xp33_ASAP7_75t_L g2301 ( 
.A(n_1931),
.B(n_1932),
.Y(n_2301)
);

NOR2xp33_ASAP7_75t_L g2302 ( 
.A(n_1863),
.B(n_1531),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1946),
.B(n_1509),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_1867),
.B(n_1531),
.Y(n_2304)
);

NOR2x1p5_ASAP7_75t_L g2305 ( 
.A(n_1750),
.B(n_1772),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_1869),
.B(n_1603),
.Y(n_2306)
);

INVx4_ASAP7_75t_SL g2307 ( 
.A(n_1912),
.Y(n_2307)
);

INVx3_ASAP7_75t_L g2308 ( 
.A(n_1976),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_1871),
.B(n_1874),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2025),
.B(n_1878),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2025),
.B(n_1884),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2016),
.B(n_1885),
.Y(n_2312)
);

O2A1O1Ixp33_ASAP7_75t_L g2313 ( 
.A1(n_2016),
.A2(n_1949),
.B(n_1960),
.C(n_1866),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2075),
.B(n_1886),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2075),
.B(n_1889),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2119),
.B(n_1905),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2131),
.B(n_1907),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2131),
.B(n_2148),
.Y(n_2318)
);

AOI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2148),
.A2(n_1943),
.B1(n_1994),
.B2(n_1983),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2022),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2042),
.B(n_1750),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2035),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_2032),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2044),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2047),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2150),
.B(n_1908),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2153),
.B(n_2272),
.Y(n_2327)
);

NAND2xp33_ASAP7_75t_L g2328 ( 
.A(n_2081),
.B(n_1780),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2272),
.B(n_1911),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2273),
.B(n_1917),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2053),
.Y(n_2331)
);

AND2x6_ASAP7_75t_L g2332 ( 
.A(n_2032),
.B(n_2077),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2018),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2018),
.Y(n_2334)
);

NAND2xp33_ASAP7_75t_L g2335 ( 
.A(n_2237),
.B(n_1829),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_2042),
.B(n_1955),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2119),
.B(n_1919),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2273),
.B(n_1921),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_SL g2339 ( 
.A(n_2023),
.B(n_1755),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2061),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2104),
.A2(n_2002),
.B1(n_1428),
.B2(n_1416),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2104),
.B(n_1922),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2070),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2281),
.B(n_2112),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2076),
.Y(n_2345)
);

BUFx6f_ASAP7_75t_L g2346 ( 
.A(n_2032),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2034),
.B(n_1924),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_L g2348 ( 
.A(n_2060),
.B(n_1416),
.Y(n_2348)
);

INVx1_ASAP7_75t_SL g2349 ( 
.A(n_2116),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2225),
.B(n_2012),
.Y(n_2350)
);

BUFx6f_ASAP7_75t_L g2351 ( 
.A(n_2032),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2225),
.B(n_1515),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_2034),
.B(n_1832),
.Y(n_2353)
);

AOI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_2182),
.A2(n_1428),
.B1(n_2009),
.B2(n_1883),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2244),
.B(n_1515),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2041),
.B(n_1957),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2244),
.B(n_1519),
.Y(n_2357)
);

INVx8_ASAP7_75t_L g2358 ( 
.A(n_2292),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2078),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_L g2360 ( 
.A1(n_2147),
.A2(n_1602),
.B1(n_1623),
.B2(n_1599),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2143),
.B(n_1519),
.Y(n_2361)
);

NOR2xp33_ASAP7_75t_L g2362 ( 
.A(n_2083),
.B(n_1261),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2091),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2149),
.B(n_1542),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2091),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2124),
.B(n_1542),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_SL g2367 ( 
.A(n_2269),
.B(n_1845),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2077),
.Y(n_2368)
);

INVx4_ASAP7_75t_L g2369 ( 
.A(n_2046),
.Y(n_2369)
);

INVx2_ASAP7_75t_SL g2370 ( 
.A(n_2095),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2020),
.B(n_1565),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2089),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2036),
.B(n_1565),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_2077),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2182),
.A2(n_1903),
.B1(n_1906),
.B2(n_1870),
.Y(n_2375)
);

CKINVDCx20_ASAP7_75t_R g2376 ( 
.A(n_2222),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2037),
.B(n_1567),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_2242),
.B(n_1865),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2037),
.B(n_1567),
.Y(n_2379)
);

AOI22xp33_ASAP7_75t_L g2380 ( 
.A1(n_2147),
.A2(n_1623),
.B1(n_1602),
.B2(n_1615),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2093),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2097),
.B(n_1539),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2140),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_2285),
.B(n_1270),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2106),
.B(n_1539),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2243),
.B(n_1880),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2279),
.B(n_2198),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2096),
.Y(n_2388)
);

INVx2_ASAP7_75t_SL g2389 ( 
.A(n_2095),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2038),
.B(n_1539),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2237),
.B(n_1568),
.Y(n_2391)
);

INVx2_ASAP7_75t_SL g2392 ( 
.A(n_2046),
.Y(n_2392)
);

A2O1A1Ixp33_ASAP7_75t_L g2393 ( 
.A1(n_2251),
.A2(n_1882),
.B(n_1876),
.C(n_1855),
.Y(n_2393)
);

INVx4_ASAP7_75t_L g2394 ( 
.A(n_2046),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2098),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2118),
.B(n_1587),
.Y(n_2396)
);

AND3x4_ASAP7_75t_L g2397 ( 
.A(n_2198),
.B(n_2279),
.C(n_2133),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2237),
.B(n_1568),
.Y(n_2398)
);

INVxp67_ASAP7_75t_SL g2399 ( 
.A(n_2178),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_2128),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_2261),
.B(n_1920),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2237),
.B(n_2126),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2167),
.B(n_1789),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_L g2404 ( 
.A1(n_2223),
.A2(n_1602),
.B1(n_1615),
.B2(n_1613),
.Y(n_2404)
);

INVx2_ASAP7_75t_SL g2405 ( 
.A(n_2048),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2101),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2237),
.B(n_1568),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2140),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2161),
.B(n_1608),
.Y(n_2409)
);

BUFx2_ASAP7_75t_L g2410 ( 
.A(n_2073),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2110),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2115),
.Y(n_2412)
);

AOI221xp5_ASAP7_75t_L g2413 ( 
.A1(n_2159),
.A2(n_1608),
.B1(n_1923),
.B2(n_1913),
.C(n_1562),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_L g2414 ( 
.A(n_2174),
.B(n_1755),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2188),
.B(n_1560),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_2077),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2189),
.B(n_1561),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2134),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2194),
.B(n_1564),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2202),
.B(n_1572),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2136),
.Y(n_2421)
);

NOR3xp33_ASAP7_75t_L g2422 ( 
.A(n_2068),
.B(n_1497),
.C(n_2005),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2232),
.B(n_2130),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2214),
.B(n_2218),
.Y(n_2424)
);

NAND2xp33_ASAP7_75t_L g2425 ( 
.A(n_2292),
.B(n_1786),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2220),
.B(n_2231),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_2167),
.B(n_2229),
.Y(n_2427)
);

AOI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_2183),
.A2(n_1838),
.B1(n_1772),
.B2(n_1760),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2232),
.B(n_1934),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2250),
.B(n_1573),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2302),
.B(n_1574),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2142),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2302),
.B(n_1575),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_SL g2434 ( 
.A(n_2229),
.B(n_1794),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2183),
.B(n_1756),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2304),
.B(n_1579),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_SL g2437 ( 
.A(n_2196),
.B(n_1756),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_2086),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2304),
.B(n_1580),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2234),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2196),
.B(n_1593),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2217),
.B(n_1604),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2217),
.B(n_1606),
.Y(n_2443)
);

NOR3xp33_ASAP7_75t_L g2444 ( 
.A(n_2270),
.B(n_1016),
.C(n_1618),
.Y(n_2444)
);

INVx3_ASAP7_75t_L g2445 ( 
.A(n_2026),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2232),
.B(n_1935),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2058),
.B(n_1760),
.Y(n_2447)
);

NAND2xp33_ASAP7_75t_L g2448 ( 
.A(n_2292),
.B(n_1779),
.Y(n_2448)
);

BUFx6f_ASAP7_75t_L g2449 ( 
.A(n_2086),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2275),
.B(n_1625),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2234),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2275),
.B(n_1626),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_L g2453 ( 
.A(n_2166),
.B(n_1982),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2030),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2284),
.B(n_1273),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2151),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2306),
.B(n_1628),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2306),
.B(n_1622),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2031),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2062),
.B(n_1622),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2103),
.B(n_1622),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_SL g2462 ( 
.A(n_2190),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2122),
.B(n_1622),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2294),
.B(n_1631),
.Y(n_2464)
);

NOR3xp33_ASAP7_75t_L g2465 ( 
.A(n_2066),
.B(n_1910),
.C(n_1585),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2154),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2303),
.B(n_1631),
.Y(n_2467)
);

BUFx6f_ASAP7_75t_L g2468 ( 
.A(n_2086),
.Y(n_2468)
);

AOI22xp33_ASAP7_75t_L g2469 ( 
.A1(n_2223),
.A2(n_1631),
.B1(n_1520),
.B2(n_1918),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2156),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2224),
.B(n_1631),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2033),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2227),
.B(n_1997),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2039),
.Y(n_2474)
);

INVx2_ASAP7_75t_SL g2475 ( 
.A(n_2190),
.Y(n_2475)
);

INVx2_ASAP7_75t_SL g2476 ( 
.A(n_2084),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_2185),
.B(n_1763),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_SL g2478 ( 
.A(n_2137),
.B(n_2155),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2166),
.B(n_2050),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2157),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2088),
.B(n_1980),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2050),
.B(n_1802),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2090),
.B(n_1779),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2181),
.B(n_1763),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_SL g2485 ( 
.A(n_2282),
.B(n_1767),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_2238),
.B(n_1804),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_SL g2487 ( 
.A(n_2297),
.B(n_1767),
.Y(n_2487)
);

AOI22xp33_ASAP7_75t_L g2488 ( 
.A1(n_2223),
.A2(n_2051),
.B1(n_2027),
.B2(n_2049),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2065),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2015),
.B(n_1839),
.Y(n_2490)
);

INVxp67_ASAP7_75t_L g2491 ( 
.A(n_2206),
.Y(n_2491)
);

INVxp67_ASAP7_75t_L g2492 ( 
.A(n_2054),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2021),
.B(n_1839),
.Y(n_2493)
);

OR2x2_ASAP7_75t_L g2494 ( 
.A(n_2102),
.B(n_1808),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2162),
.Y(n_2495)
);

INVx2_ASAP7_75t_SL g2496 ( 
.A(n_2092),
.Y(n_2496)
);

NAND2xp33_ASAP7_75t_L g2497 ( 
.A(n_2292),
.B(n_1839),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2292),
.B(n_1909),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2109),
.B(n_1915),
.Y(n_2499)
);

AND2x2_ASAP7_75t_L g2500 ( 
.A(n_2238),
.B(n_1143),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2109),
.B(n_1972),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_SL g2502 ( 
.A(n_2105),
.B(n_1811),
.Y(n_2502)
);

NOR2xp67_ASAP7_75t_L g2503 ( 
.A(n_2057),
.B(n_1818),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2238),
.B(n_1286),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2144),
.B(n_1972),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2144),
.B(n_1972),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2029),
.B(n_1859),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2029),
.B(n_1286),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_L g2509 ( 
.A(n_2268),
.B(n_1293),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2069),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2071),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2056),
.B(n_1293),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2056),
.B(n_1312),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2082),
.B(n_1312),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2074),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2094),
.Y(n_2516)
);

OAI22xp5_ASAP7_75t_L g2517 ( 
.A1(n_2263),
.A2(n_1989),
.B1(n_1976),
.B2(n_1597),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2082),
.B(n_1315),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2165),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2267),
.B(n_2264),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_SL g2521 ( 
.A(n_2105),
.B(n_1976),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2267),
.B(n_2280),
.Y(n_2522)
);

NOR2xp33_ASAP7_75t_L g2523 ( 
.A(n_2127),
.B(n_1315),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2191),
.Y(n_2524)
);

NOR2xp67_ASAP7_75t_L g2525 ( 
.A(n_2107),
.B(n_2199),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2193),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2107),
.B(n_2199),
.Y(n_2527)
);

NOR2xp33_ASAP7_75t_L g2528 ( 
.A(n_2268),
.B(n_1322),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2215),
.B(n_1976),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2067),
.B(n_1322),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_2215),
.B(n_1976),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2113),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2067),
.B(n_1325),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2158),
.B(n_1325),
.Y(n_2534)
);

BUFx5_ASAP7_75t_L g2535 ( 
.A(n_2256),
.Y(n_2535)
);

BUFx3_ASAP7_75t_L g2536 ( 
.A(n_2111),
.Y(n_2536)
);

NAND2xp33_ASAP7_75t_L g2537 ( 
.A(n_2099),
.B(n_1989),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2246),
.B(n_1520),
.Y(n_2538)
);

NAND2xp33_ASAP7_75t_L g2539 ( 
.A(n_2213),
.B(n_1989),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2063),
.B(n_1435),
.Y(n_2540)
);

INVxp67_ASAP7_75t_SL g2541 ( 
.A(n_2178),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2209),
.B(n_1144),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_2240),
.B(n_1989),
.Y(n_2543)
);

INVx5_ASAP7_75t_L g2544 ( 
.A(n_2086),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_SL g2545 ( 
.A(n_2064),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_2240),
.B(n_1989),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2128),
.Y(n_2547)
);

OAI22xp5_ASAP7_75t_L g2548 ( 
.A1(n_2079),
.A2(n_1597),
.B1(n_1551),
.B2(n_1559),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2252),
.B(n_1520),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_2289),
.B(n_1778),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2195),
.Y(n_2551)
);

NAND2x1p5_ASAP7_75t_L g2552 ( 
.A(n_2369),
.B(n_2289),
.Y(n_2552)
);

AO22x2_ASAP7_75t_L g2553 ( 
.A1(n_2542),
.A2(n_2201),
.B1(n_2203),
.B2(n_2197),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2350),
.B(n_2209),
.Y(n_2554)
);

OR2x2_ASAP7_75t_L g2555 ( 
.A(n_2492),
.B(n_2274),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_L g2556 ( 
.A(n_2318),
.B(n_2228),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2387),
.B(n_2305),
.Y(n_2557)
);

AND2x4_ASAP7_75t_L g2558 ( 
.A(n_2387),
.B(n_2064),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2320),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2327),
.B(n_2309),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2349),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2322),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2310),
.B(n_2173),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_2311),
.B(n_1144),
.Y(n_2564)
);

AO22x2_ASAP7_75t_L g2565 ( 
.A1(n_2444),
.A2(n_2399),
.B1(n_2541),
.B2(n_2500),
.Y(n_2565)
);

AO22x2_ASAP7_75t_L g2566 ( 
.A1(n_2444),
.A2(n_2205),
.B1(n_2207),
.B2(n_2204),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2454),
.Y(n_2567)
);

AO22x2_ASAP7_75t_L g2568 ( 
.A1(n_2399),
.A2(n_2212),
.B1(n_2221),
.B2(n_2210),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2324),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2325),
.Y(n_2570)
);

AO22x2_ASAP7_75t_L g2571 ( 
.A1(n_2541),
.A2(n_2248),
.B1(n_2226),
.B2(n_2160),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2331),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2321),
.B(n_2265),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2340),
.Y(n_2574)
);

NAND2xp33_ASAP7_75t_L g2575 ( 
.A(n_2329),
.B(n_2169),
.Y(n_2575)
);

INVxp67_ASAP7_75t_L g2576 ( 
.A(n_2479),
.Y(n_2576)
);

AO22x2_ASAP7_75t_L g2577 ( 
.A1(n_2514),
.A2(n_2248),
.B1(n_2226),
.B2(n_2160),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2343),
.Y(n_2578)
);

NAND2x1p5_ASAP7_75t_L g2579 ( 
.A(n_2369),
.B(n_2394),
.Y(n_2579)
);

AO22x2_ASAP7_75t_L g2580 ( 
.A1(n_2518),
.A2(n_2164),
.B1(n_2172),
.B2(n_2146),
.Y(n_2580)
);

AO22x2_ASAP7_75t_L g2581 ( 
.A1(n_2488),
.A2(n_2164),
.B1(n_2172),
.B2(n_2146),
.Y(n_2581)
);

AO22x2_ASAP7_75t_L g2582 ( 
.A1(n_2488),
.A2(n_2192),
.B1(n_2177),
.B2(n_2200),
.Y(n_2582)
);

INVx2_ASAP7_75t_SL g2583 ( 
.A(n_2397),
.Y(n_2583)
);

OAI221xp5_ASAP7_75t_L g2584 ( 
.A1(n_2341),
.A2(n_2266),
.B1(n_2169),
.B2(n_2298),
.C(n_2219),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2345),
.Y(n_2585)
);

OAI221xp5_ASAP7_75t_L g2586 ( 
.A1(n_2413),
.A2(n_2266),
.B1(n_2309),
.B2(n_2051),
.C(n_2085),
.Y(n_2586)
);

AO22x2_ASAP7_75t_L g2587 ( 
.A1(n_2402),
.A2(n_2192),
.B1(n_2177),
.B2(n_2200),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2359),
.Y(n_2588)
);

OAI221xp5_ASAP7_75t_L g2589 ( 
.A1(n_2348),
.A2(n_2266),
.B1(n_2085),
.B2(n_2079),
.C(n_2180),
.Y(n_2589)
);

INVxp67_ASAP7_75t_L g2590 ( 
.A(n_2479),
.Y(n_2590)
);

AO22x2_ASAP7_75t_L g2591 ( 
.A1(n_2508),
.A2(n_2200),
.B1(n_2293),
.B2(n_2288),
.Y(n_2591)
);

HB1xp67_ASAP7_75t_L g2592 ( 
.A(n_2491),
.Y(n_2592)
);

AOI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2336),
.A2(n_1155),
.B1(n_1157),
.B2(n_1152),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2336),
.B(n_2121),
.Y(n_2594)
);

BUFx8_ASAP7_75t_L g2595 ( 
.A(n_2462),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2459),
.Y(n_2596)
);

AOI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2384),
.A2(n_1155),
.B1(n_1157),
.B2(n_1152),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2372),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2344),
.A2(n_1175),
.B1(n_1184),
.B2(n_1163),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2396),
.B(n_2108),
.Y(n_2600)
);

OAI221xp5_ASAP7_75t_L g2601 ( 
.A1(n_2354),
.A2(n_2211),
.B1(n_2230),
.B2(n_2180),
.C(n_2152),
.Y(n_2601)
);

AOI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2344),
.A2(n_1175),
.B1(n_1184),
.B2(n_1163),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2312),
.B(n_2028),
.Y(n_2603)
);

AOI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2455),
.A2(n_1201),
.B1(n_1203),
.B2(n_1195),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2317),
.B(n_1195),
.Y(n_2605)
);

INVxp67_ASAP7_75t_L g2606 ( 
.A(n_2482),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2381),
.Y(n_2607)
);

NAND2x1p5_ASAP7_75t_L g2608 ( 
.A(n_2394),
.B(n_2028),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2472),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2474),
.Y(n_2610)
);

CKINVDCx16_ASAP7_75t_R g2611 ( 
.A(n_2376),
.Y(n_2611)
);

NAND2x1p5_ASAP7_75t_L g2612 ( 
.A(n_2427),
.B(n_2040),
.Y(n_2612)
);

AND2x2_ASAP7_75t_SL g2613 ( 
.A(n_2335),
.B(n_2027),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_2400),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2547),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2388),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2395),
.Y(n_2617)
);

AO22x2_ASAP7_75t_L g2618 ( 
.A1(n_2512),
.A2(n_2300),
.B1(n_2239),
.B2(n_2247),
.Y(n_2618)
);

NAND2x1p5_ASAP7_75t_L g2619 ( 
.A(n_2370),
.B(n_2040),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2406),
.Y(n_2620)
);

OAI221xp5_ASAP7_75t_L g2621 ( 
.A1(n_2319),
.A2(n_2230),
.B1(n_2211),
.B2(n_2152),
.C(n_1074),
.Y(n_2621)
);

OAI221xp5_ASAP7_75t_L g2622 ( 
.A1(n_2509),
.A2(n_1080),
.B1(n_1082),
.B2(n_1073),
.C(n_1071),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2409),
.B(n_2296),
.Y(n_2623)
);

NAND2x1p5_ASAP7_75t_L g2624 ( 
.A(n_2389),
.B(n_2347),
.Y(n_2624)
);

AO22x2_ASAP7_75t_L g2625 ( 
.A1(n_2513),
.A2(n_2249),
.B1(n_2253),
.B2(n_2236),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2489),
.Y(n_2626)
);

AO22x2_ASAP7_75t_L g2627 ( 
.A1(n_2530),
.A2(n_2255),
.B1(n_2295),
.B2(n_2125),
.Y(n_2627)
);

AOI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2362),
.A2(n_1203),
.B1(n_1213),
.B2(n_1201),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2411),
.Y(n_2629)
);

OAI221xp5_ASAP7_75t_L g2630 ( 
.A1(n_2509),
.A2(n_1089),
.B1(n_1090),
.B2(n_1085),
.C(n_1084),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2412),
.Y(n_2631)
);

OR2x6_ASAP7_75t_L g2632 ( 
.A(n_2358),
.B(n_2179),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2418),
.Y(n_2633)
);

NAND2x1p5_ASAP7_75t_L g2634 ( 
.A(n_2410),
.B(n_2026),
.Y(n_2634)
);

AND2x2_ASAP7_75t_SL g2635 ( 
.A(n_2528),
.B(n_2404),
.Y(n_2635)
);

NOR2x1p5_ASAP7_75t_L g2636 ( 
.A(n_2536),
.B(n_2494),
.Y(n_2636)
);

AO22x2_ASAP7_75t_L g2637 ( 
.A1(n_2533),
.A2(n_2295),
.B1(n_2125),
.B2(n_2080),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2421),
.Y(n_2638)
);

INVxp67_ASAP7_75t_L g2639 ( 
.A(n_2482),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2432),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2492),
.B(n_2296),
.Y(n_2641)
);

OR2x2_ASAP7_75t_L g2642 ( 
.A(n_2491),
.B(n_767),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2510),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2361),
.B(n_2296),
.Y(n_2644)
);

AO22x2_ASAP7_75t_L g2645 ( 
.A1(n_2477),
.A2(n_2080),
.B1(n_2132),
.B2(n_2129),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2456),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2511),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2364),
.B(n_1933),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2515),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2466),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2470),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2480),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2495),
.Y(n_2653)
);

AND2x4_ASAP7_75t_L g2654 ( 
.A(n_2525),
.B(n_1812),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2519),
.Y(n_2655)
);

AND2x2_ASAP7_75t_SL g2656 ( 
.A(n_2528),
.B(n_2049),
.Y(n_2656)
);

NAND2xp33_ASAP7_75t_L g2657 ( 
.A(n_2330),
.B(n_2100),
.Y(n_2657)
);

AO22x2_ASAP7_75t_L g2658 ( 
.A1(n_2524),
.A2(n_2129),
.B1(n_2132),
.B2(n_2117),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2526),
.Y(n_2659)
);

AO22x2_ASAP7_75t_L g2660 ( 
.A1(n_2551),
.A2(n_2163),
.B1(n_2168),
.B2(n_2139),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2516),
.Y(n_2661)
);

NAND2xp33_ASAP7_75t_L g2662 ( 
.A(n_2338),
.B(n_2100),
.Y(n_2662)
);

AO22x2_ASAP7_75t_L g2663 ( 
.A1(n_2457),
.A2(n_2186),
.B1(n_2187),
.B2(n_2175),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2342),
.B(n_1213),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2532),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2333),
.Y(n_2666)
);

AOI22xp5_ASAP7_75t_L g2667 ( 
.A1(n_2435),
.A2(n_2414),
.B1(n_2534),
.B2(n_2523),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2334),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2366),
.B(n_2179),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2363),
.Y(n_2670)
);

NAND2x1p5_ASAP7_75t_L g2671 ( 
.A(n_2544),
.B(n_2026),
.Y(n_2671)
);

OR2x2_ASAP7_75t_L g2672 ( 
.A(n_2504),
.B(n_771),
.Y(n_2672)
);

BUFx2_ASAP7_75t_L g2673 ( 
.A(n_2405),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2365),
.Y(n_2674)
);

AO22x2_ASAP7_75t_L g2675 ( 
.A1(n_2441),
.A2(n_2254),
.B1(n_2260),
.B2(n_2208),
.Y(n_2675)
);

OR2x6_ASAP7_75t_L g2676 ( 
.A(n_2358),
.B(n_2179),
.Y(n_2676)
);

AO22x2_ASAP7_75t_L g2677 ( 
.A1(n_2442),
.A2(n_2271),
.B1(n_2283),
.B2(n_2276),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2383),
.Y(n_2678)
);

OR2x2_ASAP7_75t_SL g2679 ( 
.A(n_2499),
.B(n_2111),
.Y(n_2679)
);

AO22x2_ASAP7_75t_L g2680 ( 
.A1(n_2443),
.A2(n_2257),
.B1(n_1216),
.B2(n_1217),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2408),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2440),
.Y(n_2682)
);

AOI22xp5_ASAP7_75t_SL g2683 ( 
.A1(n_2504),
.A2(n_1216),
.B1(n_1217),
.B2(n_1214),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2377),
.B(n_1214),
.Y(n_2684)
);

AO22x2_ASAP7_75t_L g2685 ( 
.A1(n_2431),
.A2(n_2257),
.B1(n_2278),
.B2(n_2024),
.Y(n_2685)
);

OAI22xp5_ASAP7_75t_SL g2686 ( 
.A1(n_2397),
.A2(n_1784),
.B1(n_1785),
.B2(n_1765),
.Y(n_2686)
);

AO22x2_ASAP7_75t_L g2687 ( 
.A1(n_2433),
.A2(n_2278),
.B1(n_2024),
.B2(n_2307),
.Y(n_2687)
);

OAI221xp5_ASAP7_75t_L g2688 ( 
.A1(n_2326),
.A2(n_1095),
.B1(n_1099),
.B2(n_1098),
.C(n_1091),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2360),
.A2(n_2356),
.B1(n_2380),
.B2(n_2375),
.Y(n_2689)
);

INVx2_ASAP7_75t_SL g2690 ( 
.A(n_2392),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2451),
.Y(n_2691)
);

NAND2x1p5_ASAP7_75t_L g2692 ( 
.A(n_2544),
.B(n_2026),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2483),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2371),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2373),
.Y(n_2695)
);

AND2x2_ASAP7_75t_SL g2696 ( 
.A(n_2404),
.B(n_2290),
.Y(n_2696)
);

AO22x2_ASAP7_75t_L g2697 ( 
.A1(n_2436),
.A2(n_2307),
.B1(n_2087),
.B2(n_2120),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2414),
.B(n_1956),
.Y(n_2698)
);

NAND2x1p5_ASAP7_75t_L g2699 ( 
.A(n_2544),
.B(n_2045),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2490),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_L g2701 ( 
.A(n_2435),
.B(n_2291),
.Y(n_2701)
);

NOR2xp67_ASAP7_75t_L g2702 ( 
.A(n_2476),
.B(n_2045),
.Y(n_2702)
);

NOR2x1_ASAP7_75t_L g2703 ( 
.A(n_2328),
.B(n_1791),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_SL g2704 ( 
.A(n_2520),
.B(n_2045),
.Y(n_2704)
);

AO22x2_ASAP7_75t_L g2705 ( 
.A1(n_2439),
.A2(n_2307),
.B1(n_2087),
.B2(n_2120),
.Y(n_2705)
);

AO22x2_ASAP7_75t_L g2706 ( 
.A1(n_2352),
.A2(n_2145),
.B1(n_2170),
.B2(n_2043),
.Y(n_2706)
);

AND2x2_ASAP7_75t_SL g2707 ( 
.A(n_2469),
.B(n_2114),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2493),
.Y(n_2708)
);

OR2x6_ASAP7_75t_L g2709 ( 
.A(n_2358),
.B(n_2286),
.Y(n_2709)
);

AOI22xp5_ASAP7_75t_L g2710 ( 
.A1(n_2360),
.A2(n_2291),
.B1(n_1904),
.B2(n_2123),
.Y(n_2710)
);

AND2x6_ASAP7_75t_L g2711 ( 
.A(n_2445),
.B(n_2135),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2481),
.Y(n_2712)
);

NAND2xp33_ASAP7_75t_L g2713 ( 
.A(n_2332),
.B(n_2277),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2471),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2473),
.Y(n_2715)
);

AND2x6_ASAP7_75t_L g2716 ( 
.A(n_2445),
.B(n_2135),
.Y(n_2716)
);

AND2x6_ASAP7_75t_L g2717 ( 
.A(n_2391),
.B(n_2135),
.Y(n_2717)
);

INVxp67_ASAP7_75t_L g2718 ( 
.A(n_2339),
.Y(n_2718)
);

CKINVDCx5p33_ASAP7_75t_R g2719 ( 
.A(n_2545),
.Y(n_2719)
);

OAI221xp5_ASAP7_75t_L g2720 ( 
.A1(n_2378),
.A2(n_1104),
.B1(n_1106),
.B2(n_1105),
.C(n_1103),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2423),
.Y(n_2721)
);

AO22x2_ASAP7_75t_L g2722 ( 
.A1(n_2355),
.A2(n_2145),
.B1(n_2170),
.B2(n_2043),
.Y(n_2722)
);

AOI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2356),
.A2(n_2380),
.B1(n_2428),
.B2(n_2401),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2379),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2535),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2535),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2522),
.B(n_2453),
.Y(n_2727)
);

AO22x2_ASAP7_75t_L g2728 ( 
.A1(n_2357),
.A2(n_2176),
.B1(n_2184),
.B2(n_2171),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2415),
.Y(n_2729)
);

AO22x2_ASAP7_75t_L g2730 ( 
.A1(n_2367),
.A2(n_2176),
.B1(n_2184),
.B2(n_2171),
.Y(n_2730)
);

NAND2x1p5_ASAP7_75t_L g2731 ( 
.A(n_2544),
.B(n_2045),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2417),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2453),
.B(n_2114),
.Y(n_2733)
);

NAND2x1p5_ASAP7_75t_L g2734 ( 
.A(n_2353),
.B(n_2052),
.Y(n_2734)
);

NAND3xp33_ASAP7_75t_L g2735 ( 
.A(n_2422),
.B(n_2259),
.C(n_2138),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2419),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2535),
.Y(n_2737)
);

AO22x2_ASAP7_75t_L g2738 ( 
.A1(n_2450),
.A2(n_2258),
.B1(n_2262),
.B2(n_2235),
.Y(n_2738)
);

AOI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2386),
.A2(n_2138),
.B1(n_2123),
.B2(n_2286),
.Y(n_2739)
);

OR2x6_ASAP7_75t_SL g2740 ( 
.A(n_2498),
.B(n_1956),
.Y(n_2740)
);

AO22x2_ASAP7_75t_L g2741 ( 
.A1(n_2452),
.A2(n_2258),
.B1(n_2262),
.B2(n_2235),
.Y(n_2741)
);

AOI22xp5_ASAP7_75t_L g2742 ( 
.A1(n_2486),
.A2(n_2286),
.B1(n_2301),
.B2(n_2233),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2420),
.Y(n_2743)
);

NAND2x1p5_ASAP7_75t_L g2744 ( 
.A(n_2503),
.B(n_2052),
.Y(n_2744)
);

NAND2x1p5_ASAP7_75t_L g2745 ( 
.A(n_2527),
.B(n_2052),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2727),
.B(n_2715),
.Y(n_2746)
);

AOI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2713),
.A2(n_2497),
.B(n_2448),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2729),
.B(n_2732),
.Y(n_2748)
);

OAI21xp5_ASAP7_75t_L g2749 ( 
.A1(n_2735),
.A2(n_2506),
.B(n_2505),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2556),
.B(n_2496),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2736),
.B(n_2314),
.Y(n_2751)
);

A2O1A1Ixp33_ASAP7_75t_L g2752 ( 
.A1(n_2656),
.A2(n_2422),
.B(n_2469),
.C(n_2390),
.Y(n_2752)
);

AOI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2657),
.A2(n_2393),
.B(n_2517),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2592),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2743),
.B(n_2315),
.Y(n_2755)
);

AOI21xp5_ASAP7_75t_L g2756 ( 
.A1(n_2662),
.A2(n_2458),
.B(n_2425),
.Y(n_2756)
);

AOI22x1_ASAP7_75t_L g2757 ( 
.A1(n_2606),
.A2(n_2639),
.B1(n_2745),
.B2(n_2475),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2559),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2576),
.B(n_2590),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2562),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2567),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2569),
.Y(n_2762)
);

INVx3_ASAP7_75t_L g2763 ( 
.A(n_2711),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2573),
.B(n_2429),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2667),
.B(n_2696),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2635),
.B(n_2465),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2724),
.B(n_2560),
.Y(n_2767)
);

O2A1O1Ixp5_ASAP7_75t_L g2768 ( 
.A1(n_2563),
.A2(n_2337),
.B(n_2316),
.C(n_2521),
.Y(n_2768)
);

OAI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2723),
.A2(n_2426),
.B1(n_2424),
.B2(n_2430),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2694),
.B(n_2437),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2570),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2695),
.B(n_2561),
.Y(n_2772)
);

OAI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2689),
.A2(n_2467),
.B1(n_2464),
.B2(n_2382),
.Y(n_2773)
);

AOI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2564),
.A2(n_2486),
.B1(n_2407),
.B2(n_2398),
.Y(n_2774)
);

AOI21xp5_ASAP7_75t_L g2775 ( 
.A1(n_2575),
.A2(n_2539),
.B(n_2537),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2693),
.B(n_2501),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_L g2777 ( 
.A(n_2605),
.B(n_2133),
.Y(n_2777)
);

AOI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2738),
.A2(n_2313),
.B(n_2461),
.Y(n_2778)
);

AOI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_2738),
.A2(n_2313),
.B(n_2463),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2712),
.B(n_2446),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2684),
.B(n_2385),
.Y(n_2781)
);

AO21x1_ASAP7_75t_L g2782 ( 
.A1(n_2733),
.A2(n_2465),
.B(n_2507),
.Y(n_2782)
);

AOI21xp5_ASAP7_75t_L g2783 ( 
.A1(n_2741),
.A2(n_2540),
.B(n_2548),
.Y(n_2783)
);

CKINVDCx20_ASAP7_75t_R g2784 ( 
.A(n_2611),
.Y(n_2784)
);

NOR2xp33_ASAP7_75t_L g2785 ( 
.A(n_2628),
.B(n_2222),
.Y(n_2785)
);

AOI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2741),
.A2(n_2687),
.B(n_2725),
.Y(n_2786)
);

BUFx6f_ASAP7_75t_L g2787 ( 
.A(n_2558),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2555),
.B(n_2485),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2687),
.A2(n_2540),
.B(n_2055),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2664),
.B(n_2487),
.Y(n_2790)
);

OR2x6_ASAP7_75t_L g2791 ( 
.A(n_2709),
.B(n_2460),
.Y(n_2791)
);

NOR2xp33_ASAP7_75t_L g2792 ( 
.A(n_2648),
.B(n_2550),
.Y(n_2792)
);

AOI22xp33_ASAP7_75t_L g2793 ( 
.A1(n_2582),
.A2(n_1520),
.B1(n_1584),
.B2(n_685),
.Y(n_2793)
);

NAND3xp33_ASAP7_75t_L g2794 ( 
.A(n_2554),
.B(n_2478),
.C(n_2484),
.Y(n_2794)
);

AOI21xp5_ASAP7_75t_L g2795 ( 
.A1(n_2726),
.A2(n_2055),
.B(n_2052),
.Y(n_2795)
);

INVx11_ASAP7_75t_L g2796 ( 
.A(n_2595),
.Y(n_2796)
);

O2A1O1Ixp33_ASAP7_75t_L g2797 ( 
.A1(n_2584),
.A2(n_2447),
.B(n_2502),
.C(n_2434),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2599),
.B(n_1107),
.Y(n_2798)
);

A2O1A1Ixp33_ASAP7_75t_L g2799 ( 
.A1(n_2589),
.A2(n_2403),
.B(n_2549),
.C(n_2538),
.Y(n_2799)
);

NOR2xp67_ASAP7_75t_L g2800 ( 
.A(n_2718),
.B(n_2055),
.Y(n_2800)
);

OAI321xp33_ASAP7_75t_L g2801 ( 
.A1(n_2586),
.A2(n_1118),
.A3(n_1114),
.B1(n_1122),
.B2(n_1116),
.C(n_1109),
.Y(n_2801)
);

AOI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_2737),
.A2(n_2059),
.B(n_2055),
.Y(n_2802)
);

AOI21xp33_ASAP7_75t_L g2803 ( 
.A1(n_2618),
.A2(n_2531),
.B(n_2529),
.Y(n_2803)
);

AOI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2697),
.A2(n_2072),
.B(n_2059),
.Y(n_2804)
);

AO21x1_ASAP7_75t_L g2805 ( 
.A1(n_2704),
.A2(n_2546),
.B(n_2543),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2697),
.A2(n_2072),
.B(n_2059),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2596),
.Y(n_2807)
);

OAI22xp5_ASAP7_75t_L g2808 ( 
.A1(n_2707),
.A2(n_2277),
.B1(n_2462),
.B2(n_2545),
.Y(n_2808)
);

AOI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2705),
.A2(n_2072),
.B(n_2059),
.Y(n_2809)
);

NOR2xp33_ASAP7_75t_L g2810 ( 
.A(n_2594),
.B(n_666),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2602),
.B(n_1123),
.Y(n_2811)
);

AOI21xp33_ASAP7_75t_L g2812 ( 
.A1(n_2618),
.A2(n_1543),
.B(n_1538),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2600),
.B(n_1075),
.Y(n_2813)
);

OAI21xp5_ASAP7_75t_L g2814 ( 
.A1(n_2623),
.A2(n_2644),
.B(n_2669),
.Y(n_2814)
);

OAI21xp33_ASAP7_75t_L g2815 ( 
.A1(n_2566),
.A2(n_671),
.B(n_670),
.Y(n_2815)
);

INVx4_ASAP7_75t_L g2816 ( 
.A(n_2557),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2572),
.Y(n_2817)
);

AOI21x1_ASAP7_75t_L g2818 ( 
.A1(n_2685),
.A2(n_1738),
.B(n_1113),
.Y(n_2818)
);

AOI21x1_ASAP7_75t_L g2819 ( 
.A1(n_2685),
.A2(n_1738),
.B(n_1113),
.Y(n_2819)
);

AOI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2705),
.A2(n_2216),
.B(n_2072),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2574),
.B(n_1127),
.Y(n_2821)
);

OAI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2622),
.A2(n_2630),
.B(n_2688),
.Y(n_2822)
);

NOR2xp33_ASAP7_75t_L g2823 ( 
.A(n_2593),
.B(n_673),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2578),
.B(n_2585),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2706),
.A2(n_2241),
.B(n_2216),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2609),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2597),
.B(n_675),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2588),
.B(n_1086),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2598),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2742),
.B(n_2603),
.Y(n_2830)
);

INVx4_ASAP7_75t_L g2831 ( 
.A(n_2719),
.Y(n_2831)
);

BUFx6f_ASAP7_75t_L g2832 ( 
.A(n_2632),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2722),
.A2(n_2241),
.B(n_2216),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2607),
.B(n_1124),
.Y(n_2834)
);

O2A1O1Ixp33_ASAP7_75t_SL g2835 ( 
.A1(n_2583),
.A2(n_1552),
.B(n_1586),
.C(n_1576),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_L g2836 ( 
.A(n_2604),
.B(n_676),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2616),
.B(n_1124),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2721),
.B(n_980),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2722),
.A2(n_2241),
.B(n_2323),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2617),
.B(n_2332),
.Y(n_2840)
);

HB1xp67_ASAP7_75t_L g2841 ( 
.A(n_2568),
.Y(n_2841)
);

O2A1O1Ixp33_ASAP7_75t_L g2842 ( 
.A1(n_2621),
.A2(n_981),
.B(n_990),
.C(n_986),
.Y(n_2842)
);

AND2x4_ASAP7_75t_SL g2843 ( 
.A(n_2632),
.B(n_2323),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2620),
.B(n_2332),
.Y(n_2844)
);

INVxp67_ASAP7_75t_L g2845 ( 
.A(n_2641),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2710),
.A2(n_2535),
.B1(n_1584),
.B2(n_681),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2672),
.B(n_991),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2629),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2631),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2633),
.B(n_2332),
.Y(n_2850)
);

OAI21xp5_ASAP7_75t_L g2851 ( 
.A1(n_2700),
.A2(n_2332),
.B(n_1543),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2610),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2728),
.A2(n_2346),
.B(n_2323),
.Y(n_2853)
);

OAI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2601),
.A2(n_684),
.B1(n_688),
.B2(n_680),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2728),
.A2(n_2613),
.B(n_2568),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2701),
.B(n_690),
.Y(n_2856)
);

AOI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2571),
.A2(n_2346),
.B(n_2323),
.Y(n_2857)
);

AOI21xp5_ASAP7_75t_L g2858 ( 
.A1(n_2571),
.A2(n_2351),
.B(n_2346),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2708),
.A2(n_2351),
.B(n_2346),
.Y(n_2859)
);

AOI33xp33_ASAP7_75t_L g2860 ( 
.A1(n_2638),
.A2(n_996),
.A3(n_993),
.B1(n_999),
.B2(n_997),
.B3(n_994),
.Y(n_2860)
);

INVxp67_ASAP7_75t_L g2861 ( 
.A(n_2673),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2626),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2640),
.B(n_2351),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2581),
.A2(n_704),
.B1(n_705),
.B2(n_696),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2646),
.B(n_2351),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2675),
.A2(n_2374),
.B(n_2368),
.Y(n_2866)
);

OAI321xp33_ASAP7_75t_L g2867 ( 
.A1(n_2739),
.A2(n_1004),
.A3(n_1000),
.B1(n_1006),
.B2(n_1005),
.C(n_1001),
.Y(n_2867)
);

INVx2_ASAP7_75t_SL g2868 ( 
.A(n_2636),
.Y(n_2868)
);

OAI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2720),
.A2(n_2714),
.B(n_2651),
.Y(n_2869)
);

OAI22x1_ASAP7_75t_L g2870 ( 
.A1(n_2650),
.A2(n_1008),
.B1(n_1009),
.B2(n_1007),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_L g2871 ( 
.A(n_2698),
.B(n_706),
.Y(n_2871)
);

O2A1O1Ixp33_ASAP7_75t_L g2872 ( 
.A1(n_2624),
.A2(n_1011),
.B(n_1014),
.C(n_772),
.Y(n_2872)
);

AOI21xp5_ASAP7_75t_L g2873 ( 
.A1(n_2675),
.A2(n_2374),
.B(n_2368),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2652),
.B(n_2368),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2653),
.B(n_2368),
.Y(n_2875)
);

OAI22xp5_ASAP7_75t_L g2876 ( 
.A1(n_2581),
.A2(n_2680),
.B1(n_2582),
.B2(n_2566),
.Y(n_2876)
);

NAND3xp33_ASAP7_75t_L g2877 ( 
.A(n_2683),
.B(n_710),
.C(n_709),
.Y(n_2877)
);

INVx1_ASAP7_75t_SL g2878 ( 
.A(n_2654),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2677),
.A2(n_2416),
.B(n_2374),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2655),
.Y(n_2880)
);

O2A1O1Ixp5_ASAP7_75t_L g2881 ( 
.A1(n_2659),
.A2(n_2299),
.B(n_2308),
.C(n_2287),
.Y(n_2881)
);

O2A1O1Ixp33_ASAP7_75t_L g2882 ( 
.A1(n_2690),
.A2(n_2017),
.B(n_2019),
.C(n_2287),
.Y(n_2882)
);

AOI21xp5_ASAP7_75t_L g2883 ( 
.A1(n_2677),
.A2(n_2416),
.B(n_2374),
.Y(n_2883)
);

AOI21xp5_ASAP7_75t_L g2884 ( 
.A1(n_2663),
.A2(n_2438),
.B(n_2416),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2553),
.B(n_2416),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2661),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2553),
.B(n_2642),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2663),
.A2(n_2449),
.B(n_2438),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2680),
.A2(n_1584),
.B1(n_2535),
.B2(n_1538),
.Y(n_2889)
);

AOI21xp5_ASAP7_75t_L g2890 ( 
.A1(n_2658),
.A2(n_2449),
.B(n_2438),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2658),
.A2(n_2449),
.B(n_2438),
.Y(n_2891)
);

AOI21x1_ASAP7_75t_L g2892 ( 
.A1(n_2627),
.A2(n_1543),
.B(n_1538),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2577),
.B(n_2449),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2645),
.A2(n_2468),
.B(n_2141),
.Y(n_2894)
);

AOI22xp33_ASAP7_75t_L g2895 ( 
.A1(n_2587),
.A2(n_2591),
.B1(n_2565),
.B2(n_2625),
.Y(n_2895)
);

AOI21xp5_ASAP7_75t_L g2896 ( 
.A1(n_2645),
.A2(n_2468),
.B(n_2141),
.Y(n_2896)
);

CKINVDCx8_ASAP7_75t_R g2897 ( 
.A(n_2614),
.Y(n_2897)
);

OAI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2565),
.A2(n_716),
.B1(n_719),
.B2(n_714),
.Y(n_2898)
);

NOR3xp33_ASAP7_75t_L g2899 ( 
.A(n_2686),
.B(n_727),
.C(n_720),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2665),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2580),
.B(n_2468),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2580),
.A2(n_2141),
.B(n_2135),
.Y(n_2902)
);

NOR2xp33_ASAP7_75t_L g2903 ( 
.A(n_2615),
.B(n_731),
.Y(n_2903)
);

OAI21xp5_ASAP7_75t_L g2904 ( 
.A1(n_2734),
.A2(n_1584),
.B(n_2299),
.Y(n_2904)
);

AO32x1_ASAP7_75t_L g2905 ( 
.A1(n_2666),
.A2(n_876),
.A3(n_880),
.B1(n_870),
.B2(n_821),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2625),
.B(n_1092),
.Y(n_2906)
);

AOI21xp5_ASAP7_75t_L g2907 ( 
.A1(n_2637),
.A2(n_2245),
.B(n_2308),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2643),
.Y(n_2908)
);

AOI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2637),
.A2(n_2245),
.B(n_2019),
.Y(n_2909)
);

AOI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2703),
.A2(n_2535),
.B1(n_1584),
.B2(n_738),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2627),
.A2(n_2245),
.B(n_2017),
.Y(n_2911)
);

NOR2x1p5_ASAP7_75t_SL g2912 ( 
.A(n_2670),
.B(n_1092),
.Y(n_2912)
);

INVx3_ASAP7_75t_SL g2913 ( 
.A(n_2679),
.Y(n_2913)
);

O2A1O1Ixp33_ASAP7_75t_L g2914 ( 
.A1(n_2552),
.A2(n_1517),
.B(n_1021),
.C(n_1023),
.Y(n_2914)
);

AOI21xp5_ASAP7_75t_L g2915 ( 
.A1(n_2671),
.A2(n_2245),
.B(n_1495),
.Y(n_2915)
);

O2A1O1Ixp33_ASAP7_75t_L g2916 ( 
.A1(n_2619),
.A2(n_1024),
.B(n_1018),
.C(n_870),
.Y(n_2916)
);

AOI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2709),
.A2(n_1584),
.B1(n_739),
.B2(n_740),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2692),
.A2(n_1489),
.B(n_1483),
.Y(n_2918)
);

AOI21xp33_ASAP7_75t_L g2919 ( 
.A1(n_2587),
.A2(n_1451),
.B(n_1102),
.Y(n_2919)
);

NOR3xp33_ASAP7_75t_L g2920 ( 
.A(n_2702),
.B(n_745),
.C(n_732),
.Y(n_2920)
);

NAND3xp33_ASAP7_75t_L g2921 ( 
.A(n_2668),
.B(n_748),
.C(n_746),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2678),
.B(n_1102),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2699),
.A2(n_1489),
.B(n_1483),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_SL g2924 ( 
.A(n_2634),
.B(n_1518),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2681),
.Y(n_2925)
);

AOI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2731),
.A2(n_1489),
.B(n_1483),
.Y(n_2926)
);

BUFx2_ASAP7_75t_L g2927 ( 
.A(n_2711),
.Y(n_2927)
);

AOI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2730),
.A2(n_1489),
.B(n_1483),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2740),
.B(n_750),
.Y(n_2929)
);

HB1xp67_ASAP7_75t_L g2930 ( 
.A(n_2730),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2682),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2660),
.A2(n_1508),
.B(n_1498),
.Y(n_2932)
);

AOI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2660),
.A2(n_1508),
.B(n_1498),
.Y(n_2933)
);

OAI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2711),
.A2(n_1466),
.B(n_876),
.Y(n_2934)
);

OA21x2_ASAP7_75t_L g2935 ( 
.A1(n_2783),
.A2(n_2691),
.B(n_2674),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2767),
.B(n_2591),
.Y(n_2936)
);

BUFx12f_ASAP7_75t_L g2937 ( 
.A(n_2831),
.Y(n_2937)
);

NOR3xp33_ASAP7_75t_SL g2938 ( 
.A(n_2777),
.B(n_755),
.C(n_751),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2746),
.B(n_2717),
.Y(n_2939)
);

AOI21xp33_ASAP7_75t_L g2940 ( 
.A1(n_2864),
.A2(n_2649),
.B(n_2647),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2747),
.A2(n_2676),
.B(n_2612),
.Y(n_2941)
);

AOI21xp33_ASAP7_75t_L g2942 ( 
.A1(n_2864),
.A2(n_2744),
.B(n_2676),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2754),
.B(n_2717),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_SL g2944 ( 
.A(n_2769),
.B(n_2579),
.Y(n_2944)
);

OAI22xp5_ASAP7_75t_L g2945 ( 
.A1(n_2765),
.A2(n_760),
.B1(n_762),
.B2(n_759),
.Y(n_2945)
);

AO32x2_ASAP7_75t_L g2946 ( 
.A1(n_2876),
.A2(n_2898),
.A3(n_2773),
.B1(n_2769),
.B2(n_2854),
.Y(n_2946)
);

OA21x2_ASAP7_75t_L g2947 ( 
.A1(n_2786),
.A2(n_2779),
.B(n_2778),
.Y(n_2947)
);

O2A1O1Ixp33_ASAP7_75t_L g2948 ( 
.A1(n_2822),
.A2(n_2608),
.B(n_821),
.C(n_903),
.Y(n_2948)
);

AOI22xp33_ASAP7_75t_L g2949 ( 
.A1(n_2822),
.A2(n_2717),
.B1(n_1102),
.B2(n_1451),
.Y(n_2949)
);

BUFx3_ASAP7_75t_L g2950 ( 
.A(n_2784),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2761),
.Y(n_2951)
);

NOR3xp33_ASAP7_75t_L g2952 ( 
.A(n_2854),
.B(n_764),
.C(n_880),
.Y(n_2952)
);

OAI22xp5_ASAP7_75t_L g2953 ( 
.A1(n_2752),
.A2(n_927),
.B1(n_929),
.B2(n_903),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2772),
.B(n_2716),
.Y(n_2954)
);

AOI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2775),
.A2(n_2716),
.B(n_1508),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2756),
.A2(n_2716),
.B(n_1508),
.Y(n_2956)
);

INVxp67_ASAP7_75t_SL g2957 ( 
.A(n_2782),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2789),
.A2(n_1514),
.B(n_1498),
.Y(n_2958)
);

AOI21xp5_ASAP7_75t_L g2959 ( 
.A1(n_2753),
.A2(n_1514),
.B(n_1498),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2764),
.B(n_927),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2758),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2808),
.B(n_1518),
.Y(n_2962)
);

O2A1O1Ixp5_ASAP7_75t_L g2963 ( 
.A1(n_2898),
.A2(n_934),
.B(n_945),
.C(n_929),
.Y(n_2963)
);

OA22x2_ASAP7_75t_L g2964 ( 
.A1(n_2815),
.A2(n_945),
.B1(n_975),
.B2(n_934),
.Y(n_2964)
);

HB1xp67_ASAP7_75t_L g2965 ( 
.A(n_2841),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2748),
.B(n_975),
.Y(n_2966)
);

AOI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2835),
.A2(n_1514),
.B(n_1518),
.Y(n_2967)
);

BUFx8_ASAP7_75t_L g2968 ( 
.A(n_2929),
.Y(n_2968)
);

OAI22x1_ASAP7_75t_L g2969 ( 
.A1(n_2913),
.A2(n_2766),
.B1(n_2887),
.B2(n_2774),
.Y(n_2969)
);

INVx1_ASAP7_75t_SL g2970 ( 
.A(n_2885),
.Y(n_2970)
);

O2A1O1Ixp33_ASAP7_75t_L g2971 ( 
.A1(n_2823),
.A2(n_998),
.B(n_1022),
.C(n_983),
.Y(n_2971)
);

INVx4_ASAP7_75t_L g2972 ( 
.A(n_2787),
.Y(n_2972)
);

OAI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2773),
.A2(n_998),
.B1(n_1022),
.B2(n_983),
.Y(n_2973)
);

OAI21xp33_ASAP7_75t_L g2974 ( 
.A1(n_2827),
.A2(n_511),
.B(n_508),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2760),
.Y(n_2975)
);

AOI21xp5_ASAP7_75t_L g2976 ( 
.A1(n_2825),
.A2(n_1466),
.B(n_1456),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2759),
.B(n_2845),
.Y(n_2977)
);

BUFx8_ASAP7_75t_L g2978 ( 
.A(n_2868),
.Y(n_2978)
);

AOI21xp5_ASAP7_75t_L g2979 ( 
.A1(n_2833),
.A2(n_1456),
.B(n_1454),
.Y(n_2979)
);

BUFx4f_ASAP7_75t_L g2980 ( 
.A(n_2832),
.Y(n_2980)
);

AOI21xp5_ASAP7_75t_L g2981 ( 
.A1(n_2749),
.A2(n_1456),
.B(n_1454),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2776),
.B(n_9),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2751),
.B(n_13),
.Y(n_2983)
);

OAI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_2749),
.A2(n_514),
.B(n_513),
.Y(n_2984)
);

O2A1O1Ixp33_ASAP7_75t_L g2985 ( 
.A1(n_2836),
.A2(n_2811),
.B(n_2798),
.C(n_2856),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2807),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2762),
.Y(n_2987)
);

BUFx2_ASAP7_75t_L g2988 ( 
.A(n_2927),
.Y(n_2988)
);

BUFx2_ASAP7_75t_L g2989 ( 
.A(n_2861),
.Y(n_2989)
);

A2O1A1Ixp33_ASAP7_75t_L g2990 ( 
.A1(n_2855),
.A2(n_519),
.B(n_521),
.C(n_517),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2826),
.Y(n_2991)
);

INVx3_ASAP7_75t_L g2992 ( 
.A(n_2763),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2771),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2755),
.B(n_2824),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2830),
.B(n_13),
.Y(n_2995)
);

OAI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2846),
.A2(n_532),
.B1(n_533),
.B2(n_523),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_R g2997 ( 
.A(n_2897),
.B(n_540),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2817),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2829),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2750),
.B(n_15),
.Y(n_3000)
);

INVx3_ASAP7_75t_L g3001 ( 
.A(n_2763),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2839),
.A2(n_1456),
.B(n_1454),
.Y(n_3002)
);

NOR2xp33_ASAP7_75t_L g3003 ( 
.A(n_2903),
.B(n_16),
.Y(n_3003)
);

OAI21x1_ASAP7_75t_L g3004 ( 
.A1(n_2818),
.A2(n_2819),
.B(n_2902),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2808),
.B(n_1454),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2757),
.B(n_1470),
.Y(n_3006)
);

BUFx3_ASAP7_75t_L g3007 ( 
.A(n_2831),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2848),
.B(n_16),
.Y(n_3008)
);

HB1xp67_ASAP7_75t_L g3009 ( 
.A(n_2863),
.Y(n_3009)
);

AOI21xp5_ASAP7_75t_L g3010 ( 
.A1(n_2804),
.A2(n_1460),
.B(n_1459),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2849),
.Y(n_3011)
);

AO32x2_ASAP7_75t_L g3012 ( 
.A1(n_2876),
.A2(n_21),
.A3(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_3012)
);

BUFx6f_ASAP7_75t_L g3013 ( 
.A(n_2832),
.Y(n_3013)
);

BUFx3_ASAP7_75t_L g3014 ( 
.A(n_2787),
.Y(n_3014)
);

AOI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2806),
.A2(n_1460),
.B(n_1459),
.Y(n_3015)
);

AOI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2809),
.A2(n_1460),
.B(n_1459),
.Y(n_3016)
);

AOI21xp5_ASAP7_75t_L g3017 ( 
.A1(n_2820),
.A2(n_1470),
.B(n_1462),
.Y(n_3017)
);

NAND2x1p5_ASAP7_75t_L g3018 ( 
.A(n_2832),
.B(n_1462),
.Y(n_3018)
);

CKINVDCx5p33_ASAP7_75t_R g3019 ( 
.A(n_2796),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2852),
.Y(n_3020)
);

OAI21x1_ASAP7_75t_L g3021 ( 
.A1(n_2907),
.A2(n_1470),
.B(n_1462),
.Y(n_3021)
);

BUFx12f_ASAP7_75t_L g3022 ( 
.A(n_2816),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2880),
.Y(n_3023)
);

OAI21x1_ASAP7_75t_L g3024 ( 
.A1(n_2866),
.A2(n_2879),
.B(n_2873),
.Y(n_3024)
);

BUFx3_ASAP7_75t_L g3025 ( 
.A(n_2787),
.Y(n_3025)
);

AOI22xp33_ASAP7_75t_L g3026 ( 
.A1(n_2895),
.A2(n_1470),
.B1(n_1462),
.B2(n_548),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2889),
.A2(n_556),
.B1(n_558),
.B2(n_545),
.Y(n_3027)
);

O2A1O1Ixp33_ASAP7_75t_L g3028 ( 
.A1(n_2797),
.A2(n_24),
.B(n_18),
.C(n_19),
.Y(n_3028)
);

AND2x4_ASAP7_75t_L g3029 ( 
.A(n_2930),
.B(n_254),
.Y(n_3029)
);

A2O1A1Ixp33_ASAP7_75t_L g3030 ( 
.A1(n_2801),
.A2(n_574),
.B(n_576),
.C(n_560),
.Y(n_3030)
);

INVx3_ASAP7_75t_L g3031 ( 
.A(n_2843),
.Y(n_3031)
);

NOR3xp33_ASAP7_75t_SL g3032 ( 
.A(n_2785),
.B(n_591),
.C(n_577),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2816),
.B(n_2871),
.Y(n_3033)
);

O2A1O1Ixp33_ASAP7_75t_L g3034 ( 
.A1(n_2799),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_3034)
);

OAI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2794),
.A2(n_597),
.B1(n_598),
.B2(n_594),
.Y(n_3035)
);

AND2x2_ASAP7_75t_L g3036 ( 
.A(n_2813),
.B(n_25),
.Y(n_3036)
);

INVx2_ASAP7_75t_SL g3037 ( 
.A(n_2878),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2925),
.Y(n_3038)
);

OAI22xp5_ASAP7_75t_L g3039 ( 
.A1(n_2781),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_3039)
);

AND2x4_ASAP7_75t_L g3040 ( 
.A(n_2893),
.B(n_255),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2851),
.A2(n_612),
.B(n_606),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2780),
.B(n_28),
.Y(n_3042)
);

AND2x2_ASAP7_75t_SL g3043 ( 
.A(n_2793),
.B(n_780),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2790),
.B(n_29),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2931),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2788),
.B(n_31),
.Y(n_3046)
);

BUFx6f_ASAP7_75t_L g3047 ( 
.A(n_2791),
.Y(n_3047)
);

A2O1A1Ixp33_ASAP7_75t_SL g3048 ( 
.A1(n_2810),
.A2(n_36),
.B(n_33),
.C(n_34),
.Y(n_3048)
);

NOR2x1_ASAP7_75t_R g3049 ( 
.A(n_2770),
.B(n_614),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2814),
.B(n_33),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2886),
.Y(n_3051)
);

OAI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_2792),
.A2(n_621),
.B1(n_630),
.B2(n_616),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2768),
.B(n_635),
.Y(n_3053)
);

OAI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_2910),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_3054)
);

INVx2_ASAP7_75t_SL g3055 ( 
.A(n_2847),
.Y(n_3055)
);

AOI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_2851),
.A2(n_661),
.B(n_660),
.Y(n_3056)
);

BUFx4f_ASAP7_75t_SL g3057 ( 
.A(n_2838),
.Y(n_3057)
);

BUFx2_ASAP7_75t_SL g3058 ( 
.A(n_2800),
.Y(n_3058)
);

AOI21xp5_ASAP7_75t_L g3059 ( 
.A1(n_2928),
.A2(n_674),
.B(n_664),
.Y(n_3059)
);

AOI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2853),
.A2(n_687),
.B(n_686),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2894),
.A2(n_699),
.B(n_689),
.Y(n_3061)
);

NOR3xp33_ASAP7_75t_SL g3062 ( 
.A(n_2814),
.B(n_701),
.C(n_700),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2865),
.B(n_37),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2874),
.B(n_39),
.Y(n_3064)
);

AOI21x1_ASAP7_75t_L g3065 ( 
.A1(n_2906),
.A2(n_794),
.B(n_780),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2875),
.B(n_40),
.Y(n_3066)
);

OAI22xp5_ASAP7_75t_SL g3067 ( 
.A1(n_2877),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_3067)
);

OAI21xp5_ASAP7_75t_L g3068 ( 
.A1(n_2869),
.A2(n_707),
.B(n_702),
.Y(n_3068)
);

BUFx6f_ASAP7_75t_L g3069 ( 
.A(n_2791),
.Y(n_3069)
);

NAND2xp33_ASAP7_75t_SL g3070 ( 
.A(n_2840),
.B(n_725),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2896),
.A2(n_737),
.B(n_726),
.Y(n_3071)
);

O2A1O1Ixp33_ASAP7_75t_L g3072 ( 
.A1(n_2899),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2900),
.Y(n_3073)
);

BUFx6f_ASAP7_75t_L g3074 ( 
.A(n_2791),
.Y(n_3074)
);

O2A1O1Ixp33_ASAP7_75t_L g3075 ( 
.A1(n_2869),
.A2(n_47),
.B(n_44),
.C(n_46),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2828),
.B(n_48),
.Y(n_3076)
);

AOI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_2934),
.A2(n_753),
.B(n_744),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2834),
.B(n_48),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2837),
.B(n_49),
.Y(n_3079)
);

BUFx2_ASAP7_75t_L g3080 ( 
.A(n_2844),
.Y(n_3080)
);

INVx3_ASAP7_75t_L g3081 ( 
.A(n_2850),
.Y(n_3081)
);

INVx2_ASAP7_75t_SL g3082 ( 
.A(n_2901),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2862),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2908),
.B(n_50),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2921),
.B(n_52),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2922),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_2857),
.B(n_256),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2892),
.Y(n_3088)
);

NOR2x1_ASAP7_75t_L g3089 ( 
.A(n_2882),
.B(n_780),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2821),
.Y(n_3090)
);

A2O1A1Ixp33_ASAP7_75t_L g3091 ( 
.A1(n_2867),
.A2(n_756),
.B(n_794),
.C(n_780),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_SL g3092 ( 
.A(n_2805),
.B(n_794),
.Y(n_3092)
);

CKINVDCx5p33_ASAP7_75t_R g3093 ( 
.A(n_2859),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2858),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2890),
.Y(n_3095)
);

O2A1O1Ixp33_ASAP7_75t_L g3096 ( 
.A1(n_2803),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_3096)
);

OR2x2_ASAP7_75t_L g3097 ( 
.A(n_2891),
.B(n_54),
.Y(n_3097)
);

INVx3_ASAP7_75t_SL g3098 ( 
.A(n_2924),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2870),
.Y(n_3099)
);

OAI21xp33_ASAP7_75t_SL g3100 ( 
.A1(n_2917),
.A2(n_55),
.B(n_58),
.Y(n_3100)
);

AOI21xp5_ASAP7_75t_L g3101 ( 
.A1(n_2934),
.A2(n_805),
.B(n_794),
.Y(n_3101)
);

NOR3xp33_ASAP7_75t_SL g3102 ( 
.A(n_2872),
.B(n_59),
.C(n_60),
.Y(n_3102)
);

AOI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2795),
.A2(n_805),
.B(n_794),
.Y(n_3103)
);

OAI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2904),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2883),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2802),
.A2(n_836),
.B(n_805),
.Y(n_3106)
);

O2A1O1Ixp33_ASAP7_75t_L g3107 ( 
.A1(n_2920),
.A2(n_64),
.B(n_61),
.C(n_63),
.Y(n_3107)
);

AOI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_2904),
.A2(n_836),
.B1(n_906),
.B2(n_805),
.Y(n_3108)
);

INVx2_ASAP7_75t_L g3109 ( 
.A(n_2881),
.Y(n_3109)
);

AOI21xp5_ASAP7_75t_L g3110 ( 
.A1(n_2911),
.A2(n_836),
.B(n_805),
.Y(n_3110)
);

OR2x2_ASAP7_75t_L g3111 ( 
.A(n_2884),
.B(n_64),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2860),
.B(n_2909),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2905),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2905),
.Y(n_3114)
);

NOR2x1_ASAP7_75t_L g3115 ( 
.A(n_2888),
.B(n_2914),
.Y(n_3115)
);

O2A1O1Ixp33_ASAP7_75t_L g3116 ( 
.A1(n_2842),
.A2(n_69),
.B(n_65),
.C(n_67),
.Y(n_3116)
);

NOR2xp33_ASAP7_75t_L g3117 ( 
.A(n_2916),
.B(n_71),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2919),
.B(n_71),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2932),
.A2(n_906),
.B(n_836),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2905),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2812),
.B(n_72),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2933),
.B(n_72),
.Y(n_3122)
);

BUFx2_ASAP7_75t_L g3123 ( 
.A(n_2912),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2915),
.Y(n_3124)
);

NAND3xp33_ASAP7_75t_L g3125 ( 
.A(n_2918),
.B(n_906),
.C(n_836),
.Y(n_3125)
);

A2O1A1Ixp33_ASAP7_75t_L g3126 ( 
.A1(n_2923),
.A2(n_909),
.B(n_961),
.C(n_906),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2926),
.B(n_73),
.Y(n_3127)
);

OAI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_2765),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2747),
.A2(n_909),
.B(n_906),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_2747),
.A2(n_961),
.B(n_909),
.Y(n_3130)
);

AOI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2747),
.A2(n_961),
.B(n_909),
.Y(n_3131)
);

BUFx6f_ASAP7_75t_L g3132 ( 
.A(n_2832),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_2750),
.B(n_74),
.Y(n_3133)
);

AOI21x1_ASAP7_75t_SL g3134 ( 
.A1(n_2929),
.A2(n_76),
.B(n_78),
.Y(n_3134)
);

BUFx2_ASAP7_75t_L g3135 ( 
.A(n_2988),
.Y(n_3135)
);

AND2x4_ASAP7_75t_L g3136 ( 
.A(n_3082),
.B(n_78),
.Y(n_3136)
);

INVx3_ASAP7_75t_L g3137 ( 
.A(n_3081),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_3038),
.Y(n_3138)
);

CKINVDCx11_ASAP7_75t_R g3139 ( 
.A(n_2937),
.Y(n_3139)
);

AND2x4_ASAP7_75t_L g3140 ( 
.A(n_3080),
.B(n_79),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2961),
.Y(n_3141)
);

OAI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_3039),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3142)
);

AND2x4_ASAP7_75t_L g3143 ( 
.A(n_2965),
.B(n_3081),
.Y(n_3143)
);

OAI22xp5_ASAP7_75t_L g3144 ( 
.A1(n_3039),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_3144)
);

BUFx2_ASAP7_75t_SL g3145 ( 
.A(n_2950),
.Y(n_3145)
);

INVx1_ASAP7_75t_SL g3146 ( 
.A(n_3093),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2975),
.Y(n_3147)
);

INVx4_ASAP7_75t_L g3148 ( 
.A(n_3098),
.Y(n_3148)
);

AOI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_2956),
.A2(n_961),
.B(n_909),
.Y(n_3149)
);

OAI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_2985),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2994),
.B(n_3009),
.Y(n_3151)
);

INVx5_ASAP7_75t_L g3152 ( 
.A(n_3087),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2957),
.B(n_85),
.Y(n_3153)
);

OR2x6_ASAP7_75t_SL g3154 ( 
.A(n_3019),
.B(n_86),
.Y(n_3154)
);

AOI222xp33_ASAP7_75t_L g3155 ( 
.A1(n_3003),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.C1(n_92),
.C2(n_93),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2987),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2989),
.B(n_92),
.Y(n_3157)
);

BUFx12f_ASAP7_75t_L g3158 ( 
.A(n_2968),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_3045),
.Y(n_3159)
);

BUFx2_ASAP7_75t_L g3160 ( 
.A(n_2943),
.Y(n_3160)
);

CKINVDCx5p33_ASAP7_75t_R g3161 ( 
.A(n_2997),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_3051),
.Y(n_3162)
);

AND2x4_ASAP7_75t_L g3163 ( 
.A(n_2970),
.B(n_94),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2993),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2998),
.B(n_94),
.Y(n_3165)
);

AOI21x1_ASAP7_75t_L g3166 ( 
.A1(n_3092),
.A2(n_963),
.B(n_961),
.Y(n_3166)
);

INVxp67_ASAP7_75t_SL g3167 ( 
.A(n_3088),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2999),
.B(n_95),
.Y(n_3168)
);

NAND2x1p5_ASAP7_75t_L g3169 ( 
.A(n_2944),
.B(n_963),
.Y(n_3169)
);

AOI22xp33_ASAP7_75t_L g3170 ( 
.A1(n_2952),
.A2(n_984),
.B1(n_995),
.B2(n_963),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_3011),
.B(n_95),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_3023),
.B(n_96),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_3073),
.Y(n_3173)
);

BUFx3_ASAP7_75t_L g3174 ( 
.A(n_3007),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2936),
.Y(n_3175)
);

INVxp67_ASAP7_75t_SL g3176 ( 
.A(n_2947),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_3124),
.B(n_96),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_3057),
.B(n_97),
.Y(n_3178)
);

AOI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_3068),
.A2(n_3043),
.B1(n_3067),
.B2(n_3055),
.Y(n_3179)
);

BUFx2_ASAP7_75t_L g3180 ( 
.A(n_3022),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3086),
.Y(n_3181)
);

BUFx6f_ASAP7_75t_L g3182 ( 
.A(n_3013),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_3090),
.B(n_2947),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2977),
.B(n_97),
.Y(n_3184)
);

INVx4_ASAP7_75t_L g3185 ( 
.A(n_2992),
.Y(n_3185)
);

AOI22xp5_ASAP7_75t_L g3186 ( 
.A1(n_3067),
.A2(n_3128),
.B1(n_2974),
.B2(n_2969),
.Y(n_3186)
);

AOI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_3128),
.A2(n_984),
.B1(n_963),
.B2(n_995),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2960),
.B(n_2970),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2954),
.B(n_98),
.Y(n_3189)
);

CKINVDCx5p33_ASAP7_75t_R g3190 ( 
.A(n_2968),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2951),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2986),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2991),
.Y(n_3193)
);

CKINVDCx6p67_ASAP7_75t_R g3194 ( 
.A(n_3036),
.Y(n_3194)
);

HB1xp67_ASAP7_75t_L g3195 ( 
.A(n_3094),
.Y(n_3195)
);

AOI22xp33_ASAP7_75t_L g3196 ( 
.A1(n_3068),
.A2(n_984),
.B1(n_995),
.B2(n_963),
.Y(n_3196)
);

BUFx4f_ASAP7_75t_SL g3197 ( 
.A(n_2978),
.Y(n_3197)
);

CKINVDCx5p33_ASAP7_75t_R g3198 ( 
.A(n_2978),
.Y(n_3198)
);

INVx6_ASAP7_75t_L g3199 ( 
.A(n_3013),
.Y(n_3199)
);

AND2x4_ASAP7_75t_SL g3200 ( 
.A(n_3031),
.B(n_984),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_3020),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3083),
.Y(n_3202)
);

INVx4_ASAP7_75t_L g3203 ( 
.A(n_2992),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2966),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3008),
.Y(n_3205)
);

INVxp67_ASAP7_75t_L g3206 ( 
.A(n_3095),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3111),
.Y(n_3207)
);

OAI22xp33_ASAP7_75t_L g3208 ( 
.A1(n_3104),
.A2(n_102),
.B1(n_98),
.B2(n_100),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3097),
.Y(n_3209)
);

AND2x4_ASAP7_75t_L g3210 ( 
.A(n_3047),
.B(n_100),
.Y(n_3210)
);

INVx5_ASAP7_75t_L g3211 ( 
.A(n_3087),
.Y(n_3211)
);

BUFx2_ASAP7_75t_L g3212 ( 
.A(n_3001),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3105),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2935),
.Y(n_3214)
);

OAI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_3034),
.A2(n_103),
.B(n_104),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_3001),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_2972),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3050),
.B(n_103),
.Y(n_3218)
);

BUFx3_ASAP7_75t_L g3219 ( 
.A(n_3037),
.Y(n_3219)
);

AND2x4_ASAP7_75t_L g3220 ( 
.A(n_3047),
.B(n_105),
.Y(n_3220)
);

INVx5_ASAP7_75t_L g3221 ( 
.A(n_3047),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3033),
.B(n_105),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_3121),
.B(n_108),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2935),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_2938),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_3000),
.B(n_108),
.Y(n_3226)
);

INVx2_ASAP7_75t_L g3227 ( 
.A(n_3024),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2939),
.Y(n_3228)
);

HB1xp67_ASAP7_75t_L g3229 ( 
.A(n_3004),
.Y(n_3229)
);

INVx2_ASAP7_75t_SL g3230 ( 
.A(n_3014),
.Y(n_3230)
);

INVx2_ASAP7_75t_SL g3231 ( 
.A(n_3025),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3084),
.Y(n_3232)
);

BUFx6f_ASAP7_75t_L g3233 ( 
.A(n_3013),
.Y(n_3233)
);

BUFx2_ASAP7_75t_L g3234 ( 
.A(n_2972),
.Y(n_3234)
);

AOI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_2955),
.A2(n_995),
.B(n_984),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_2964),
.A2(n_995),
.B1(n_115),
.B2(n_109),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2946),
.Y(n_3237)
);

NAND2x1_ASAP7_75t_L g3238 ( 
.A(n_3123),
.B(n_114),
.Y(n_3238)
);

BUFx2_ASAP7_75t_L g3239 ( 
.A(n_3069),
.Y(n_3239)
);

AND2x6_ASAP7_75t_L g3240 ( 
.A(n_3029),
.B(n_257),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3133),
.B(n_114),
.Y(n_3241)
);

BUFx2_ASAP7_75t_L g3242 ( 
.A(n_3069),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_3069),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2946),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2946),
.Y(n_3245)
);

OR2x6_ASAP7_75t_L g3246 ( 
.A(n_3005),
.B(n_258),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_3040),
.Y(n_3247)
);

INVx3_ASAP7_75t_L g3248 ( 
.A(n_3074),
.Y(n_3248)
);

INVx3_ASAP7_75t_L g3249 ( 
.A(n_3074),
.Y(n_3249)
);

INVx3_ASAP7_75t_L g3250 ( 
.A(n_3074),
.Y(n_3250)
);

AND2x4_ASAP7_75t_L g3251 ( 
.A(n_3132),
.B(n_115),
.Y(n_3251)
);

OR2x2_ASAP7_75t_L g3252 ( 
.A(n_3042),
.B(n_118),
.Y(n_3252)
);

AND2x4_ASAP7_75t_L g3253 ( 
.A(n_3132),
.B(n_3040),
.Y(n_3253)
);

AOI22xp33_ASAP7_75t_SL g3254 ( 
.A1(n_3029),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_3046),
.B(n_121),
.Y(n_3255)
);

BUFx2_ASAP7_75t_L g3256 ( 
.A(n_3132),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_2980),
.Y(n_3257)
);

NAND2x1p5_ASAP7_75t_L g3258 ( 
.A(n_2962),
.B(n_262),
.Y(n_3258)
);

BUFx3_ASAP7_75t_L g3259 ( 
.A(n_2980),
.Y(n_3259)
);

HB1xp67_ASAP7_75t_L g3260 ( 
.A(n_3109),
.Y(n_3260)
);

OAI22xp5_ASAP7_75t_L g3261 ( 
.A1(n_3104),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_3261)
);

INVx2_ASAP7_75t_SL g3262 ( 
.A(n_3031),
.Y(n_3262)
);

BUFx6f_ASAP7_75t_L g3263 ( 
.A(n_3018),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2982),
.B(n_122),
.Y(n_3264)
);

AND2x4_ASAP7_75t_L g3265 ( 
.A(n_2941),
.B(n_3115),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3122),
.Y(n_3266)
);

BUFx2_ASAP7_75t_L g3267 ( 
.A(n_3063),
.Y(n_3267)
);

BUFx2_ASAP7_75t_L g3268 ( 
.A(n_3064),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2983),
.B(n_125),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_2995),
.B(n_127),
.Y(n_3270)
);

AND2x2_ASAP7_75t_L g3271 ( 
.A(n_3044),
.B(n_128),
.Y(n_3271)
);

AND2x2_ASAP7_75t_L g3272 ( 
.A(n_3066),
.B(n_128),
.Y(n_3272)
);

INVx3_ASAP7_75t_L g3273 ( 
.A(n_3021),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3012),
.Y(n_3274)
);

BUFx2_ASAP7_75t_L g3275 ( 
.A(n_3070),
.Y(n_3275)
);

AND2x4_ASAP7_75t_L g3276 ( 
.A(n_3099),
.B(n_129),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_2973),
.B(n_129),
.Y(n_3277)
);

AOI22xp33_ASAP7_75t_L g3278 ( 
.A1(n_2974),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2973),
.B(n_133),
.Y(n_3279)
);

BUFx8_ASAP7_75t_SL g3280 ( 
.A(n_3076),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3012),
.Y(n_3281)
);

AND2x2_ASAP7_75t_L g3282 ( 
.A(n_3012),
.B(n_133),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3112),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3118),
.B(n_134),
.Y(n_3284)
);

BUFx6f_ASAP7_75t_L g3285 ( 
.A(n_3127),
.Y(n_3285)
);

BUFx3_ASAP7_75t_L g3286 ( 
.A(n_3078),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3113),
.Y(n_3287)
);

AOI22xp5_ASAP7_75t_L g3288 ( 
.A1(n_3054),
.A2(n_2945),
.B1(n_3085),
.B2(n_3102),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_3089),
.B(n_135),
.Y(n_3289)
);

OA22x2_ASAP7_75t_L g3290 ( 
.A1(n_2984),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_3114),
.Y(n_3291)
);

AO22x1_ASAP7_75t_L g3292 ( 
.A1(n_2984),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_3292)
);

BUFx6f_ASAP7_75t_L g3293 ( 
.A(n_3006),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3079),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2958),
.B(n_142),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3120),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2953),
.B(n_142),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3096),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_3058),
.B(n_143),
.Y(n_3299)
);

HB1xp67_ASAP7_75t_L g3300 ( 
.A(n_3065),
.Y(n_3300)
);

AO21x2_ASAP7_75t_L g3301 ( 
.A1(n_3110),
.A2(n_143),
.B(n_144),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3075),
.Y(n_3302)
);

OR2x6_ASAP7_75t_L g3303 ( 
.A(n_3002),
.B(n_263),
.Y(n_3303)
);

NOR2xp67_ASAP7_75t_SL g3304 ( 
.A(n_3053),
.B(n_144),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3032),
.B(n_2942),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2953),
.B(n_147),
.Y(n_3306)
);

BUFx6f_ASAP7_75t_L g3307 ( 
.A(n_3117),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3062),
.B(n_147),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_2940),
.Y(n_3309)
);

BUFx3_ASAP7_75t_L g3310 ( 
.A(n_3049),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_2963),
.Y(n_3311)
);

BUFx6f_ASAP7_75t_L g3312 ( 
.A(n_3125),
.Y(n_3312)
);

BUFx2_ASAP7_75t_R g3313 ( 
.A(n_3134),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3108),
.Y(n_3314)
);

CKINVDCx8_ASAP7_75t_R g3315 ( 
.A(n_2945),
.Y(n_3315)
);

CKINVDCx5p33_ASAP7_75t_R g3316 ( 
.A(n_3052),
.Y(n_3316)
);

AOI22xp33_ASAP7_75t_L g3317 ( 
.A1(n_3054),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_3317)
);

AND2x4_ASAP7_75t_L g3318 ( 
.A(n_2979),
.B(n_148),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2981),
.B(n_149),
.Y(n_3319)
);

NOR2xp33_ASAP7_75t_L g3320 ( 
.A(n_3035),
.B(n_151),
.Y(n_3320)
);

INVx2_ASAP7_75t_L g3321 ( 
.A(n_3108),
.Y(n_3321)
);

BUFx3_ASAP7_75t_L g3322 ( 
.A(n_3125),
.Y(n_3322)
);

AOI22xp33_ASAP7_75t_L g3323 ( 
.A1(n_3100),
.A2(n_151),
.B1(n_152),
.B2(n_155),
.Y(n_3323)
);

INVx3_ASAP7_75t_L g3324 ( 
.A(n_3010),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_3028),
.B(n_152),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2959),
.B(n_155),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3107),
.Y(n_3327)
);

BUFx3_ASAP7_75t_L g3328 ( 
.A(n_2996),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_2990),
.B(n_156),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2948),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_3048),
.Y(n_3331)
);

AND2x2_ASAP7_75t_L g3332 ( 
.A(n_2949),
.B(n_156),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3015),
.B(n_157),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3116),
.Y(n_3334)
);

INVx3_ASAP7_75t_L g3335 ( 
.A(n_3016),
.Y(n_3335)
);

INVx2_ASAP7_75t_SL g3336 ( 
.A(n_3060),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_2971),
.Y(n_3337)
);

INVx3_ASAP7_75t_L g3338 ( 
.A(n_3017),
.Y(n_3338)
);

BUFx2_ASAP7_75t_L g3339 ( 
.A(n_3126),
.Y(n_3339)
);

AOI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_3101),
.A2(n_158),
.B(n_159),
.Y(n_3340)
);

AOI221xp5_ASAP7_75t_L g3341 ( 
.A1(n_3072),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.C(n_162),
.Y(n_3341)
);

BUFx2_ASAP7_75t_L g3342 ( 
.A(n_3030),
.Y(n_3342)
);

NOR2x1_ASAP7_75t_L g3343 ( 
.A(n_3061),
.B(n_161),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3041),
.B(n_162),
.Y(n_3344)
);

AND2x2_ASAP7_75t_L g3345 ( 
.A(n_3135),
.B(n_3071),
.Y(n_3345)
);

NOR2x1_ASAP7_75t_SL g3346 ( 
.A(n_3152),
.B(n_3059),
.Y(n_3346)
);

AOI22xp5_ASAP7_75t_L g3347 ( 
.A1(n_3186),
.A2(n_3026),
.B1(n_3027),
.B2(n_3056),
.Y(n_3347)
);

NOR3xp33_ASAP7_75t_L g3348 ( 
.A(n_3150),
.B(n_3077),
.C(n_3129),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3266),
.B(n_3130),
.Y(n_3349)
);

BUFx3_ASAP7_75t_L g3350 ( 
.A(n_3158),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3181),
.Y(n_3351)
);

AOI22xp33_ASAP7_75t_L g3352 ( 
.A1(n_3342),
.A2(n_3119),
.B1(n_3106),
.B2(n_3103),
.Y(n_3352)
);

AOI21xp5_ASAP7_75t_L g3353 ( 
.A1(n_3340),
.A2(n_3211),
.B(n_3152),
.Y(n_3353)
);

INVx5_ASAP7_75t_L g3354 ( 
.A(n_3240),
.Y(n_3354)
);

OR2x2_ASAP7_75t_L g3355 ( 
.A(n_3151),
.B(n_3131),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3151),
.B(n_3237),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3141),
.Y(n_3357)
);

CKINVDCx20_ASAP7_75t_R g3358 ( 
.A(n_3139),
.Y(n_3358)
);

AOI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3340),
.A2(n_2976),
.B(n_2967),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3147),
.Y(n_3360)
);

INVx1_ASAP7_75t_SL g3361 ( 
.A(n_3146),
.Y(n_3361)
);

INVxp67_ASAP7_75t_SL g3362 ( 
.A(n_3183),
.Y(n_3362)
);

BUFx2_ASAP7_75t_SL g3363 ( 
.A(n_3174),
.Y(n_3363)
);

A2O1A1Ixp33_ASAP7_75t_L g3364 ( 
.A1(n_3288),
.A2(n_3091),
.B(n_164),
.C(n_165),
.Y(n_3364)
);

CKINVDCx5p33_ASAP7_75t_R g3365 ( 
.A(n_3198),
.Y(n_3365)
);

INVx1_ASAP7_75t_SL g3366 ( 
.A(n_3146),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3156),
.Y(n_3367)
);

O2A1O1Ixp5_ASAP7_75t_L g3368 ( 
.A1(n_3150),
.A2(n_163),
.B(n_164),
.C(n_165),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3244),
.B(n_163),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_3138),
.Y(n_3370)
);

INVx1_ASAP7_75t_SL g3371 ( 
.A(n_3145),
.Y(n_3371)
);

BUFx4_ASAP7_75t_SL g3372 ( 
.A(n_3190),
.Y(n_3372)
);

AND2x4_ASAP7_75t_L g3373 ( 
.A(n_3143),
.B(n_166),
.Y(n_3373)
);

AOI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_3152),
.A2(n_166),
.B(n_168),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3160),
.B(n_169),
.Y(n_3375)
);

OA21x2_ASAP7_75t_L g3376 ( 
.A1(n_3183),
.A2(n_170),
.B(n_171),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_3143),
.B(n_170),
.Y(n_3377)
);

OAI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_3315),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_3378)
);

INVx5_ASAP7_75t_L g3379 ( 
.A(n_3240),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_SL g3380 ( 
.A(n_3152),
.B(n_175),
.Y(n_3380)
);

HB1xp67_ASAP7_75t_L g3381 ( 
.A(n_3195),
.Y(n_3381)
);

INVx3_ASAP7_75t_L g3382 ( 
.A(n_3285),
.Y(n_3382)
);

BUFx2_ASAP7_75t_L g3383 ( 
.A(n_3148),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3245),
.B(n_175),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3205),
.B(n_176),
.Y(n_3385)
);

OR2x2_ASAP7_75t_L g3386 ( 
.A(n_3188),
.B(n_176),
.Y(n_3386)
);

AND2x4_ASAP7_75t_L g3387 ( 
.A(n_3211),
.B(n_178),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_3211),
.A2(n_180),
.B(n_181),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_3164),
.Y(n_3389)
);

BUFx2_ASAP7_75t_L g3390 ( 
.A(n_3148),
.Y(n_3390)
);

OR2x6_ASAP7_75t_L g3391 ( 
.A(n_3140),
.B(n_183),
.Y(n_3391)
);

INVx1_ASAP7_75t_SL g3392 ( 
.A(n_3194),
.Y(n_3392)
);

AOI21xp5_ASAP7_75t_L g3393 ( 
.A1(n_3211),
.A2(n_185),
.B(n_186),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3294),
.B(n_185),
.Y(n_3394)
);

BUFx6f_ASAP7_75t_L g3395 ( 
.A(n_3263),
.Y(n_3395)
);

HB1xp67_ASAP7_75t_L g3396 ( 
.A(n_3195),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3267),
.B(n_187),
.Y(n_3397)
);

BUFx6f_ASAP7_75t_L g3398 ( 
.A(n_3263),
.Y(n_3398)
);

OAI22xp5_ASAP7_75t_L g3399 ( 
.A1(n_3179),
.A2(n_3254),
.B1(n_3313),
.B2(n_3328),
.Y(n_3399)
);

INVx3_ASAP7_75t_L g3400 ( 
.A(n_3285),
.Y(n_3400)
);

INVx1_ASAP7_75t_SL g3401 ( 
.A(n_3280),
.Y(n_3401)
);

INVx3_ASAP7_75t_L g3402 ( 
.A(n_3285),
.Y(n_3402)
);

OAI21x1_ASAP7_75t_L g3403 ( 
.A1(n_3273),
.A2(n_3227),
.B(n_3149),
.Y(n_3403)
);

BUFx3_ASAP7_75t_L g3404 ( 
.A(n_3161),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3268),
.B(n_190),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3283),
.B(n_190),
.Y(n_3406)
);

INVx3_ASAP7_75t_L g3407 ( 
.A(n_3185),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3159),
.Y(n_3408)
);

NAND2x1p5_ASAP7_75t_L g3409 ( 
.A(n_3140),
.B(n_3257),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3297),
.A2(n_192),
.B(n_193),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3162),
.Y(n_3411)
);

AOI22xp33_ASAP7_75t_L g3412 ( 
.A1(n_3282),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_3412)
);

AOI21xp33_ASAP7_75t_SL g3413 ( 
.A1(n_3241),
.A2(n_194),
.B(n_195),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3137),
.B(n_197),
.Y(n_3414)
);

INVx2_ASAP7_75t_SL g3415 ( 
.A(n_3219),
.Y(n_3415)
);

AND2x4_ASAP7_75t_L g3416 ( 
.A(n_3137),
.B(n_198),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_3297),
.A2(n_198),
.B(n_199),
.Y(n_3417)
);

AND2x4_ASAP7_75t_L g3418 ( 
.A(n_3212),
.B(n_199),
.Y(n_3418)
);

NAND2x1_ASAP7_75t_SL g3419 ( 
.A(n_3265),
.B(n_200),
.Y(n_3419)
);

BUFx3_ASAP7_75t_L g3420 ( 
.A(n_3197),
.Y(n_3420)
);

INVx3_ASAP7_75t_L g3421 ( 
.A(n_3185),
.Y(n_3421)
);

AND2x4_ASAP7_75t_L g3422 ( 
.A(n_3216),
.B(n_3228),
.Y(n_3422)
);

INVx2_ASAP7_75t_SL g3423 ( 
.A(n_3199),
.Y(n_3423)
);

INVx1_ASAP7_75t_SL g3424 ( 
.A(n_3180),
.Y(n_3424)
);

BUFx2_ASAP7_75t_L g3425 ( 
.A(n_3217),
.Y(n_3425)
);

INVxp67_ASAP7_75t_L g3426 ( 
.A(n_3286),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3173),
.Y(n_3427)
);

CKINVDCx20_ASAP7_75t_R g3428 ( 
.A(n_3310),
.Y(n_3428)
);

OAI22xp5_ASAP7_75t_L g3429 ( 
.A1(n_3254),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_3306),
.A2(n_3265),
.B(n_3215),
.Y(n_3430)
);

BUFx2_ASAP7_75t_L g3431 ( 
.A(n_3234),
.Y(n_3431)
);

AOI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_3306),
.A2(n_203),
.B(n_204),
.Y(n_3432)
);

OAI22xp5_ASAP7_75t_L g3433 ( 
.A1(n_3313),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_3433)
);

AOI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_3215),
.A2(n_205),
.B(n_207),
.Y(n_3434)
);

INVxp67_ASAP7_75t_L g3435 ( 
.A(n_3184),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3213),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3232),
.B(n_207),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_SL g3438 ( 
.A(n_3307),
.B(n_208),
.Y(n_3438)
);

OR2x6_ASAP7_75t_L g3439 ( 
.A(n_3253),
.B(n_210),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3207),
.B(n_211),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3209),
.B(n_212),
.Y(n_3441)
);

BUFx10_ASAP7_75t_L g3442 ( 
.A(n_3178),
.Y(n_3442)
);

CKINVDCx14_ASAP7_75t_R g3443 ( 
.A(n_3154),
.Y(n_3443)
);

BUFx12f_ASAP7_75t_L g3444 ( 
.A(n_3225),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3206),
.B(n_3153),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3206),
.B(n_214),
.Y(n_3446)
);

OAI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_3290),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_3447)
);

A2O1A1Ixp33_ASAP7_75t_L g3448 ( 
.A1(n_3302),
.A2(n_215),
.B(n_217),
.C(n_218),
.Y(n_3448)
);

OR2x2_ASAP7_75t_L g3449 ( 
.A(n_3188),
.B(n_218),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3175),
.Y(n_3450)
);

AO21x1_ASAP7_75t_L g3451 ( 
.A1(n_3153),
.A2(n_219),
.B(n_220),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3296),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_3191),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3287),
.Y(n_3454)
);

INVx2_ASAP7_75t_L g3455 ( 
.A(n_3201),
.Y(n_3455)
);

AOI222xp33_ASAP7_75t_L g3456 ( 
.A1(n_3334),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.C1(n_226),
.C2(n_227),
.Y(n_3456)
);

CKINVDCx8_ASAP7_75t_R g3457 ( 
.A(n_3316),
.Y(n_3457)
);

INVx2_ASAP7_75t_SL g3458 ( 
.A(n_3199),
.Y(n_3458)
);

AND2x2_ASAP7_75t_L g3459 ( 
.A(n_3216),
.B(n_222),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3230),
.B(n_3231),
.Y(n_3460)
);

INVx1_ASAP7_75t_SL g3461 ( 
.A(n_3222),
.Y(n_3461)
);

CKINVDCx8_ASAP7_75t_R g3462 ( 
.A(n_3307),
.Y(n_3462)
);

AND2x4_ASAP7_75t_L g3463 ( 
.A(n_3203),
.B(n_226),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3192),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3176),
.A2(n_227),
.B(n_228),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3274),
.B(n_229),
.Y(n_3466)
);

OAI21xp33_ASAP7_75t_L g3467 ( 
.A1(n_3155),
.A2(n_229),
.B(n_230),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3281),
.B(n_231),
.Y(n_3468)
);

A2O1A1Ixp33_ASAP7_75t_L g3469 ( 
.A1(n_3327),
.A2(n_232),
.B(n_233),
.C(n_234),
.Y(n_3469)
);

NOR2xp67_ASAP7_75t_SL g3470 ( 
.A(n_3275),
.B(n_234),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3291),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3204),
.B(n_235),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3260),
.Y(n_3473)
);

AND2x4_ASAP7_75t_L g3474 ( 
.A(n_3203),
.B(n_237),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_3262),
.B(n_238),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3260),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3177),
.B(n_238),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_3193),
.Y(n_3478)
);

NAND2x1p5_ASAP7_75t_L g3479 ( 
.A(n_3259),
.B(n_239),
.Y(n_3479)
);

OR2x2_ASAP7_75t_L g3480 ( 
.A(n_3309),
.B(n_240),
.Y(n_3480)
);

INVx3_ASAP7_75t_L g3481 ( 
.A(n_3199),
.Y(n_3481)
);

NOR2xp33_ASAP7_75t_L g3482 ( 
.A(n_3184),
.B(n_3252),
.Y(n_3482)
);

BUFx3_ASAP7_75t_L g3483 ( 
.A(n_3239),
.Y(n_3483)
);

INVx2_ASAP7_75t_SL g3484 ( 
.A(n_3182),
.Y(n_3484)
);

OAI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3290),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_3485)
);

AND2x4_ASAP7_75t_L g3486 ( 
.A(n_3256),
.B(n_243),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3167),
.Y(n_3487)
);

NAND2x1p5_ASAP7_75t_L g3488 ( 
.A(n_3221),
.B(n_243),
.Y(n_3488)
);

AND2x4_ASAP7_75t_L g3489 ( 
.A(n_3243),
.B(n_245),
.Y(n_3489)
);

AOI21x1_ASAP7_75t_L g3490 ( 
.A1(n_3177),
.A2(n_246),
.B(n_247),
.Y(n_3490)
);

BUFx2_ASAP7_75t_L g3491 ( 
.A(n_3182),
.Y(n_3491)
);

HB1xp67_ASAP7_75t_L g3492 ( 
.A(n_3167),
.Y(n_3492)
);

OAI22xp5_ASAP7_75t_L g3493 ( 
.A1(n_3317),
.A2(n_3261),
.B1(n_3307),
.B2(n_3208),
.Y(n_3493)
);

AOI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_3176),
.A2(n_247),
.B(n_248),
.Y(n_3494)
);

BUFx2_ASAP7_75t_L g3495 ( 
.A(n_3182),
.Y(n_3495)
);

OAI22xp5_ASAP7_75t_L g3496 ( 
.A1(n_3261),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3163),
.B(n_250),
.Y(n_3497)
);

AND2x4_ASAP7_75t_L g3498 ( 
.A(n_3243),
.B(n_264),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3157),
.B(n_267),
.Y(n_3499)
);

AND2x4_ASAP7_75t_L g3500 ( 
.A(n_3248),
.B(n_268),
.Y(n_3500)
);

AND2x4_ASAP7_75t_L g3501 ( 
.A(n_3248),
.B(n_270),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3202),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3319),
.A2(n_271),
.B(n_272),
.Y(n_3503)
);

INVx3_ASAP7_75t_L g3504 ( 
.A(n_3233),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3163),
.B(n_273),
.Y(n_3505)
);

AOI21xp33_ASAP7_75t_L g3506 ( 
.A1(n_3298),
.A2(n_274),
.B(n_276),
.Y(n_3506)
);

INVx2_ASAP7_75t_SL g3507 ( 
.A(n_3233),
.Y(n_3507)
);

INVx4_ASAP7_75t_L g3508 ( 
.A(n_3233),
.Y(n_3508)
);

AND2x4_ASAP7_75t_L g3509 ( 
.A(n_3249),
.B(n_278),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3189),
.B(n_286),
.Y(n_3510)
);

INVx3_ASAP7_75t_L g3511 ( 
.A(n_3249),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3165),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3224),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3214),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3473),
.Y(n_3515)
);

INVx1_ASAP7_75t_SL g3516 ( 
.A(n_3425),
.Y(n_3516)
);

AOI22xp33_ASAP7_75t_L g3517 ( 
.A1(n_3399),
.A2(n_3331),
.B1(n_3336),
.B2(n_3240),
.Y(n_3517)
);

BUFx3_ASAP7_75t_L g3518 ( 
.A(n_3358),
.Y(n_3518)
);

BUFx2_ASAP7_75t_L g3519 ( 
.A(n_3383),
.Y(n_3519)
);

CKINVDCx5p33_ASAP7_75t_R g3520 ( 
.A(n_3372),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3362),
.B(n_3165),
.Y(n_3521)
);

BUFx6f_ASAP7_75t_L g3522 ( 
.A(n_3420),
.Y(n_3522)
);

AND2x2_ASAP7_75t_L g3523 ( 
.A(n_3431),
.B(n_3229),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3473),
.Y(n_3524)
);

CKINVDCx20_ASAP7_75t_R g3525 ( 
.A(n_3428),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3467),
.A2(n_3240),
.B1(n_3325),
.B2(n_3155),
.Y(n_3526)
);

AOI22xp33_ASAP7_75t_L g3527 ( 
.A1(n_3433),
.A2(n_3240),
.B1(n_3325),
.B2(n_3208),
.Y(n_3527)
);

BUFx10_ASAP7_75t_L g3528 ( 
.A(n_3365),
.Y(n_3528)
);

CKINVDCx11_ASAP7_75t_R g3529 ( 
.A(n_3457),
.Y(n_3529)
);

CKINVDCx11_ASAP7_75t_R g3530 ( 
.A(n_3444),
.Y(n_3530)
);

INVx1_ASAP7_75t_SL g3531 ( 
.A(n_3361),
.Y(n_3531)
);

INVx6_ASAP7_75t_L g3532 ( 
.A(n_3354),
.Y(n_3532)
);

AND2x2_ASAP7_75t_L g3533 ( 
.A(n_3483),
.B(n_3229),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3452),
.Y(n_3534)
);

AOI22xp33_ASAP7_75t_SL g3535 ( 
.A1(n_3354),
.A2(n_3276),
.B1(n_3142),
.B2(n_3144),
.Y(n_3535)
);

INVx8_ASAP7_75t_L g3536 ( 
.A(n_3439),
.Y(n_3536)
);

HB1xp67_ASAP7_75t_L g3537 ( 
.A(n_3381),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3447),
.A2(n_3144),
.B1(n_3142),
.B2(n_3292),
.Y(n_3538)
);

CKINVDCx11_ASAP7_75t_R g3539 ( 
.A(n_3401),
.Y(n_3539)
);

CKINVDCx11_ASAP7_75t_R g3540 ( 
.A(n_3442),
.Y(n_3540)
);

CKINVDCx11_ASAP7_75t_R g3541 ( 
.A(n_3442),
.Y(n_3541)
);

NAND2x1p5_ASAP7_75t_L g3542 ( 
.A(n_3354),
.B(n_3221),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3452),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3476),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3357),
.Y(n_3545)
);

BUFx3_ASAP7_75t_L g3546 ( 
.A(n_3404),
.Y(n_3546)
);

CKINVDCx14_ASAP7_75t_R g3547 ( 
.A(n_3443),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3476),
.Y(n_3548)
);

AOI22xp33_ASAP7_75t_L g3549 ( 
.A1(n_3485),
.A2(n_3343),
.B1(n_3341),
.B2(n_3329),
.Y(n_3549)
);

BUFx3_ASAP7_75t_L g3550 ( 
.A(n_3350),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3357),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3514),
.Y(n_3552)
);

AOI22xp33_ASAP7_75t_L g3553 ( 
.A1(n_3348),
.A2(n_3451),
.B1(n_3434),
.B2(n_3347),
.Y(n_3553)
);

INVx6_ASAP7_75t_L g3554 ( 
.A(n_3379),
.Y(n_3554)
);

INVx5_ASAP7_75t_SL g3555 ( 
.A(n_3439),
.Y(n_3555)
);

CKINVDCx6p67_ASAP7_75t_R g3556 ( 
.A(n_3391),
.Y(n_3556)
);

AOI22xp33_ASAP7_75t_SL g3557 ( 
.A1(n_3379),
.A2(n_3493),
.B1(n_3376),
.B2(n_3430),
.Y(n_3557)
);

AOI22xp33_ASAP7_75t_L g3558 ( 
.A1(n_3376),
.A2(n_3341),
.B1(n_3344),
.B2(n_3305),
.Y(n_3558)
);

CKINVDCx6p67_ASAP7_75t_R g3559 ( 
.A(n_3391),
.Y(n_3559)
);

CKINVDCx11_ASAP7_75t_R g3560 ( 
.A(n_3424),
.Y(n_3560)
);

BUFx10_ASAP7_75t_L g3561 ( 
.A(n_3463),
.Y(n_3561)
);

OAI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3368),
.A2(n_3344),
.B(n_3319),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3367),
.Y(n_3563)
);

AOI22xp33_ASAP7_75t_L g3564 ( 
.A1(n_3429),
.A2(n_3247),
.B1(n_3330),
.B2(n_3320),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3367),
.Y(n_3565)
);

INVxp67_ASAP7_75t_L g3566 ( 
.A(n_3445),
.Y(n_3566)
);

BUFx6f_ASAP7_75t_L g3567 ( 
.A(n_3379),
.Y(n_3567)
);

INVx2_ASAP7_75t_SL g3568 ( 
.A(n_3460),
.Y(n_3568)
);

INVx6_ASAP7_75t_L g3569 ( 
.A(n_3387),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3389),
.Y(n_3570)
);

INVx3_ASAP7_75t_L g3571 ( 
.A(n_3407),
.Y(n_3571)
);

AOI22xp33_ASAP7_75t_L g3572 ( 
.A1(n_3482),
.A2(n_3255),
.B1(n_3276),
.B2(n_3304),
.Y(n_3572)
);

AOI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_3496),
.A2(n_3271),
.B1(n_3226),
.B2(n_3308),
.Y(n_3573)
);

BUFx6f_ASAP7_75t_L g3574 ( 
.A(n_3387),
.Y(n_3574)
);

BUFx3_ASAP7_75t_L g3575 ( 
.A(n_3415),
.Y(n_3575)
);

OAI22xp33_ASAP7_75t_L g3576 ( 
.A1(n_3353),
.A2(n_3246),
.B1(n_3480),
.B2(n_3461),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3389),
.Y(n_3577)
);

BUFx2_ASAP7_75t_L g3578 ( 
.A(n_3390),
.Y(n_3578)
);

AOI22xp33_ASAP7_75t_L g3579 ( 
.A1(n_3456),
.A2(n_3323),
.B1(n_3332),
.B2(n_3136),
.Y(n_3579)
);

AND2x4_ASAP7_75t_L g3580 ( 
.A(n_3382),
.B(n_3136),
.Y(n_3580)
);

AOI22xp5_ASAP7_75t_L g3581 ( 
.A1(n_3380),
.A2(n_3210),
.B1(n_3220),
.B2(n_3253),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3408),
.Y(n_3582)
);

NAND2xp33_ASAP7_75t_R g3583 ( 
.A(n_3418),
.B(n_3299),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3513),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3408),
.Y(n_3585)
);

BUFx2_ASAP7_75t_L g3586 ( 
.A(n_3481),
.Y(n_3586)
);

INVx1_ASAP7_75t_SL g3587 ( 
.A(n_3366),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3427),
.Y(n_3588)
);

INVx1_ASAP7_75t_SL g3589 ( 
.A(n_3371),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3427),
.Y(n_3590)
);

INVx1_ASAP7_75t_SL g3591 ( 
.A(n_3363),
.Y(n_3591)
);

INVx6_ASAP7_75t_L g3592 ( 
.A(n_3395),
.Y(n_3592)
);

CKINVDCx5p33_ASAP7_75t_R g3593 ( 
.A(n_3392),
.Y(n_3593)
);

BUFx3_ASAP7_75t_L g3594 ( 
.A(n_3409),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3436),
.Y(n_3595)
);

OAI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_3412),
.A2(n_3278),
.B1(n_3223),
.B2(n_3289),
.Y(n_3596)
);

CKINVDCx20_ASAP7_75t_R g3597 ( 
.A(n_3462),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3396),
.B(n_3168),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3487),
.Y(n_3599)
);

OAI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_3374),
.A2(n_3246),
.B1(n_3393),
.B2(n_3388),
.Y(n_3600)
);

AOI22xp33_ASAP7_75t_SL g3601 ( 
.A1(n_3375),
.A2(n_3284),
.B1(n_3223),
.B2(n_3210),
.Y(n_3601)
);

AOI22xp33_ASAP7_75t_L g3602 ( 
.A1(n_3465),
.A2(n_3301),
.B1(n_3337),
.B2(n_3321),
.Y(n_3602)
);

INVx2_ASAP7_75t_L g3603 ( 
.A(n_3487),
.Y(n_3603)
);

INVx6_ASAP7_75t_L g3604 ( 
.A(n_3395),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3492),
.Y(n_3605)
);

AOI22xp5_ASAP7_75t_L g3606 ( 
.A1(n_3378),
.A2(n_3220),
.B1(n_3272),
.B2(n_3218),
.Y(n_3606)
);

BUFx2_ASAP7_75t_L g3607 ( 
.A(n_3481),
.Y(n_3607)
);

CKINVDCx6p67_ASAP7_75t_R g3608 ( 
.A(n_3486),
.Y(n_3608)
);

AOI22xp33_ASAP7_75t_L g3609 ( 
.A1(n_3494),
.A2(n_3301),
.B1(n_3314),
.B2(n_3218),
.Y(n_3609)
);

OAI22xp5_ASAP7_75t_L g3610 ( 
.A1(n_3446),
.A2(n_3289),
.B1(n_3279),
.B2(n_3277),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3351),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3454),
.Y(n_3612)
);

OAI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_3448),
.A2(n_3279),
.B1(n_3277),
.B2(n_3295),
.Y(n_3613)
);

OAI21xp5_ASAP7_75t_SL g3614 ( 
.A1(n_3413),
.A2(n_3270),
.B(n_3269),
.Y(n_3614)
);

OAI22xp5_ASAP7_75t_L g3615 ( 
.A1(n_3469),
.A2(n_3295),
.B1(n_3333),
.B2(n_3326),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_3410),
.A2(n_3236),
.B1(n_3311),
.B2(n_3339),
.Y(n_3616)
);

AOI22xp33_ASAP7_75t_SL g3617 ( 
.A1(n_3466),
.A2(n_3322),
.B1(n_3251),
.B2(n_3246),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3351),
.Y(n_3618)
);

INVx2_ASAP7_75t_SL g3619 ( 
.A(n_3422),
.Y(n_3619)
);

BUFx10_ASAP7_75t_L g3620 ( 
.A(n_3463),
.Y(n_3620)
);

BUFx12f_ASAP7_75t_L g3621 ( 
.A(n_3479),
.Y(n_3621)
);

BUFx3_ASAP7_75t_L g3622 ( 
.A(n_3373),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3454),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3471),
.Y(n_3624)
);

OAI22xp5_ASAP7_75t_L g3625 ( 
.A1(n_3435),
.A2(n_3333),
.B1(n_3326),
.B2(n_3189),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3360),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3370),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3411),
.Y(n_3628)
);

OAI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_3468),
.A2(n_3270),
.B1(n_3269),
.B2(n_3264),
.Y(n_3629)
);

AOI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3417),
.A2(n_3293),
.B1(n_3318),
.B2(n_3242),
.Y(n_3630)
);

BUFx3_ASAP7_75t_L g3631 ( 
.A(n_3373),
.Y(n_3631)
);

CKINVDCx20_ASAP7_75t_R g3632 ( 
.A(n_3426),
.Y(n_3632)
);

INVx6_ASAP7_75t_L g3633 ( 
.A(n_3395),
.Y(n_3633)
);

CKINVDCx8_ASAP7_75t_R g3634 ( 
.A(n_3418),
.Y(n_3634)
);

OAI22xp5_ASAP7_75t_L g3635 ( 
.A1(n_3386),
.A2(n_3264),
.B1(n_3171),
.B2(n_3172),
.Y(n_3635)
);

OAI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3449),
.A2(n_3369),
.B1(n_3384),
.B2(n_3364),
.Y(n_3636)
);

OAI22xp5_ASAP7_75t_SL g3637 ( 
.A1(n_3397),
.A2(n_3238),
.B1(n_3171),
.B2(n_3168),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3422),
.B(n_3250),
.Y(n_3638)
);

INVx4_ASAP7_75t_L g3639 ( 
.A(n_3474),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3450),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3471),
.Y(n_3641)
);

INVx1_ASAP7_75t_SL g3642 ( 
.A(n_3419),
.Y(n_3642)
);

AOI22xp33_ASAP7_75t_L g3643 ( 
.A1(n_3432),
.A2(n_3293),
.B1(n_3318),
.B2(n_3312),
.Y(n_3643)
);

INVx1_ASAP7_75t_SL g3644 ( 
.A(n_3382),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3512),
.Y(n_3645)
);

BUFx4f_ASAP7_75t_SL g3646 ( 
.A(n_3486),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3512),
.B(n_3250),
.Y(n_3647)
);

AOI22xp33_ASAP7_75t_L g3648 ( 
.A1(n_3503),
.A2(n_3293),
.B1(n_3312),
.B2(n_3187),
.Y(n_3648)
);

AOI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3356),
.A2(n_3312),
.B1(n_3251),
.B2(n_3303),
.Y(n_3649)
);

INVx2_ASAP7_75t_L g3650 ( 
.A(n_3515),
.Y(n_3650)
);

BUFx3_ASAP7_75t_L g3651 ( 
.A(n_3525),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_SL g3652 ( 
.A(n_3557),
.B(n_3567),
.Y(n_3652)
);

HB1xp67_ASAP7_75t_L g3653 ( 
.A(n_3537),
.Y(n_3653)
);

HB1xp67_ASAP7_75t_L g3654 ( 
.A(n_3521),
.Y(n_3654)
);

INVxp67_ASAP7_75t_L g3655 ( 
.A(n_3519),
.Y(n_3655)
);

INVx3_ASAP7_75t_L g3656 ( 
.A(n_3639),
.Y(n_3656)
);

HB1xp67_ASAP7_75t_L g3657 ( 
.A(n_3521),
.Y(n_3657)
);

BUFx6f_ASAP7_75t_L g3658 ( 
.A(n_3530),
.Y(n_3658)
);

OAI21x1_ASAP7_75t_L g3659 ( 
.A1(n_3571),
.A2(n_3403),
.B(n_3355),
.Y(n_3659)
);

BUFx4f_ASAP7_75t_SL g3660 ( 
.A(n_3518),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3625),
.B(n_3349),
.Y(n_3661)
);

HB1xp67_ASAP7_75t_L g3662 ( 
.A(n_3605),
.Y(n_3662)
);

CKINVDCx6p67_ASAP7_75t_R g3663 ( 
.A(n_3539),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3524),
.Y(n_3664)
);

OA21x2_ASAP7_75t_L g3665 ( 
.A1(n_3553),
.A2(n_3414),
.B(n_3406),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3545),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3551),
.Y(n_3667)
);

INVx1_ASAP7_75t_SL g3668 ( 
.A(n_3560),
.Y(n_3668)
);

AOI22xp33_ASAP7_75t_SL g3669 ( 
.A1(n_3636),
.A2(n_3346),
.B1(n_3497),
.B2(n_3499),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3625),
.B(n_3345),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3563),
.Y(n_3671)
);

BUFx6f_ASAP7_75t_L g3672 ( 
.A(n_3567),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3565),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3570),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3516),
.B(n_3423),
.Y(n_3675)
);

OR2x2_ASAP7_75t_L g3676 ( 
.A(n_3598),
.B(n_3566),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3544),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3577),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3611),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3618),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_3548),
.Y(n_3681)
);

AOI22xp33_ASAP7_75t_L g3682 ( 
.A1(n_3526),
.A2(n_3506),
.B1(n_3470),
.B2(n_3438),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3645),
.Y(n_3683)
);

OR2x2_ASAP7_75t_L g3684 ( 
.A(n_3598),
.B(n_3516),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3534),
.Y(n_3685)
);

BUFx6f_ASAP7_75t_L g3686 ( 
.A(n_3567),
.Y(n_3686)
);

OAI22xp5_ASAP7_75t_L g3687 ( 
.A1(n_3535),
.A2(n_3416),
.B1(n_3474),
.B2(n_3488),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3543),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3599),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3582),
.Y(n_3690)
);

INVx2_ASAP7_75t_L g3691 ( 
.A(n_3603),
.Y(n_3691)
);

OR2x6_ASAP7_75t_L g3692 ( 
.A(n_3536),
.B(n_3359),
.Y(n_3692)
);

AND2x4_ASAP7_75t_L g3693 ( 
.A(n_3639),
.B(n_3407),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3612),
.Y(n_3694)
);

BUFx8_ASAP7_75t_SL g3695 ( 
.A(n_3520),
.Y(n_3695)
);

INVx4_ASAP7_75t_L g3696 ( 
.A(n_3522),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3623),
.Y(n_3697)
);

BUFx2_ASAP7_75t_L g3698 ( 
.A(n_3547),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3624),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3585),
.Y(n_3700)
);

BUFx2_ASAP7_75t_L g3701 ( 
.A(n_3523),
.Y(n_3701)
);

INVx3_ASAP7_75t_L g3702 ( 
.A(n_3634),
.Y(n_3702)
);

BUFx2_ASAP7_75t_L g3703 ( 
.A(n_3578),
.Y(n_3703)
);

INVx1_ASAP7_75t_SL g3704 ( 
.A(n_3529),
.Y(n_3704)
);

BUFx2_ASAP7_75t_L g3705 ( 
.A(n_3597),
.Y(n_3705)
);

AO21x2_ASAP7_75t_L g3706 ( 
.A1(n_3562),
.A2(n_3477),
.B(n_3472),
.Y(n_3706)
);

OR2x2_ASAP7_75t_L g3707 ( 
.A(n_3531),
.B(n_3587),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3610),
.B(n_3405),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3588),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3586),
.B(n_3458),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3552),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3584),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3590),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3595),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3641),
.Y(n_3715)
);

OAI21x1_ASAP7_75t_SL g3716 ( 
.A1(n_3517),
.A2(n_3614),
.B(n_3610),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3626),
.Y(n_3717)
);

INVx6_ASAP7_75t_L g3718 ( 
.A(n_3536),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3640),
.Y(n_3719)
);

INVx2_ASAP7_75t_L g3720 ( 
.A(n_3647),
.Y(n_3720)
);

BUFx2_ASAP7_75t_L g3721 ( 
.A(n_3533),
.Y(n_3721)
);

INVx2_ASAP7_75t_SL g3722 ( 
.A(n_3561),
.Y(n_3722)
);

OR2x6_ASAP7_75t_L g3723 ( 
.A(n_3536),
.B(n_3169),
.Y(n_3723)
);

INVx6_ASAP7_75t_L g3724 ( 
.A(n_3528),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3627),
.Y(n_3725)
);

CKINVDCx5p33_ASAP7_75t_R g3726 ( 
.A(n_3593),
.Y(n_3726)
);

BUFx3_ASAP7_75t_L g3727 ( 
.A(n_3522),
.Y(n_3727)
);

OAI21x1_ASAP7_75t_L g3728 ( 
.A1(n_3571),
.A2(n_3421),
.B(n_3402),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3628),
.Y(n_3729)
);

CKINVDCx16_ASAP7_75t_R g3730 ( 
.A(n_3583),
.Y(n_3730)
);

AND2x4_ASAP7_75t_L g3731 ( 
.A(n_3574),
.B(n_3421),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3569),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3635),
.Y(n_3733)
);

INVx3_ASAP7_75t_L g3734 ( 
.A(n_3532),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3558),
.A2(n_3478),
.B1(n_3464),
.B2(n_3502),
.Y(n_3735)
);

BUFx3_ASAP7_75t_L g3736 ( 
.A(n_3522),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3635),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3629),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3569),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3629),
.Y(n_3740)
);

BUFx3_ASAP7_75t_L g3741 ( 
.A(n_3528),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3531),
.Y(n_3742)
);

BUFx3_ASAP7_75t_L g3743 ( 
.A(n_3540),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3607),
.B(n_3491),
.Y(n_3744)
);

INVx2_ASAP7_75t_SL g3745 ( 
.A(n_3561),
.Y(n_3745)
);

OAI22xp5_ASAP7_75t_L g3746 ( 
.A1(n_3527),
.A2(n_3416),
.B1(n_3489),
.B2(n_3377),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3587),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3576),
.Y(n_3748)
);

BUFx6f_ASAP7_75t_L g3749 ( 
.A(n_3541),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3589),
.Y(n_3750)
);

AOI21x1_ASAP7_75t_L g3751 ( 
.A1(n_3636),
.A2(n_3437),
.B(n_3385),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3589),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3580),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3580),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3615),
.Y(n_3755)
);

OAI21x1_ASAP7_75t_L g3756 ( 
.A1(n_3542),
.A2(n_3400),
.B(n_3402),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3615),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3569),
.Y(n_3758)
);

AOI22xp33_ASAP7_75t_L g3759 ( 
.A1(n_3549),
.A2(n_3400),
.B1(n_3505),
.B2(n_3510),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3644),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3644),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3568),
.B(n_3495),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3562),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3532),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3613),
.Y(n_3765)
);

OR2x6_ASAP7_75t_L g3766 ( 
.A(n_3532),
.B(n_3169),
.Y(n_3766)
);

AOI21x1_ASAP7_75t_L g3767 ( 
.A1(n_3596),
.A2(n_3394),
.B(n_3441),
.Y(n_3767)
);

BUFx2_ASAP7_75t_SL g3768 ( 
.A(n_3591),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3554),
.Y(n_3769)
);

INVx3_ASAP7_75t_L g3770 ( 
.A(n_3554),
.Y(n_3770)
);

BUFx2_ASAP7_75t_L g3771 ( 
.A(n_3646),
.Y(n_3771)
);

INVx3_ASAP7_75t_L g3772 ( 
.A(n_3554),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3638),
.B(n_3511),
.Y(n_3773)
);

BUFx2_ASAP7_75t_L g3774 ( 
.A(n_3608),
.Y(n_3774)
);

BUFx6f_ASAP7_75t_L g3775 ( 
.A(n_3550),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3690),
.Y(n_3776)
);

AND2x2_ASAP7_75t_L g3777 ( 
.A(n_3701),
.B(n_3591),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3690),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3707),
.Y(n_3779)
);

OA21x2_ASAP7_75t_L g3780 ( 
.A1(n_3659),
.A2(n_3609),
.B(n_3602),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3707),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3734),
.B(n_3620),
.Y(n_3782)
);

AND2x2_ASAP7_75t_L g3783 ( 
.A(n_3734),
.B(n_3620),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3706),
.Y(n_3784)
);

INVx2_ASAP7_75t_L g3785 ( 
.A(n_3706),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3700),
.Y(n_3786)
);

BUFx2_ASAP7_75t_L g3787 ( 
.A(n_3698),
.Y(n_3787)
);

AND2x4_ASAP7_75t_L g3788 ( 
.A(n_3692),
.B(n_3574),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3706),
.Y(n_3789)
);

AND2x2_ASAP7_75t_L g3790 ( 
.A(n_3734),
.B(n_3770),
.Y(n_3790)
);

BUFx3_ASAP7_75t_L g3791 ( 
.A(n_3658),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3767),
.Y(n_3792)
);

BUFx10_ASAP7_75t_L g3793 ( 
.A(n_3658),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3767),
.Y(n_3794)
);

OR2x2_ASAP7_75t_L g3795 ( 
.A(n_3763),
.B(n_3613),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3765),
.B(n_3614),
.Y(n_3796)
);

BUFx4f_ASAP7_75t_L g3797 ( 
.A(n_3658),
.Y(n_3797)
);

BUFx6f_ASAP7_75t_L g3798 ( 
.A(n_3658),
.Y(n_3798)
);

HB1xp67_ASAP7_75t_L g3799 ( 
.A(n_3755),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3751),
.Y(n_3800)
);

AND2x4_ASAP7_75t_L g3801 ( 
.A(n_3692),
.B(n_3574),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3700),
.Y(n_3802)
);

INVx2_ASAP7_75t_SL g3803 ( 
.A(n_3698),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3666),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3667),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3671),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_3770),
.B(n_3594),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3659),
.A2(n_3542),
.B(n_3649),
.Y(n_3808)
);

AO21x2_ASAP7_75t_L g3809 ( 
.A1(n_3716),
.A2(n_3490),
.B(n_3596),
.Y(n_3809)
);

BUFx2_ASAP7_75t_L g3810 ( 
.A(n_3749),
.Y(n_3810)
);

INVx3_ASAP7_75t_L g3811 ( 
.A(n_3672),
.Y(n_3811)
);

OAI21x1_ASAP7_75t_L g3812 ( 
.A1(n_3728),
.A2(n_3511),
.B(n_3630),
.Y(n_3812)
);

INVx3_ASAP7_75t_L g3813 ( 
.A(n_3672),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3673),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3751),
.Y(n_3815)
);

HB1xp67_ASAP7_75t_L g3816 ( 
.A(n_3757),
.Y(n_3816)
);

INVx3_ASAP7_75t_L g3817 ( 
.A(n_3672),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3674),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3678),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3665),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3679),
.Y(n_3821)
);

INVx2_ASAP7_75t_L g3822 ( 
.A(n_3665),
.Y(n_3822)
);

INVx3_ASAP7_75t_L g3823 ( 
.A(n_3672),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3665),
.Y(n_3824)
);

BUFx3_ASAP7_75t_L g3825 ( 
.A(n_3658),
.Y(n_3825)
);

AOI21x1_ASAP7_75t_L g3826 ( 
.A1(n_3652),
.A2(n_3440),
.B(n_3300),
.Y(n_3826)
);

INVxp67_ASAP7_75t_L g3827 ( 
.A(n_3768),
.Y(n_3827)
);

INVx3_ASAP7_75t_L g3828 ( 
.A(n_3672),
.Y(n_3828)
);

OA21x2_ASAP7_75t_L g3829 ( 
.A1(n_3716),
.A2(n_3643),
.B(n_3564),
.Y(n_3829)
);

HB1xp67_ASAP7_75t_L g3830 ( 
.A(n_3653),
.Y(n_3830)
);

AO31x2_ASAP7_75t_L g3831 ( 
.A1(n_3713),
.A2(n_3455),
.A3(n_3453),
.B(n_3172),
.Y(n_3831)
);

INVx2_ASAP7_75t_SL g3832 ( 
.A(n_3749),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3713),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3770),
.B(n_3622),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3680),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3685),
.Y(n_3836)
);

CKINVDCx6p67_ASAP7_75t_R g3837 ( 
.A(n_3663),
.Y(n_3837)
);

BUFx2_ASAP7_75t_L g3838 ( 
.A(n_3749),
.Y(n_3838)
);

OA21x2_ASAP7_75t_L g3839 ( 
.A1(n_3652),
.A2(n_3661),
.B(n_3728),
.Y(n_3839)
);

OAI21x1_ASAP7_75t_L g3840 ( 
.A1(n_3756),
.A2(n_3504),
.B(n_3324),
.Y(n_3840)
);

OAI21x1_ASAP7_75t_L g3841 ( 
.A1(n_3756),
.A2(n_3504),
.B(n_3324),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3715),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3715),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3650),
.Y(n_3844)
);

AO21x2_ASAP7_75t_L g3845 ( 
.A1(n_3708),
.A2(n_3538),
.B(n_3600),
.Y(n_3845)
);

AO21x2_ASAP7_75t_L g3846 ( 
.A1(n_3670),
.A2(n_3573),
.B(n_3606),
.Y(n_3846)
);

HB1xp67_ASAP7_75t_L g3847 ( 
.A(n_3684),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3688),
.Y(n_3848)
);

OAI21x1_ASAP7_75t_L g3849 ( 
.A1(n_3772),
.A2(n_3335),
.B(n_3338),
.Y(n_3849)
);

OA21x2_ASAP7_75t_L g3850 ( 
.A1(n_3738),
.A2(n_3616),
.B(n_3648),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3650),
.Y(n_3851)
);

HB1xp67_ASAP7_75t_L g3852 ( 
.A(n_3684),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3709),
.Y(n_3853)
);

OA21x2_ASAP7_75t_L g3854 ( 
.A1(n_3740),
.A2(n_3737),
.B(n_3733),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3714),
.Y(n_3855)
);

HB1xp67_ASAP7_75t_L g3856 ( 
.A(n_3654),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3717),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3664),
.Y(n_3858)
);

BUFx3_ASAP7_75t_L g3859 ( 
.A(n_3663),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3772),
.B(n_3631),
.Y(n_3860)
);

BUFx3_ASAP7_75t_L g3861 ( 
.A(n_3695),
.Y(n_3861)
);

NOR2xp33_ASAP7_75t_L g3862 ( 
.A(n_3695),
.B(n_3749),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3719),
.Y(n_3863)
);

BUFx2_ASAP7_75t_L g3864 ( 
.A(n_3749),
.Y(n_3864)
);

BUFx2_ASAP7_75t_L g3865 ( 
.A(n_3743),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3772),
.B(n_3575),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3664),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3677),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3677),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3683),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3725),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3657),
.Y(n_3872)
);

OR2x6_ASAP7_75t_L g3873 ( 
.A(n_3692),
.B(n_3723),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3681),
.Y(n_3874)
);

OA21x2_ASAP7_75t_L g3875 ( 
.A1(n_3689),
.A2(n_3581),
.B(n_3572),
.Y(n_3875)
);

AO21x2_ASAP7_75t_L g3876 ( 
.A1(n_3694),
.A2(n_3149),
.B(n_3166),
.Y(n_3876)
);

OR2x2_ASAP7_75t_L g3877 ( 
.A(n_3676),
.B(n_3662),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3681),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3676),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3689),
.Y(n_3880)
);

OR2x2_ASAP7_75t_L g3881 ( 
.A(n_3703),
.B(n_3619),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3691),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3701),
.B(n_3556),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3691),
.Y(n_3884)
);

INVx3_ASAP7_75t_L g3885 ( 
.A(n_3686),
.Y(n_3885)
);

AO21x2_ASAP7_75t_L g3886 ( 
.A1(n_3694),
.A2(n_3235),
.B(n_3459),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3742),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3697),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3747),
.Y(n_3889)
);

BUFx2_ASAP7_75t_L g3890 ( 
.A(n_3743),
.Y(n_3890)
);

AND2x4_ASAP7_75t_L g3891 ( 
.A(n_3692),
.B(n_3632),
.Y(n_3891)
);

HB1xp67_ASAP7_75t_L g3892 ( 
.A(n_3703),
.Y(n_3892)
);

AND2x2_ASAP7_75t_L g3893 ( 
.A(n_3721),
.B(n_3559),
.Y(n_3893)
);

HB1xp67_ASAP7_75t_L g3894 ( 
.A(n_3760),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3750),
.Y(n_3895)
);

INVx3_ASAP7_75t_L g3896 ( 
.A(n_3686),
.Y(n_3896)
);

AND2x2_ASAP7_75t_L g3897 ( 
.A(n_3721),
.B(n_3546),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3697),
.Y(n_3898)
);

CKINVDCx5p33_ASAP7_75t_R g3899 ( 
.A(n_3837),
.Y(n_3899)
);

AND2x4_ASAP7_75t_L g3900 ( 
.A(n_3803),
.B(n_3702),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_3787),
.B(n_3768),
.Y(n_3901)
);

AND2x4_ASAP7_75t_L g3902 ( 
.A(n_3803),
.B(n_3702),
.Y(n_3902)
);

OAI211xp5_ASAP7_75t_L g3903 ( 
.A1(n_3799),
.A2(n_3682),
.B(n_3669),
.C(n_3702),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3787),
.B(n_3656),
.Y(n_3904)
);

AND2x4_ASAP7_75t_L g3905 ( 
.A(n_3803),
.B(n_3774),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3865),
.Y(n_3906)
);

INVx3_ASAP7_75t_L g3907 ( 
.A(n_3798),
.Y(n_3907)
);

A2O1A1Ixp33_ASAP7_75t_L g3908 ( 
.A1(n_3800),
.A2(n_3642),
.B(n_3759),
.C(n_3735),
.Y(n_3908)
);

AO21x2_ASAP7_75t_L g3909 ( 
.A1(n_3820),
.A2(n_3748),
.B(n_3739),
.Y(n_3909)
);

AO32x2_ASAP7_75t_L g3910 ( 
.A1(n_3832),
.A2(n_3745),
.A3(n_3722),
.B1(n_3696),
.B2(n_3746),
.Y(n_3910)
);

O2A1O1Ixp33_ASAP7_75t_L g3911 ( 
.A1(n_3809),
.A2(n_3687),
.B(n_3752),
.C(n_3642),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3891),
.B(n_3656),
.Y(n_3912)
);

AND2x4_ASAP7_75t_L g3913 ( 
.A(n_3891),
.B(n_3883),
.Y(n_3913)
);

OAI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3795),
.A2(n_3730),
.B1(n_3718),
.B2(n_3774),
.Y(n_3914)
);

O2A1O1Ixp33_ASAP7_75t_L g3915 ( 
.A1(n_3809),
.A2(n_3745),
.B(n_3722),
.C(n_3771),
.Y(n_3915)
);

OR2x2_ASAP7_75t_L g3916 ( 
.A(n_3795),
.B(n_3655),
.Y(n_3916)
);

BUFx3_ASAP7_75t_L g3917 ( 
.A(n_3861),
.Y(n_3917)
);

NOR2x1_ASAP7_75t_SL g3918 ( 
.A(n_3873),
.B(n_3686),
.Y(n_3918)
);

OAI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_3826),
.A2(n_3617),
.B(n_3732),
.Y(n_3919)
);

A2O1A1Ixp33_ASAP7_75t_L g3920 ( 
.A1(n_3800),
.A2(n_3705),
.B(n_3579),
.C(n_3651),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3776),
.Y(n_3921)
);

AND2x4_ASAP7_75t_L g3922 ( 
.A(n_3891),
.B(n_3771),
.Y(n_3922)
);

A2O1A1Ixp33_ASAP7_75t_L g3923 ( 
.A1(n_3800),
.A2(n_3705),
.B(n_3651),
.C(n_3601),
.Y(n_3923)
);

BUFx6f_ASAP7_75t_L g3924 ( 
.A(n_3861),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3891),
.B(n_3656),
.Y(n_3925)
);

NOR2xp33_ASAP7_75t_L g3926 ( 
.A(n_3861),
.B(n_3704),
.Y(n_3926)
);

CKINVDCx20_ASAP7_75t_R g3927 ( 
.A(n_3837),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3776),
.Y(n_3928)
);

OR2x2_ASAP7_75t_L g3929 ( 
.A(n_3796),
.B(n_3732),
.Y(n_3929)
);

AND2x2_ASAP7_75t_L g3930 ( 
.A(n_3897),
.B(n_3696),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3865),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3778),
.Y(n_3932)
);

BUFx2_ASAP7_75t_L g3933 ( 
.A(n_3890),
.Y(n_3933)
);

NOR2x1_ASAP7_75t_R g3934 ( 
.A(n_3859),
.B(n_3724),
.Y(n_3934)
);

AND2x2_ASAP7_75t_L g3935 ( 
.A(n_3897),
.B(n_3696),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3778),
.Y(n_3936)
);

HB1xp67_ASAP7_75t_L g3937 ( 
.A(n_3892),
.Y(n_3937)
);

NOR2x1_ASAP7_75t_SL g3938 ( 
.A(n_3873),
.B(n_3686),
.Y(n_3938)
);

OR2x2_ASAP7_75t_L g3939 ( 
.A(n_3796),
.B(n_3739),
.Y(n_3939)
);

AO21x2_ASAP7_75t_L g3940 ( 
.A1(n_3820),
.A2(n_3758),
.B(n_3764),
.Y(n_3940)
);

OAI22xp5_ASAP7_75t_L g3941 ( 
.A1(n_3829),
.A2(n_3718),
.B1(n_3758),
.B2(n_3555),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3883),
.B(n_3693),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3893),
.B(n_3693),
.Y(n_3943)
);

INVxp33_ASAP7_75t_SL g3944 ( 
.A(n_3862),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3845),
.B(n_3720),
.Y(n_3945)
);

A2O1A1Ixp33_ASAP7_75t_L g3946 ( 
.A1(n_3815),
.A2(n_3668),
.B(n_3741),
.C(n_3769),
.Y(n_3946)
);

INVx3_ASAP7_75t_L g3947 ( 
.A(n_3798),
.Y(n_3947)
);

OAI22xp5_ASAP7_75t_SL g3948 ( 
.A1(n_3798),
.A2(n_3718),
.B1(n_3724),
.B2(n_3621),
.Y(n_3948)
);

HB1xp67_ASAP7_75t_L g3949 ( 
.A(n_3892),
.Y(n_3949)
);

NOR2xp33_ASAP7_75t_L g3950 ( 
.A(n_3837),
.B(n_3718),
.Y(n_3950)
);

BUFx6f_ASAP7_75t_L g3951 ( 
.A(n_3798),
.Y(n_3951)
);

AND2x2_ASAP7_75t_SL g3952 ( 
.A(n_3829),
.B(n_3775),
.Y(n_3952)
);

OR2x2_ASAP7_75t_L g3953 ( 
.A(n_3877),
.B(n_3760),
.Y(n_3953)
);

HB1xp67_ASAP7_75t_L g3954 ( 
.A(n_3777),
.Y(n_3954)
);

OR2x2_ASAP7_75t_L g3955 ( 
.A(n_3877),
.B(n_3761),
.Y(n_3955)
);

NOR2xp33_ASAP7_75t_L g3956 ( 
.A(n_3859),
.B(n_3798),
.Y(n_3956)
);

OAI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3826),
.A2(n_3761),
.B(n_3675),
.Y(n_3957)
);

AOI221xp5_ASAP7_75t_L g3958 ( 
.A1(n_3792),
.A2(n_3637),
.B1(n_3729),
.B2(n_3699),
.C(n_3711),
.Y(n_3958)
);

AND2x4_ASAP7_75t_L g3959 ( 
.A(n_3893),
.B(n_3727),
.Y(n_3959)
);

AO21x2_ASAP7_75t_L g3960 ( 
.A1(n_3820),
.A2(n_3764),
.B(n_3769),
.Y(n_3960)
);

OAI22xp5_ASAP7_75t_L g3961 ( 
.A1(n_3829),
.A2(n_3555),
.B1(n_3754),
.B2(n_3753),
.Y(n_3961)
);

NOR2x1_ASAP7_75t_SL g3962 ( 
.A(n_3873),
.B(n_3686),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3777),
.B(n_3693),
.Y(n_3963)
);

CKINVDCx6p67_ASAP7_75t_R g3964 ( 
.A(n_3859),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3845),
.B(n_3720),
.Y(n_3965)
);

A2O1A1Ixp33_ASAP7_75t_L g3966 ( 
.A1(n_3815),
.A2(n_3741),
.B(n_3727),
.C(n_3736),
.Y(n_3966)
);

INVxp67_ASAP7_75t_L g3967 ( 
.A(n_3890),
.Y(n_3967)
);

AO21x1_ASAP7_75t_L g3968 ( 
.A1(n_3815),
.A2(n_3675),
.B(n_3475),
.Y(n_3968)
);

OAI22xp5_ASAP7_75t_L g3969 ( 
.A1(n_3829),
.A2(n_3555),
.B1(n_3724),
.B2(n_3736),
.Y(n_3969)
);

AO21x2_ASAP7_75t_L g3970 ( 
.A1(n_3822),
.A2(n_3699),
.B(n_3729),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3845),
.B(n_3799),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3777),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3866),
.B(n_3775),
.Y(n_3973)
);

AND2x4_ASAP7_75t_L g3974 ( 
.A(n_3832),
.B(n_3775),
.Y(n_3974)
);

HB1xp67_ASAP7_75t_L g3975 ( 
.A(n_3830),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3811),
.Y(n_3976)
);

OR2x2_ASAP7_75t_L g3977 ( 
.A(n_3816),
.B(n_3775),
.Y(n_3977)
);

AND2x2_ASAP7_75t_L g3978 ( 
.A(n_3866),
.B(n_3775),
.Y(n_3978)
);

AOI211xp5_ASAP7_75t_L g3979 ( 
.A1(n_3816),
.A2(n_3794),
.B(n_3792),
.C(n_3822),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3807),
.B(n_3724),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_3811),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3855),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3845),
.B(n_3744),
.Y(n_3983)
);

AOI221xp5_ASAP7_75t_L g3984 ( 
.A1(n_3792),
.A2(n_3711),
.B1(n_3712),
.B2(n_3489),
.C(n_3762),
.Y(n_3984)
);

AND2x2_ASAP7_75t_SL g3985 ( 
.A(n_3829),
.B(n_3731),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3809),
.A2(n_3723),
.B1(n_3712),
.B2(n_3766),
.Y(n_3986)
);

A2O1A1Ixp33_ASAP7_75t_L g3987 ( 
.A1(n_3794),
.A2(n_3726),
.B(n_3731),
.C(n_3762),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3807),
.B(n_3731),
.Y(n_3988)
);

NOR2xp33_ASAP7_75t_L g3989 ( 
.A(n_3798),
.B(n_3726),
.Y(n_3989)
);

INVx5_ASAP7_75t_L g3990 ( 
.A(n_3798),
.Y(n_3990)
);

OR2x6_ASAP7_75t_L g3991 ( 
.A(n_3832),
.B(n_3723),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3786),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3855),
.Y(n_3993)
);

NOR2xp33_ASAP7_75t_L g3994 ( 
.A(n_3791),
.B(n_3660),
.Y(n_3994)
);

OAI221xp5_ASAP7_75t_SL g3995 ( 
.A1(n_3794),
.A2(n_3723),
.B1(n_3766),
.B2(n_3744),
.C(n_3710),
.Y(n_3995)
);

INVxp67_ASAP7_75t_L g3996 ( 
.A(n_3810),
.Y(n_3996)
);

AOI221xp5_ASAP7_75t_L g3997 ( 
.A1(n_3809),
.A2(n_3352),
.B1(n_3196),
.B2(n_3710),
.C(n_3773),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3834),
.B(n_3773),
.Y(n_3998)
);

OAI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3839),
.A2(n_3824),
.B(n_3822),
.Y(n_3999)
);

A2O1A1Ixp33_ASAP7_75t_L g4000 ( 
.A1(n_3824),
.A2(n_3509),
.B(n_3501),
.C(n_3498),
.Y(n_4000)
);

AOI221xp5_ASAP7_75t_L g4001 ( 
.A1(n_3824),
.A2(n_3785),
.B1(n_3784),
.B2(n_3789),
.C(n_3779),
.Y(n_4001)
);

AND2x4_ASAP7_75t_L g4002 ( 
.A(n_3827),
.B(n_3484),
.Y(n_4002)
);

AOI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3846),
.A2(n_3766),
.B1(n_3633),
.B2(n_3604),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_L g4004 ( 
.A1(n_3846),
.A2(n_3780),
.B1(n_3850),
.B2(n_3875),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3786),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3834),
.B(n_3507),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3860),
.B(n_3508),
.Y(n_4007)
);

BUFx2_ASAP7_75t_L g4008 ( 
.A(n_3791),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3847),
.B(n_3592),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3860),
.B(n_3508),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3782),
.B(n_3783),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3811),
.Y(n_4012)
);

AO32x2_ASAP7_75t_L g4013 ( 
.A1(n_3846),
.A2(n_3766),
.A3(n_3633),
.B1(n_3604),
.B2(n_3592),
.Y(n_4013)
);

INVx5_ASAP7_75t_SL g4014 ( 
.A(n_3797),
.Y(n_4014)
);

O2A1O1Ixp33_ASAP7_75t_SL g4015 ( 
.A1(n_3827),
.A2(n_3633),
.B(n_3604),
.C(n_3592),
.Y(n_4015)
);

INVx1_ASAP7_75t_SL g4016 ( 
.A(n_3791),
.Y(n_4016)
);

AOI21xp5_ASAP7_75t_SL g4017 ( 
.A1(n_3839),
.A2(n_3509),
.B(n_3501),
.Y(n_4017)
);

AND2x4_ASAP7_75t_L g4018 ( 
.A(n_3922),
.B(n_3810),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3922),
.B(n_3838),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3937),
.Y(n_4020)
);

AND2x2_ASAP7_75t_L g4021 ( 
.A(n_3901),
.B(n_3838),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3949),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3970),
.Y(n_4023)
);

NAND4xp25_ASAP7_75t_L g4024 ( 
.A(n_3915),
.B(n_3864),
.C(n_3825),
.D(n_3790),
.Y(n_4024)
);

AOI22xp33_ASAP7_75t_L g4025 ( 
.A1(n_3952),
.A2(n_3846),
.B1(n_3780),
.B2(n_3850),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3975),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3921),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_3913),
.B(n_3864),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3933),
.B(n_3854),
.Y(n_4029)
);

INVx4_ASAP7_75t_L g4030 ( 
.A(n_3924),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3913),
.B(n_3825),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3921),
.Y(n_4032)
);

AND2x4_ASAP7_75t_L g4033 ( 
.A(n_3900),
.B(n_3825),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3900),
.B(n_3790),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3928),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3928),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3902),
.B(n_3793),
.Y(n_4037)
);

NAND2x1p5_ASAP7_75t_L g4038 ( 
.A(n_3990),
.B(n_3797),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3970),
.Y(n_4039)
);

HB1xp67_ASAP7_75t_L g4040 ( 
.A(n_3999),
.Y(n_4040)
);

OAI22xp5_ASAP7_75t_L g4041 ( 
.A1(n_3903),
.A2(n_3839),
.B1(n_3854),
.B2(n_3847),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3932),
.Y(n_4042)
);

AOI22xp33_ASAP7_75t_L g4043 ( 
.A1(n_3985),
.A2(n_3780),
.B1(n_3850),
.B2(n_3854),
.Y(n_4043)
);

OR2x2_ASAP7_75t_L g4044 ( 
.A(n_3954),
.B(n_3916),
.Y(n_4044)
);

OR2x2_ASAP7_75t_L g4045 ( 
.A(n_3972),
.B(n_3779),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_L g4046 ( 
.A(n_3971),
.B(n_3854),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3967),
.B(n_3854),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3906),
.B(n_3852),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3960),
.Y(n_4049)
);

INVx1_ASAP7_75t_SL g4050 ( 
.A(n_3927),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3902),
.B(n_3793),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3932),
.Y(n_4052)
);

NAND2x1p5_ASAP7_75t_L g4053 ( 
.A(n_3990),
.B(n_3797),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3973),
.B(n_3793),
.Y(n_4054)
);

OR2x2_ASAP7_75t_L g4055 ( 
.A(n_3953),
.B(n_3779),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3931),
.B(n_3852),
.Y(n_4056)
);

AO21x2_ASAP7_75t_L g4057 ( 
.A1(n_3946),
.A2(n_3785),
.B(n_3784),
.Y(n_4057)
);

AND2x4_ASAP7_75t_L g4058 ( 
.A(n_3905),
.B(n_3781),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3978),
.B(n_3793),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_3988),
.B(n_3797),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3960),
.Y(n_4061)
);

OAI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_3911),
.A2(n_3839),
.B(n_3780),
.Y(n_4062)
);

INVx2_ASAP7_75t_SL g4063 ( 
.A(n_3917),
.Y(n_4063)
);

AND2x4_ASAP7_75t_L g4064 ( 
.A(n_3905),
.B(n_3781),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3940),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3980),
.B(n_3782),
.Y(n_4066)
);

INVxp67_ASAP7_75t_L g4067 ( 
.A(n_3926),
.Y(n_4067)
);

BUFx3_ASAP7_75t_L g4068 ( 
.A(n_3924),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_3942),
.B(n_3783),
.Y(n_4069)
);

HB1xp67_ASAP7_75t_L g4070 ( 
.A(n_3979),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_3940),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3951),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3936),
.Y(n_4073)
);

OR2x2_ASAP7_75t_L g4074 ( 
.A(n_3955),
.B(n_3781),
.Y(n_4074)
);

INVx2_ASAP7_75t_SL g4075 ( 
.A(n_3924),
.Y(n_4075)
);

OR2x2_ASAP7_75t_L g4076 ( 
.A(n_3929),
.B(n_3879),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3936),
.Y(n_4077)
);

INVx3_ASAP7_75t_L g4078 ( 
.A(n_3951),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3943),
.B(n_3839),
.Y(n_4079)
);

INVxp67_ASAP7_75t_L g4080 ( 
.A(n_3956),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3951),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_3963),
.B(n_3856),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3992),
.Y(n_4083)
);

BUFx2_ASAP7_75t_L g4084 ( 
.A(n_3899),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_4008),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_4013),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3992),
.Y(n_4087)
);

AOI22xp5_ASAP7_75t_L g4088 ( 
.A1(n_4004),
.A2(n_3850),
.B1(n_3780),
.B2(n_3875),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_4013),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_4016),
.B(n_3879),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4005),
.Y(n_4091)
);

BUFx2_ASAP7_75t_L g4092 ( 
.A(n_3964),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_4005),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_4011),
.B(n_3894),
.Y(n_4094)
);

OAI222xp33_ASAP7_75t_L g4095 ( 
.A1(n_3986),
.A2(n_3873),
.B1(n_3784),
.B2(n_3785),
.C1(n_3789),
.C2(n_3894),
.Y(n_4095)
);

BUFx2_ASAP7_75t_L g4096 ( 
.A(n_3959),
.Y(n_4096)
);

OR2x2_ASAP7_75t_L g4097 ( 
.A(n_3939),
.B(n_3830),
.Y(n_4097)
);

OR2x2_ASAP7_75t_L g4098 ( 
.A(n_3983),
.B(n_3887),
.Y(n_4098)
);

AND2x4_ASAP7_75t_L g4099 ( 
.A(n_3959),
.B(n_3788),
.Y(n_4099)
);

BUFx6f_ASAP7_75t_L g4100 ( 
.A(n_3990),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3982),
.Y(n_4101)
);

OR2x2_ASAP7_75t_L g4102 ( 
.A(n_3977),
.B(n_3887),
.Y(n_4102)
);

HB1xp67_ASAP7_75t_L g4103 ( 
.A(n_3996),
.Y(n_4103)
);

AND2x2_ASAP7_75t_L g4104 ( 
.A(n_3930),
.B(n_3856),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3993),
.Y(n_4105)
);

OR2x2_ASAP7_75t_L g4106 ( 
.A(n_4009),
.B(n_3889),
.Y(n_4106)
);

BUFx3_ASAP7_75t_L g4107 ( 
.A(n_3944),
.Y(n_4107)
);

HB1xp67_ASAP7_75t_L g4108 ( 
.A(n_3904),
.Y(n_4108)
);

CKINVDCx20_ASAP7_75t_R g4109 ( 
.A(n_3994),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_4001),
.Y(n_4110)
);

AOI221xp5_ASAP7_75t_L g4111 ( 
.A1(n_4070),
.A2(n_3920),
.B1(n_3958),
.B2(n_3923),
.C(n_3969),
.Y(n_4111)
);

NOR2xp33_ASAP7_75t_L g4112 ( 
.A(n_4107),
.B(n_3934),
.Y(n_4112)
);

AOI22xp33_ASAP7_75t_L g4113 ( 
.A1(n_4040),
.A2(n_3968),
.B1(n_3909),
.B2(n_3850),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_4050),
.B(n_3935),
.Y(n_4114)
);

NAND3xp33_ASAP7_75t_L g4115 ( 
.A(n_4070),
.B(n_3966),
.C(n_3908),
.Y(n_4115)
);

AOI21xp5_ASAP7_75t_SL g4116 ( 
.A1(n_4041),
.A2(n_3914),
.B(n_3987),
.Y(n_4116)
);

OAI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_4043),
.A2(n_4025),
.B1(n_4040),
.B2(n_4017),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_4058),
.B(n_3945),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_4033),
.B(n_3788),
.Y(n_4119)
);

OAI221xp5_ASAP7_75t_SL g4120 ( 
.A1(n_4043),
.A2(n_4003),
.B1(n_3965),
.B2(n_3984),
.C(n_3997),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_L g4121 ( 
.A1(n_4025),
.A2(n_3909),
.B1(n_3961),
.B2(n_3941),
.Y(n_4121)
);

OAI21xp5_ASAP7_75t_SL g4122 ( 
.A1(n_4024),
.A2(n_3957),
.B(n_3950),
.Y(n_4122)
);

NOR2xp33_ASAP7_75t_L g4123 ( 
.A(n_4107),
.B(n_3989),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_4058),
.B(n_3889),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_4058),
.B(n_3895),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_4064),
.B(n_3895),
.Y(n_4126)
);

NAND3xp33_ASAP7_75t_L g4127 ( 
.A(n_4062),
.B(n_3789),
.C(n_3919),
.Y(n_4127)
);

AND2x2_ASAP7_75t_SL g4128 ( 
.A(n_4103),
.B(n_3974),
.Y(n_4128)
);

NOR3xp33_ASAP7_75t_L g4129 ( 
.A(n_4110),
.B(n_3995),
.C(n_3947),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_4096),
.B(n_4084),
.Y(n_4130)
);

NOR3xp33_ASAP7_75t_L g4131 ( 
.A(n_4046),
.B(n_3947),
.C(n_3907),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_4031),
.B(n_3912),
.Y(n_4132)
);

NAND3xp33_ASAP7_75t_L g4133 ( 
.A(n_4088),
.B(n_3981),
.C(n_3976),
.Y(n_4133)
);

NOR3xp33_ASAP7_75t_L g4134 ( 
.A(n_4047),
.B(n_3907),
.C(n_3872),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4064),
.B(n_3872),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_4064),
.B(n_3857),
.Y(n_4136)
);

OAI22xp5_ASAP7_75t_L g4137 ( 
.A1(n_4109),
.A2(n_4014),
.B1(n_3788),
.B2(n_3801),
.Y(n_4137)
);

NAND3xp33_ASAP7_75t_L g4138 ( 
.A(n_4067),
.B(n_4012),
.C(n_3974),
.Y(n_4138)
);

INVx4_ASAP7_75t_L g4139 ( 
.A(n_4030),
.Y(n_4139)
);

NOR3xp33_ASAP7_75t_L g4140 ( 
.A(n_4029),
.B(n_3948),
.C(n_3813),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_4094),
.B(n_3857),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_4094),
.B(n_4108),
.Y(n_4142)
);

AOI22xp33_ASAP7_75t_SL g4143 ( 
.A1(n_4079),
.A2(n_3918),
.B1(n_3938),
.B2(n_3962),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_4108),
.B(n_3863),
.Y(n_4144)
);

NOR2xp33_ASAP7_75t_L g4145 ( 
.A(n_4109),
.B(n_4030),
.Y(n_4145)
);

NOR3xp33_ASAP7_75t_L g4146 ( 
.A(n_4030),
.B(n_3813),
.C(n_3811),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_L g4147 ( 
.A1(n_4049),
.A2(n_4061),
.B1(n_4071),
.B2(n_4065),
.Y(n_4147)
);

NAND3xp33_ASAP7_75t_L g4148 ( 
.A(n_4103),
.B(n_3925),
.C(n_3817),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_4031),
.B(n_4028),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_4028),
.B(n_3998),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_SL g4151 ( 
.A(n_4033),
.B(n_3788),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4092),
.B(n_4014),
.Y(n_4152)
);

NAND3xp33_ASAP7_75t_L g4153 ( 
.A(n_4080),
.B(n_3817),
.C(n_3813),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_4085),
.B(n_3863),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_4019),
.B(n_4007),
.Y(n_4155)
);

NOR2xp33_ASAP7_75t_L g4156 ( 
.A(n_4068),
.B(n_3801),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4085),
.B(n_3871),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_SL g4158 ( 
.A(n_4033),
.B(n_3801),
.Y(n_4158)
);

NAND3xp33_ASAP7_75t_L g4159 ( 
.A(n_4063),
.B(n_3817),
.C(n_3813),
.Y(n_4159)
);

NAND3xp33_ASAP7_75t_L g4160 ( 
.A(n_4063),
.B(n_3823),
.C(n_3817),
.Y(n_4160)
);

OA21x2_ASAP7_75t_L g4161 ( 
.A1(n_4023),
.A2(n_3812),
.B(n_3808),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_4019),
.B(n_4010),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_4082),
.B(n_3871),
.Y(n_4163)
);

OAI221xp5_ASAP7_75t_SL g4164 ( 
.A1(n_4079),
.A2(n_4000),
.B1(n_3873),
.B2(n_3991),
.C(n_3910),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_4128),
.Y(n_4165)
);

HB1xp67_ASAP7_75t_L g4166 ( 
.A(n_4130),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_4128),
.B(n_4104),
.Y(n_4167)
);

INVxp67_ASAP7_75t_L g4168 ( 
.A(n_4145),
.Y(n_4168)
);

AND2x2_ASAP7_75t_SL g4169 ( 
.A(n_4152),
.B(n_4113),
.Y(n_4169)
);

NOR2xp33_ASAP7_75t_L g4170 ( 
.A(n_4139),
.B(n_4068),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4141),
.Y(n_4171)
);

INVx4_ASAP7_75t_L g4172 ( 
.A(n_4139),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_4149),
.B(n_4034),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4142),
.Y(n_4174)
);

INVx2_ASAP7_75t_L g4175 ( 
.A(n_4161),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_4161),
.Y(n_4176)
);

AND2x4_ASAP7_75t_L g4177 ( 
.A(n_4150),
.B(n_4018),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_4118),
.B(n_4104),
.Y(n_4178)
);

OR2x6_ASAP7_75t_L g4179 ( 
.A(n_4116),
.B(n_4075),
.Y(n_4179)
);

OAI211xp5_ASAP7_75t_SL g4180 ( 
.A1(n_4122),
.A2(n_4056),
.B(n_4048),
.C(n_4044),
.Y(n_4180)
);

OR2x2_ASAP7_75t_L g4181 ( 
.A(n_4163),
.B(n_4076),
.Y(n_4181)
);

AOI22xp33_ASAP7_75t_L g4182 ( 
.A1(n_4127),
.A2(n_4071),
.B1(n_4049),
.B2(n_4061),
.Y(n_4182)
);

NAND3xp33_ASAP7_75t_L g4183 ( 
.A(n_4113),
.B(n_4026),
.C(n_4022),
.Y(n_4183)
);

OAI33xp33_ASAP7_75t_L g4184 ( 
.A1(n_4117),
.A2(n_4115),
.A3(n_4135),
.B1(n_4020),
.B2(n_4144),
.B3(n_4133),
.Y(n_4184)
);

HB1xp67_ASAP7_75t_L g4185 ( 
.A(n_4114),
.Y(n_4185)
);

AND2x2_ASAP7_75t_L g4186 ( 
.A(n_4132),
.B(n_4034),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_4124),
.B(n_4075),
.Y(n_4187)
);

INVx4_ASAP7_75t_L g4188 ( 
.A(n_4155),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_SL g4189 ( 
.A(n_4123),
.B(n_4018),
.Y(n_4189)
);

NOR2x1p5_ASAP7_75t_L g4190 ( 
.A(n_4138),
.B(n_4090),
.Y(n_4190)
);

AND2x4_ASAP7_75t_L g4191 ( 
.A(n_4162),
.B(n_4018),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4154),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_4156),
.B(n_4021),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4157),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4125),
.B(n_4097),
.Y(n_4195)
);

INVx5_ASAP7_75t_L g4196 ( 
.A(n_4112),
.Y(n_4196)
);

OAI211xp5_ASAP7_75t_L g4197 ( 
.A1(n_4111),
.A2(n_4098),
.B(n_4051),
.C(n_4037),
.Y(n_4197)
);

OAI31xp33_ASAP7_75t_SL g4198 ( 
.A1(n_4143),
.A2(n_4099),
.A3(n_4051),
.B(n_4037),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4136),
.Y(n_4199)
);

OR2x2_ASAP7_75t_L g4200 ( 
.A(n_4126),
.B(n_4055),
.Y(n_4200)
);

INVx2_ASAP7_75t_L g4201 ( 
.A(n_4119),
.Y(n_4201)
);

AND2x4_ASAP7_75t_L g4202 ( 
.A(n_4151),
.B(n_4099),
.Y(n_4202)
);

INVx2_ASAP7_75t_L g4203 ( 
.A(n_4158),
.Y(n_4203)
);

BUFx2_ASAP7_75t_L g4204 ( 
.A(n_4137),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4129),
.B(n_4021),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_4140),
.B(n_4099),
.Y(n_4206)
);

NOR2x1_ASAP7_75t_SL g4207 ( 
.A(n_4148),
.B(n_4100),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4147),
.Y(n_4208)
);

INVx2_ASAP7_75t_L g4209 ( 
.A(n_4159),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_4140),
.B(n_4069),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_4160),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_4153),
.Y(n_4212)
);

AND2x2_ASAP7_75t_L g4213 ( 
.A(n_4129),
.B(n_4069),
.Y(n_4213)
);

OR2x2_ASAP7_75t_L g4214 ( 
.A(n_4134),
.B(n_4074),
.Y(n_4214)
);

NAND4xp25_ASAP7_75t_L g4215 ( 
.A(n_4134),
.B(n_4060),
.C(n_4054),
.D(n_4066),
.Y(n_4215)
);

INVx1_ASAP7_75t_SL g4216 ( 
.A(n_4164),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4185),
.Y(n_4217)
);

INVx2_ASAP7_75t_L g4218 ( 
.A(n_4169),
.Y(n_4218)
);

HB1xp67_ASAP7_75t_L g4219 ( 
.A(n_4166),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4173),
.B(n_4121),
.Y(n_4220)
);

AND2x4_ASAP7_75t_L g4221 ( 
.A(n_4177),
.B(n_4054),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4175),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_4169),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4175),
.Y(n_4224)
);

OR2x2_ASAP7_75t_L g4225 ( 
.A(n_4200),
.B(n_4045),
.Y(n_4225)
);

OAI22xp5_ASAP7_75t_L g4226 ( 
.A1(n_4179),
.A2(n_4120),
.B1(n_4106),
.B2(n_3801),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_4200),
.B(n_4102),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_4176),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_4176),
.Y(n_4229)
);

AND2x4_ASAP7_75t_L g4230 ( 
.A(n_4177),
.B(n_4191),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_4173),
.B(n_4072),
.Y(n_4231)
);

AND2x2_ASAP7_75t_L g4232 ( 
.A(n_4179),
.B(n_4059),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4181),
.Y(n_4233)
);

OR2x2_ASAP7_75t_L g4234 ( 
.A(n_4214),
.B(n_4101),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4188),
.B(n_4213),
.Y(n_4235)
);

INVx1_ASAP7_75t_SL g4236 ( 
.A(n_4193),
.Y(n_4236)
);

INVx3_ASAP7_75t_L g4237 ( 
.A(n_4179),
.Y(n_4237)
);

INVx2_ASAP7_75t_SL g4238 ( 
.A(n_4177),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_4188),
.B(n_3910),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4186),
.Y(n_4240)
);

OAI221xp5_ASAP7_75t_L g4241 ( 
.A1(n_4179),
.A2(n_4086),
.B1(n_4089),
.B2(n_4065),
.C(n_4131),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4186),
.Y(n_4242)
);

INVxp67_ASAP7_75t_L g4243 ( 
.A(n_4189),
.Y(n_4243)
);

HB1xp67_ASAP7_75t_L g4244 ( 
.A(n_4183),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4165),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4165),
.Y(n_4246)
);

AND2x2_ASAP7_75t_L g4247 ( 
.A(n_4188),
.B(n_3910),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4213),
.B(n_4072),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_4193),
.B(n_4081),
.Y(n_4249)
);

INVx4_ASAP7_75t_L g4250 ( 
.A(n_4172),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4210),
.B(n_4081),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_4210),
.B(n_4105),
.Y(n_4252)
);

OAI21xp33_ASAP7_75t_L g4253 ( 
.A1(n_4205),
.A2(n_4146),
.B(n_4131),
.Y(n_4253)
);

AND2x2_ASAP7_75t_L g4254 ( 
.A(n_4191),
.B(n_4038),
.Y(n_4254)
);

OR2x2_ASAP7_75t_L g4255 ( 
.A(n_4178),
.B(n_4027),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_4230),
.Y(n_4256)
);

INVxp67_ASAP7_75t_SL g4257 ( 
.A(n_4244),
.Y(n_4257)
);

OAI22xp5_ASAP7_75t_L g4258 ( 
.A1(n_4244),
.A2(n_4167),
.B1(n_4190),
.B2(n_4212),
.Y(n_4258)
);

OR2x2_ASAP7_75t_L g4259 ( 
.A(n_4236),
.B(n_4195),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4219),
.Y(n_4260)
);

AND2x4_ASAP7_75t_L g4261 ( 
.A(n_4230),
.B(n_4191),
.Y(n_4261)
);

INVx2_ASAP7_75t_L g4262 ( 
.A(n_4230),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_4238),
.B(n_4201),
.Y(n_4263)
);

OR2x2_ASAP7_75t_L g4264 ( 
.A(n_4227),
.B(n_4174),
.Y(n_4264)
);

OR2x2_ASAP7_75t_L g4265 ( 
.A(n_4240),
.B(n_4201),
.Y(n_4265)
);

OR2x2_ASAP7_75t_L g4266 ( 
.A(n_4242),
.B(n_4203),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4219),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4225),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4218),
.B(n_4192),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4228),
.Y(n_4270)
);

OR2x2_ASAP7_75t_L g4271 ( 
.A(n_4235),
.B(n_4203),
.Y(n_4271)
);

INVx2_ASAP7_75t_L g4272 ( 
.A(n_4237),
.Y(n_4272)
);

INVxp33_ASAP7_75t_L g4273 ( 
.A(n_4232),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_4237),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_R g4275 ( 
.A(n_4238),
.B(n_4196),
.Y(n_4275)
);

INVx2_ASAP7_75t_SL g4276 ( 
.A(n_4221),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4228),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_4218),
.B(n_4194),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4223),
.B(n_4171),
.Y(n_4279)
);

NAND2x1p5_ASAP7_75t_L g4280 ( 
.A(n_4237),
.B(n_4196),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4249),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_4261),
.B(n_4239),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_4261),
.B(n_4221),
.Y(n_4283)
);

OAI22xp33_ASAP7_75t_L g4284 ( 
.A1(n_4257),
.A2(n_4223),
.B1(n_4220),
.B2(n_4216),
.Y(n_4284)
);

AOI22xp5_ASAP7_75t_L g4285 ( 
.A1(n_4258),
.A2(n_4184),
.B1(n_4208),
.B2(n_4247),
.Y(n_4285)
);

INVx2_ASAP7_75t_SL g4286 ( 
.A(n_4276),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4281),
.B(n_4221),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_4265),
.Y(n_4288)
);

INVxp67_ASAP7_75t_SL g4289 ( 
.A(n_4263),
.Y(n_4289)
);

AOI22xp5_ASAP7_75t_L g4290 ( 
.A1(n_4258),
.A2(n_4247),
.B1(n_4245),
.B2(n_4246),
.Y(n_4290)
);

OAI211xp5_ASAP7_75t_L g4291 ( 
.A1(n_4275),
.A2(n_4253),
.B(n_4198),
.C(n_4243),
.Y(n_4291)
);

AND2x4_ASAP7_75t_L g4292 ( 
.A(n_4256),
.B(n_4196),
.Y(n_4292)
);

INVx2_ASAP7_75t_SL g4293 ( 
.A(n_4262),
.Y(n_4293)
);

AND2x4_ASAP7_75t_L g4294 ( 
.A(n_4268),
.B(n_4196),
.Y(n_4294)
);

AOI321xp33_ASAP7_75t_L g4295 ( 
.A1(n_4272),
.A2(n_4226),
.A3(n_4241),
.B1(n_4182),
.B2(n_4248),
.C(n_4206),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4266),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_4259),
.Y(n_4297)
);

OR2x2_ASAP7_75t_L g4298 ( 
.A(n_4264),
.B(n_4271),
.Y(n_4298)
);

HB1xp67_ASAP7_75t_L g4299 ( 
.A(n_4280),
.Y(n_4299)
);

AND2x4_ASAP7_75t_L g4300 ( 
.A(n_4260),
.B(n_4196),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4270),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4298),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4283),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4292),
.B(n_4249),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4287),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_4289),
.Y(n_4306)
);

OAI22x1_ASAP7_75t_L g4307 ( 
.A1(n_4285),
.A2(n_4204),
.B1(n_4168),
.B2(n_4217),
.Y(n_4307)
);

NOR2x1_ASAP7_75t_R g4308 ( 
.A(n_4286),
.B(n_4172),
.Y(n_4308)
);

INVx2_ASAP7_75t_SL g4309 ( 
.A(n_4294),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4282),
.Y(n_4310)
);

XNOR2x1_ASAP7_75t_L g4311 ( 
.A(n_4284),
.B(n_4280),
.Y(n_4311)
);

XNOR2xp5_ASAP7_75t_L g4312 ( 
.A(n_4290),
.B(n_4232),
.Y(n_4312)
);

AO22x2_ASAP7_75t_L g4313 ( 
.A1(n_4291),
.A2(n_4277),
.B1(n_4222),
.B2(n_4229),
.Y(n_4313)
);

XOR2x2_ASAP7_75t_L g4314 ( 
.A(n_4297),
.B(n_4251),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4288),
.Y(n_4315)
);

NOR2x1_ASAP7_75t_L g4316 ( 
.A(n_4296),
.B(n_4172),
.Y(n_4316)
);

INVx1_ASAP7_75t_SL g4317 ( 
.A(n_4294),
.Y(n_4317)
);

XOR2x2_ASAP7_75t_L g4318 ( 
.A(n_4293),
.B(n_4279),
.Y(n_4318)
);

CKINVDCx16_ASAP7_75t_R g4319 ( 
.A(n_4312),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4318),
.Y(n_4320)
);

INVx2_ASAP7_75t_L g4321 ( 
.A(n_4302),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4302),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4304),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4314),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_4303),
.B(n_4202),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4313),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4313),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_4305),
.B(n_4273),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_L g4329 ( 
.A(n_4317),
.B(n_4267),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4316),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_4319),
.B(n_4292),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_4325),
.Y(n_4332)
);

NAND3xp33_ASAP7_75t_L g4333 ( 
.A(n_4326),
.B(n_4311),
.C(n_4299),
.Y(n_4333)
);

INVx1_ASAP7_75t_SL g4334 ( 
.A(n_4329),
.Y(n_4334)
);

OAI22xp33_ASAP7_75t_L g4335 ( 
.A1(n_4327),
.A2(n_4322),
.B1(n_4321),
.B2(n_4278),
.Y(n_4335)
);

AO21x1_ASAP7_75t_L g4336 ( 
.A1(n_4329),
.A2(n_4250),
.B(n_4300),
.Y(n_4336)
);

INVx2_ASAP7_75t_L g4337 ( 
.A(n_4320),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4328),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_SL g4339 ( 
.A1(n_4331),
.A2(n_4300),
.B(n_4307),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4334),
.B(n_4274),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_L g4341 ( 
.A(n_4332),
.B(n_4206),
.Y(n_4341)
);

OAI22xp5_ASAP7_75t_L g4342 ( 
.A1(n_4338),
.A2(n_4328),
.B1(n_4279),
.B2(n_4315),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4336),
.Y(n_4343)
);

AOI21xp33_ASAP7_75t_L g4344 ( 
.A1(n_4335),
.A2(n_4324),
.B(n_4278),
.Y(n_4344)
);

AOI221xp5_ASAP7_75t_L g4345 ( 
.A1(n_4337),
.A2(n_4224),
.B1(n_4269),
.B2(n_4301),
.C(n_4182),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4333),
.Y(n_4346)
);

NOR2xp33_ASAP7_75t_L g4347 ( 
.A(n_4334),
.B(n_4310),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4334),
.B(n_4254),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_SL g4349 ( 
.A1(n_4334),
.A2(n_4269),
.B(n_4306),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4334),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_4334),
.B(n_4202),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4348),
.B(n_4233),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4351),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4345),
.B(n_4252),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4350),
.B(n_4254),
.Y(n_4355)
);

INVx2_ASAP7_75t_L g4356 ( 
.A(n_4340),
.Y(n_4356)
);

AND2x4_ASAP7_75t_L g4357 ( 
.A(n_4346),
.B(n_4309),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4341),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4347),
.B(n_4202),
.Y(n_4359)
);

INVx1_ASAP7_75t_SL g4360 ( 
.A(n_4343),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4342),
.Y(n_4361)
);

BUFx12f_ASAP7_75t_L g4362 ( 
.A(n_4339),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4344),
.B(n_4170),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4349),
.B(n_4170),
.Y(n_4364)
);

AND2x2_ASAP7_75t_L g4365 ( 
.A(n_4348),
.B(n_4231),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_4348),
.B(n_4323),
.Y(n_4366)
);

AOI222xp33_ASAP7_75t_L g4367 ( 
.A1(n_4345),
.A2(n_4147),
.B1(n_4023),
.B2(n_4039),
.C1(n_4180),
.C2(n_4295),
.Y(n_4367)
);

AND2x2_ASAP7_75t_L g4368 ( 
.A(n_4348),
.B(n_4207),
.Y(n_4368)
);

INVx2_ASAP7_75t_SL g4369 ( 
.A(n_4348),
.Y(n_4369)
);

NOR2xp33_ASAP7_75t_L g4370 ( 
.A(n_4351),
.B(n_4234),
.Y(n_4370)
);

AOI22xp5_ASAP7_75t_L g4371 ( 
.A1(n_4345),
.A2(n_4330),
.B1(n_4199),
.B2(n_4250),
.Y(n_4371)
);

INVx2_ASAP7_75t_SL g4372 ( 
.A(n_4348),
.Y(n_4372)
);

OR2x2_ASAP7_75t_L g4373 ( 
.A(n_4351),
.B(n_4215),
.Y(n_4373)
);

INVx1_ASAP7_75t_SL g4374 ( 
.A(n_4359),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4365),
.Y(n_4375)
);

AOI221xp5_ASAP7_75t_L g4376 ( 
.A1(n_4360),
.A2(n_4250),
.B1(n_4197),
.B2(n_4187),
.C(n_4212),
.Y(n_4376)
);

INVx2_ASAP7_75t_SL g4377 ( 
.A(n_4362),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4368),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4352),
.Y(n_4379)
);

AOI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_4356),
.A2(n_4211),
.B1(n_4209),
.B2(n_4255),
.Y(n_4380)
);

NAND4xp75_ASAP7_75t_L g4381 ( 
.A(n_4366),
.B(n_4308),
.C(n_4211),
.D(n_4209),
.Y(n_4381)
);

OAI322xp33_ASAP7_75t_L g4382 ( 
.A1(n_4360),
.A2(n_4039),
.A3(n_4086),
.B1(n_4089),
.B2(n_4093),
.C1(n_4091),
.C2(n_4036),
.Y(n_4382)
);

AOI22xp5_ASAP7_75t_L g4383 ( 
.A1(n_4370),
.A2(n_4078),
.B1(n_4057),
.B2(n_4146),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_4352),
.Y(n_4384)
);

NAND2x1_ASAP7_75t_SL g4385 ( 
.A(n_4355),
.B(n_4078),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4357),
.Y(n_4386)
);

AO22x2_ASAP7_75t_L g4387 ( 
.A1(n_4369),
.A2(n_4372),
.B1(n_4357),
.B2(n_4353),
.Y(n_4387)
);

INVx1_ASAP7_75t_SL g4388 ( 
.A(n_4364),
.Y(n_4388)
);

AND4x1_ASAP7_75t_L g4389 ( 
.A(n_4363),
.B(n_4073),
.C(n_4042),
.D(n_4087),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4373),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4361),
.Y(n_4391)
);

AO22x2_ASAP7_75t_L g4392 ( 
.A1(n_4358),
.A2(n_4032),
.B1(n_4052),
.B2(n_4083),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_4354),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4371),
.Y(n_4394)
);

AOI221xp5_ASAP7_75t_L g4395 ( 
.A1(n_4371),
.A2(n_4095),
.B1(n_4057),
.B2(n_4078),
.C(n_4077),
.Y(n_4395)
);

AOI22xp5_ASAP7_75t_L g4396 ( 
.A1(n_4367),
.A2(n_4100),
.B1(n_4035),
.B2(n_4038),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4367),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4365),
.Y(n_4398)
);

AOI22xp5_ASAP7_75t_L g4399 ( 
.A1(n_4356),
.A2(n_4100),
.B1(n_4053),
.B2(n_3828),
.Y(n_4399)
);

NOR3xp33_ASAP7_75t_L g4400 ( 
.A(n_4377),
.B(n_3828),
.C(n_3823),
.Y(n_4400)
);

NOR2xp33_ASAP7_75t_L g4401 ( 
.A(n_4374),
.B(n_4100),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4387),
.B(n_4053),
.Y(n_4402)
);

INVx2_ASAP7_75t_L g4403 ( 
.A(n_4387),
.Y(n_4403)
);

NOR3xp33_ASAP7_75t_L g4404 ( 
.A(n_4386),
.B(n_3828),
.C(n_3823),
.Y(n_4404)
);

NOR3xp33_ASAP7_75t_L g4405 ( 
.A(n_4375),
.B(n_3828),
.C(n_3823),
.Y(n_4405)
);

AND3x1_ASAP7_75t_L g4406 ( 
.A(n_4376),
.B(n_3896),
.C(n_3885),
.Y(n_4406)
);

INVxp67_ASAP7_75t_L g4407 ( 
.A(n_4381),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4385),
.Y(n_4408)
);

NOR3x1_ASAP7_75t_L g4409 ( 
.A(n_4379),
.B(n_3812),
.C(n_3840),
.Y(n_4409)
);

NOR3xp33_ASAP7_75t_L g4410 ( 
.A(n_4398),
.B(n_3896),
.C(n_3885),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_4388),
.B(n_3833),
.Y(n_4411)
);

INVxp67_ASAP7_75t_L g4412 ( 
.A(n_4384),
.Y(n_4412)
);

AND4x1_ASAP7_75t_L g4413 ( 
.A(n_4394),
.B(n_4013),
.C(n_4015),
.D(n_4006),
.Y(n_4413)
);

O2A1O1Ixp33_ASAP7_75t_SL g4414 ( 
.A1(n_4390),
.A2(n_3885),
.B(n_3896),
.C(n_3881),
.Y(n_4414)
);

AOI21xp5_ASAP7_75t_L g4415 ( 
.A1(n_4378),
.A2(n_3842),
.B(n_3833),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4392),
.Y(n_4416)
);

AND2x2_ASAP7_75t_L g4417 ( 
.A(n_4380),
.B(n_4391),
.Y(n_4417)
);

NOR3xp33_ASAP7_75t_L g4418 ( 
.A(n_4397),
.B(n_3896),
.C(n_3885),
.Y(n_4418)
);

XNOR2xp5_ASAP7_75t_L g4419 ( 
.A(n_4389),
.B(n_3873),
.Y(n_4419)
);

AOI21xp33_ASAP7_75t_L g4420 ( 
.A1(n_4393),
.A2(n_3844),
.B(n_3851),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4396),
.B(n_3833),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_SL g4422 ( 
.A(n_4399),
.B(n_4002),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4392),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_4402),
.B(n_4383),
.Y(n_4424)
);

NOR2x1p5_ASAP7_75t_SL g4425 ( 
.A(n_4403),
.B(n_4382),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_4408),
.B(n_4395),
.Y(n_4426)
);

NAND4xp25_ASAP7_75t_L g4427 ( 
.A(n_4401),
.B(n_4417),
.C(n_4407),
.D(n_4412),
.Y(n_4427)
);

AOI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_4423),
.A2(n_3842),
.B(n_3843),
.Y(n_4428)
);

NOR4xp25_ASAP7_75t_L g4429 ( 
.A(n_4416),
.B(n_3843),
.C(n_3842),
.D(n_3802),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_4413),
.B(n_4002),
.Y(n_4430)
);

AND3x2_ASAP7_75t_L g4431 ( 
.A(n_4418),
.B(n_3843),
.C(n_3802),
.Y(n_4431)
);

NOR2xp33_ASAP7_75t_L g4432 ( 
.A(n_4419),
.B(n_3844),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4411),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_SL g4434 ( 
.A(n_4406),
.B(n_3804),
.Y(n_4434)
);

AOI21xp5_ASAP7_75t_L g4435 ( 
.A1(n_4421),
.A2(n_3819),
.B(n_3821),
.Y(n_4435)
);

AO22x2_ASAP7_75t_L g4436 ( 
.A1(n_4422),
.A2(n_3868),
.B1(n_3898),
.B2(n_3888),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_4415),
.B(n_3844),
.Y(n_4437)
);

NAND4xp75_ASAP7_75t_L g4438 ( 
.A(n_4420),
.B(n_3875),
.C(n_3819),
.D(n_3821),
.Y(n_4438)
);

NOR3xp33_ASAP7_75t_L g4439 ( 
.A(n_4400),
.B(n_4404),
.C(n_4410),
.Y(n_4439)
);

AND2x2_ASAP7_75t_L g4440 ( 
.A(n_4405),
.B(n_3991),
.Y(n_4440)
);

OAI211xp5_ASAP7_75t_SL g4441 ( 
.A1(n_4424),
.A2(n_4414),
.B(n_4409),
.C(n_3881),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4425),
.B(n_3851),
.Y(n_4442)
);

NOR2xp33_ASAP7_75t_L g4443 ( 
.A(n_4427),
.B(n_3851),
.Y(n_4443)
);

NAND2xp33_ASAP7_75t_SL g4444 ( 
.A(n_4426),
.B(n_3804),
.Y(n_4444)
);

NOR2x1_ASAP7_75t_L g4445 ( 
.A(n_4433),
.B(n_3805),
.Y(n_4445)
);

NAND3x1_ASAP7_75t_L g4446 ( 
.A(n_4439),
.B(n_3853),
.C(n_3805),
.Y(n_4446)
);

AND2x2_ASAP7_75t_L g4447 ( 
.A(n_4430),
.B(n_3806),
.Y(n_4447)
);

NAND3xp33_ASAP7_75t_SL g4448 ( 
.A(n_4432),
.B(n_3898),
.C(n_3888),
.Y(n_4448)
);

NAND4xp25_ASAP7_75t_L g4449 ( 
.A(n_4428),
.B(n_3170),
.C(n_3888),
.D(n_3884),
.Y(n_4449)
);

AOI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_4434),
.A2(n_3898),
.B(n_3858),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_4440),
.B(n_3858),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_4436),
.Y(n_4452)
);

NAND3xp33_ASAP7_75t_SL g4453 ( 
.A(n_4429),
.B(n_3884),
.C(n_3882),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4431),
.B(n_3858),
.Y(n_4454)
);

NOR4xp25_ASAP7_75t_L g4455 ( 
.A(n_4437),
.B(n_3853),
.C(n_3814),
.D(n_3818),
.Y(n_4455)
);

AOI322xp5_ASAP7_75t_L g4456 ( 
.A1(n_4443),
.A2(n_4436),
.A3(n_4438),
.B1(n_4435),
.B2(n_3806),
.C1(n_3814),
.C2(n_3818),
.Y(n_4456)
);

AOI222xp33_ASAP7_75t_L g4457 ( 
.A1(n_4442),
.A2(n_3868),
.B1(n_3884),
.B2(n_3882),
.C1(n_3874),
.C2(n_3869),
.Y(n_4457)
);

OAI221xp5_ASAP7_75t_L g4458 ( 
.A1(n_4441),
.A2(n_3836),
.B1(n_3835),
.B2(n_3848),
.C(n_3870),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4454),
.Y(n_4459)
);

O2A1O1Ixp33_ASAP7_75t_L g4460 ( 
.A1(n_4452),
.A2(n_3835),
.B(n_3836),
.C(n_3848),
.Y(n_4460)
);

OAI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_4446),
.A2(n_3870),
.B1(n_3882),
.B2(n_3874),
.Y(n_4461)
);

AOI211xp5_ASAP7_75t_L g4462 ( 
.A1(n_4444),
.A2(n_3812),
.B(n_3841),
.C(n_3840),
.Y(n_4462)
);

BUFx8_ASAP7_75t_SL g4463 ( 
.A(n_4447),
.Y(n_4463)
);

AOI22xp5_ASAP7_75t_L g4464 ( 
.A1(n_4445),
.A2(n_4451),
.B1(n_4453),
.B2(n_4448),
.Y(n_4464)
);

NOR3xp33_ASAP7_75t_L g4465 ( 
.A(n_4450),
.B(n_3808),
.C(n_3840),
.Y(n_4465)
);

OAI21xp33_ASAP7_75t_L g4466 ( 
.A1(n_4455),
.A2(n_3808),
.B(n_3869),
.Y(n_4466)
);

XOR2x2_ASAP7_75t_L g4467 ( 
.A(n_4449),
.B(n_3875),
.Y(n_4467)
);

AOI221xp5_ASAP7_75t_L g4468 ( 
.A1(n_4441),
.A2(n_3867),
.B1(n_3868),
.B2(n_3874),
.C(n_3869),
.Y(n_4468)
);

OAI311xp33_ASAP7_75t_L g4469 ( 
.A1(n_4442),
.A2(n_3880),
.A3(n_3878),
.B1(n_3875),
.C1(n_3841),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_4442),
.B(n_3867),
.Y(n_4470)
);

OAI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_4446),
.A2(n_3867),
.B1(n_3880),
.B2(n_3878),
.Y(n_4471)
);

AOI221xp5_ASAP7_75t_L g4472 ( 
.A1(n_4441),
.A2(n_3886),
.B1(n_3498),
.B2(n_3500),
.C(n_3876),
.Y(n_4472)
);

NAND2x1_ASAP7_75t_L g4473 ( 
.A(n_4445),
.B(n_3500),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_4463),
.B(n_3886),
.Y(n_4474)
);

INVx2_ASAP7_75t_L g4475 ( 
.A(n_4473),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4470),
.Y(n_4476)
);

NOR2x1_ASAP7_75t_L g4477 ( 
.A(n_4459),
.B(n_3886),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4464),
.B(n_3886),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4467),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4471),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4460),
.Y(n_4481)
);

BUFx4f_ASAP7_75t_SL g4482 ( 
.A(n_4456),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4461),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4458),
.Y(n_4484)
);

AOI22xp33_ASAP7_75t_L g4485 ( 
.A1(n_4466),
.A2(n_3841),
.B1(n_3849),
.B2(n_3876),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4468),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_4457),
.B(n_3831),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_SL g4488 ( 
.A(n_4472),
.B(n_3849),
.Y(n_4488)
);

AOI22xp5_ASAP7_75t_L g4489 ( 
.A1(n_4465),
.A2(n_3849),
.B1(n_3876),
.B2(n_3303),
.Y(n_4489)
);

AOI22xp5_ASAP7_75t_L g4490 ( 
.A1(n_4462),
.A2(n_4469),
.B1(n_3876),
.B2(n_3303),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4475),
.Y(n_4491)
);

CKINVDCx5p33_ASAP7_75t_R g4492 ( 
.A(n_4479),
.Y(n_4492)
);

NAND3x1_ASAP7_75t_L g4493 ( 
.A(n_4481),
.B(n_288),
.C(n_291),
.Y(n_4493)
);

AND3x4_ASAP7_75t_L g4494 ( 
.A(n_4482),
.B(n_292),
.C(n_293),
.Y(n_4494)
);

NOR4xp25_ASAP7_75t_L g4495 ( 
.A(n_4476),
.B(n_294),
.C(n_295),
.D(n_298),
.Y(n_4495)
);

AOI211xp5_ASAP7_75t_L g4496 ( 
.A1(n_4486),
.A2(n_299),
.B(n_300),
.C(n_302),
.Y(n_4496)
);

OAI311xp33_ASAP7_75t_L g4497 ( 
.A1(n_4474),
.A2(n_311),
.A3(n_315),
.B1(n_316),
.C1(n_318),
.Y(n_4497)
);

AOI211xp5_ASAP7_75t_L g4498 ( 
.A1(n_4484),
.A2(n_320),
.B(n_321),
.C(n_324),
.Y(n_4498)
);

OR2x2_ASAP7_75t_L g4499 ( 
.A(n_4478),
.B(n_3831),
.Y(n_4499)
);

OAI221xp5_ASAP7_75t_L g4500 ( 
.A1(n_4483),
.A2(n_3258),
.B1(n_326),
.B2(n_327),
.C(n_328),
.Y(n_4500)
);

NAND4xp75_ASAP7_75t_L g4501 ( 
.A(n_4480),
.B(n_325),
.C(n_329),
.D(n_330),
.Y(n_4501)
);

AOI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_4491),
.A2(n_4488),
.B1(n_4487),
.B2(n_4490),
.Y(n_4502)
);

NAND2xp33_ASAP7_75t_SL g4503 ( 
.A(n_4494),
.B(n_4485),
.Y(n_4503)
);

NAND4xp75_ASAP7_75t_L g4504 ( 
.A(n_4492),
.B(n_4489),
.C(n_4477),
.D(n_335),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_4493),
.B(n_331),
.Y(n_4505)
);

NOR2x1_ASAP7_75t_L g4506 ( 
.A(n_4501),
.B(n_332),
.Y(n_4506)
);

NOR2xp33_ASAP7_75t_L g4507 ( 
.A(n_4497),
.B(n_336),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4507),
.B(n_4495),
.Y(n_4508)
);

INVx1_ASAP7_75t_SL g4509 ( 
.A(n_4503),
.Y(n_4509)
);

HB1xp67_ASAP7_75t_L g4510 ( 
.A(n_4502),
.Y(n_4510)
);

AO22x2_ASAP7_75t_L g4511 ( 
.A1(n_4509),
.A2(n_4508),
.B1(n_4504),
.B2(n_4505),
.Y(n_4511)
);

AO22x2_ASAP7_75t_L g4512 ( 
.A1(n_4510),
.A2(n_4506),
.B1(n_4498),
.B2(n_4496),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4511),
.Y(n_4513)
);

AOI22xp33_ASAP7_75t_L g4514 ( 
.A1(n_4513),
.A2(n_4512),
.B1(n_4499),
.B2(n_4500),
.Y(n_4514)
);

INVx3_ASAP7_75t_SL g4515 ( 
.A(n_4514),
.Y(n_4515)
);

OAI22x1_ASAP7_75t_L g4516 ( 
.A1(n_4515),
.A2(n_337),
.B1(n_342),
.B2(n_349),
.Y(n_4516)
);

XNOR2xp5_ASAP7_75t_L g4517 ( 
.A(n_4516),
.B(n_352),
.Y(n_4517)
);

NOR2xp33_ASAP7_75t_L g4518 ( 
.A(n_4517),
.B(n_354),
.Y(n_4518)
);

OAI22xp33_ASAP7_75t_L g4519 ( 
.A1(n_4518),
.A2(n_3221),
.B1(n_3258),
.B2(n_3398),
.Y(n_4519)
);

NAND3xp33_ASAP7_75t_L g4520 ( 
.A(n_4519),
.B(n_359),
.C(n_362),
.Y(n_4520)
);

AOI22xp5_ASAP7_75t_L g4521 ( 
.A1(n_4520),
.A2(n_3200),
.B1(n_3221),
.B2(n_3398),
.Y(n_4521)
);

OA21x2_ASAP7_75t_L g4522 ( 
.A1(n_4521),
.A2(n_364),
.B(n_366),
.Y(n_4522)
);

OAI221xp5_ASAP7_75t_R g4523 ( 
.A1(n_4522),
.A2(n_372),
.B1(n_374),
.B2(n_379),
.C(n_381),
.Y(n_4523)
);

AOI21xp5_ASAP7_75t_L g4524 ( 
.A1(n_4523),
.A2(n_384),
.B(n_389),
.Y(n_4524)
);

AOI211xp5_ASAP7_75t_L g4525 ( 
.A1(n_4524),
.A2(n_394),
.B(n_395),
.C(n_396),
.Y(n_4525)
);


endmodule