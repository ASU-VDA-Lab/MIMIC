module fake_jpeg_26058_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_44),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_33),
.B1(n_18),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_54),
.B1(n_60),
.B2(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_49),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_57),
.Y(n_68)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_33),
.B1(n_24),
.B2(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_62),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_56),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_33),
.B1(n_27),
.B2(n_30),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_34),
.B1(n_32),
.B2(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_21),
.B1(n_32),
.B2(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_71),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_25),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_35),
.B1(n_16),
.B2(n_19),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_86),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_78),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_76),
.B(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_36),
.B1(n_56),
.B2(n_29),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_35),
.B1(n_19),
.B2(n_28),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_80),
.A2(n_94),
.B1(n_99),
.B2(n_0),
.Y(n_129)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_25),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_92),
.B(n_93),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_20),
.B(n_26),
.C(n_31),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_106),
.B1(n_56),
.B2(n_46),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_26),
.B(n_31),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_20),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_54),
.B1(n_45),
.B2(n_28),
.Y(n_94)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_36),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_0),
.Y(n_128)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_101),
.Y(n_130)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_28),
.B1(n_23),
.B2(n_29),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_60),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_0),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_29),
.B1(n_23),
.B2(n_38),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_129),
.B1(n_95),
.B2(n_93),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_114),
.B1(n_121),
.B2(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_23),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_26),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_103),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_20),
.B1(n_8),
.B2(n_2),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_93),
.B1(n_103),
.B2(n_79),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_8),
.B1(n_14),
.B2(n_3),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_7),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_72),
.C(n_68),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_79),
.B(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_89),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_132),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_155),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_137),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_117),
.B1(n_118),
.B2(n_114),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_143),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_86),
.C(n_104),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_160),
.C(n_102),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_147),
.A2(n_152),
.B1(n_81),
.B2(n_123),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_151),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_164),
.B1(n_146),
.B2(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_120),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_73),
.Y(n_153)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_127),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_120),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_97),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_84),
.B1(n_76),
.B2(n_70),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_118),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_84),
.B1(n_73),
.B2(n_87),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_74),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_167),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_121),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_82),
.Y(n_165)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_105),
.B1(n_83),
.B2(n_77),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_169),
.A2(n_81),
.B1(n_158),
.B2(n_82),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_169),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_120),
.C(n_128),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_190),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_177),
.A2(n_178),
.B1(n_193),
.B2(n_151),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_124),
.B1(n_112),
.B2(n_108),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_122),
.B(n_109),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_162),
.B(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_189),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_147),
.A2(n_106),
.B1(n_122),
.B2(n_109),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_195),
.B1(n_139),
.B2(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_98),
.B1(n_134),
.B2(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_142),
.B(n_134),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_188),
.B1(n_192),
.B2(n_186),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_160),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_205),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_141),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_217),
.C(n_202),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_207),
.B1(n_219),
.B2(n_220),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_197),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_208),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_210),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_136),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_215),
.B(n_178),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_156),
.C(n_158),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_184),
.CI(n_170),
.CON(n_238),
.SN(n_238)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_222),
.A2(n_192),
.B1(n_186),
.B2(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_227),
.B1(n_222),
.B2(n_212),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_220),
.B1(n_210),
.B2(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_203),
.C(n_215),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_236),
.C(n_242),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_182),
.C(n_172),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_206),
.B(n_176),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_168),
.C(n_187),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_207),
.A2(n_184),
.B1(n_135),
.B2(n_1),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_1),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_205),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_247),
.B(n_257),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_258),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_237),
.Y(n_264)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_256),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_135),
.C(n_5),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_229),
.C(n_228),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_227),
.A2(n_135),
.B1(n_6),
.B2(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_225),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_258)
);

INVxp33_ASAP7_75t_SL g259 ( 
.A(n_241),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_236),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_249),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_233),
.B(n_224),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_250),
.B(n_243),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_240),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_234),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_249),
.C(n_252),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_278),
.C(n_282),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_235),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_232),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_251),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_234),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_247),
.B1(n_255),
.B2(n_257),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_280),
.A2(n_261),
.B1(n_270),
.B2(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_254),
.C(n_232),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_262),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_285),
.A2(n_292),
.B1(n_278),
.B2(n_274),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_263),
.C(n_272),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_267),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_242),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_296),
.B(n_297),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_291),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_286),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_281),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_295),
.B(n_289),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_303),
.A2(n_300),
.B1(n_302),
.B2(n_299),
.Y(n_304)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_10),
.B(n_13),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_13),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_15),
.B1(n_223),
.B2(n_204),
.Y(n_307)
);


endmodule