module fake_jpeg_841_n_109 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_17),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_37),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_32),
.B1(n_38),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_51),
.B1(n_44),
.B2(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_32),
.B1(n_38),
.B2(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_30),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_35),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_57),
.B1(n_35),
.B2(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_36),
.B1(n_44),
.B2(n_35),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_0),
.C(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_60),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_6),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_72),
.B(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_3),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_5),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_3),
.B(n_4),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_8),
.B(n_9),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_78),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_19),
.C(n_26),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_15),
.C(n_23),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_83),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_7),
.Y(n_83)
);

OAI22x1_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_20),
.B1(n_25),
.B2(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_27),
.C(n_22),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_11),
.B(n_16),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_94),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_85),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_99),
.C(n_90),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_87),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_88),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_97),
.B(n_93),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_106),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_95),
.B1(n_99),
.B2(n_101),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_93),
.Y(n_109)
);


endmodule