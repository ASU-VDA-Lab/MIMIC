module real_aes_7146_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
INVx1_ASAP7_75t_L g525 ( .A(n_1), .Y(n_525) );
INVx1_ASAP7_75t_L g147 ( .A(n_2), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_3), .A2(n_36), .B1(n_172), .B2(n_471), .Y(n_494) );
AOI21xp33_ASAP7_75t_L g179 ( .A1(n_4), .A2(n_163), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_5), .B(n_161), .Y(n_537) );
AND2x6_ASAP7_75t_L g140 ( .A(n_6), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_7), .A2(n_250), .B(n_251), .Y(n_249) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_8), .B(n_37), .Y(n_437) );
INVx1_ASAP7_75t_L g185 ( .A(n_9), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_10), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g132 ( .A(n_11), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_12), .B(n_153), .Y(n_480) );
INVx1_ASAP7_75t_L g256 ( .A(n_13), .Y(n_256) );
INVx1_ASAP7_75t_L g519 ( .A(n_14), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_15), .B(n_128), .Y(n_508) );
AO32x2_ASAP7_75t_L g492 ( .A1(n_16), .A2(n_127), .A3(n_161), .B1(n_473), .B2(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_17), .B(n_172), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_18), .B(n_168), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_19), .B(n_128), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_20), .A2(n_48), .B1(n_172), .B2(n_471), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_21), .B(n_163), .Y(n_213) );
OAI222xp33_ASAP7_75t_L g442 ( .A1(n_22), .A2(n_443), .B1(n_727), .B2(n_728), .C1(n_733), .C2(n_737), .Y(n_442) );
INVx1_ASAP7_75t_L g727 ( .A(n_22), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_23), .A2(n_73), .B1(n_153), .B2(n_172), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_24), .B(n_172), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_25), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_26), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_28), .B(n_158), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_29), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g200 ( .A(n_30), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_31), .B(n_158), .Y(n_464) );
INVx2_ASAP7_75t_L g138 ( .A(n_32), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_33), .B(n_172), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_34), .B(n_158), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_35), .A2(n_140), .B(n_143), .C(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_37), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g198 ( .A(n_38), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_39), .B(n_151), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_40), .B(n_172), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_41), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_42), .A2(n_83), .B1(n_220), .B2(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_43), .B(n_172), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_44), .B(n_172), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_45), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_46), .B(n_524), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_47), .B(n_163), .Y(n_244) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_49), .A2(n_59), .B1(n_153), .B2(n_172), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_50), .A2(n_143), .B1(n_153), .B2(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_51), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_52), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_53), .B(n_172), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_54), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_55), .B(n_172), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_56), .A2(n_171), .B(n_183), .C(n_184), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_57), .Y(n_233) );
INVx1_ASAP7_75t_L g181 ( .A(n_58), .Y(n_181) );
INVx1_ASAP7_75t_L g141 ( .A(n_60), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_61), .B(n_172), .Y(n_526) );
INVx1_ASAP7_75t_L g131 ( .A(n_62), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_63), .Y(n_115) );
AO32x2_ASAP7_75t_L g468 ( .A1(n_64), .A2(n_161), .A3(n_236), .B1(n_469), .B2(n_473), .Y(n_468) );
INVx1_ASAP7_75t_L g544 ( .A(n_65), .Y(n_544) );
INVx1_ASAP7_75t_L g459 ( .A(n_66), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_67), .A2(n_168), .B(n_169), .C(n_171), .Y(n_167) );
INVxp67_ASAP7_75t_L g170 ( .A(n_68), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_69), .B(n_153), .Y(n_460) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_71), .Y(n_203) );
INVx1_ASAP7_75t_L g226 ( .A(n_72), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_74), .A2(n_140), .B(n_143), .C(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_75), .B(n_471), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_76), .B(n_153), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_77), .B(n_148), .Y(n_216) );
INVx2_ASAP7_75t_L g129 ( .A(n_78), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_79), .B(n_168), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_80), .B(n_153), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_81), .A2(n_140), .B(n_143), .C(n_146), .Y(n_142) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_82), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g434 ( .A(n_82), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g447 ( .A(n_82), .B(n_436), .Y(n_447) );
INVx2_ASAP7_75t_L g726 ( .A(n_82), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_84), .A2(n_98), .B1(n_153), .B2(n_154), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_85), .A2(n_118), .B1(n_119), .B2(n_432), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_85), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_86), .B(n_158), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_87), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_88), .A2(n_100), .B1(n_111), .B2(n_738), .Y(n_99) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_89), .A2(n_140), .B(n_143), .C(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_90), .Y(n_246) );
INVx1_ASAP7_75t_L g166 ( .A(n_91), .Y(n_166) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_92), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_93), .B(n_148), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_94), .B(n_153), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_95), .B(n_161), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_97), .A2(n_163), .B(n_164), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx5_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_103), .Y(n_739) );
OR2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g436 ( .A(n_107), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_116), .B(n_441), .Y(n_111) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_112), .A2(n_438), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_433), .B(n_438), .Y(n_116) );
INVx1_ASAP7_75t_L g432 ( .A(n_119), .Y(n_432) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_120), .A2(n_445), .B1(n_448), .B2(n_723), .Y(n_444) );
INVx1_ASAP7_75t_L g731 ( .A(n_120), .Y(n_731) );
NAND2x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_348), .Y(n_120) );
NOR5xp2_ASAP7_75t_L g121 ( .A(n_122), .B(n_271), .C(n_303), .D(n_318), .E(n_335), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_187), .B(n_208), .C(n_259), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_159), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_124), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_124), .B(n_323), .Y(n_386) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_125), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_125), .B(n_205), .Y(n_272) );
AND2x2_ASAP7_75t_L g313 ( .A(n_125), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_125), .B(n_282), .Y(n_317) );
OR2x2_ASAP7_75t_L g354 ( .A(n_125), .B(n_193), .Y(n_354) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g192 ( .A(n_126), .B(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g262 ( .A(n_126), .Y(n_262) );
OR2x2_ASAP7_75t_L g425 ( .A(n_126), .B(n_265), .Y(n_425) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_133), .B(n_155), .Y(n_126) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_127), .A2(n_194), .B(n_202), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_127), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g221 ( .A(n_127), .Y(n_221) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_129), .B(n_130), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B(n_142), .Y(n_133) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_135), .A2(n_173), .B1(n_195), .B2(n_201), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_135), .A2(n_226), .B(n_227), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
AND2x4_ASAP7_75t_L g163 ( .A(n_136), .B(n_140), .Y(n_163) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g524 ( .A(n_137), .Y(n_524) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx3_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_139), .Y(n_151) );
INVx1_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
INVx4_ASAP7_75t_SL g173 ( .A(n_140), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_140), .A2(n_458), .B(n_461), .Y(n_457) );
BUFx3_ASAP7_75t_L g473 ( .A(n_140), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_140), .A2(n_478), .B(n_482), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_140), .A2(n_518), .B(n_522), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_140), .A2(n_531), .B(n_534), .Y(n_530) );
INVx5_ASAP7_75t_L g165 ( .A(n_143), .Y(n_165) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
BUFx3_ASAP7_75t_L g220 ( .A(n_144), .Y(n_220) );
INVx1_ASAP7_75t_L g471 ( .A(n_144), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_150), .C(n_152), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_SL g458 ( .A1(n_148), .A2(n_171), .B(n_459), .C(n_460), .Y(n_458) );
INVx2_ASAP7_75t_L g495 ( .A(n_148), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_148), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_148), .A2(n_541), .B(n_542), .Y(n_540) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_149), .B(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_149), .B(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_149), .A2(n_151), .B1(n_470), .B2(n_472), .Y(n_469) );
INVx2_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx4_ASAP7_75t_L g242 ( .A(n_151), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_151), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_151), .A2(n_495), .B1(n_511), .B2(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_152), .A2(n_519), .B(n_520), .C(n_521), .Y(n_518) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_157), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_157), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_158), .A2(n_249), .B(n_258), .Y(n_248) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_158), .A2(n_457), .B(n_464), .Y(n_456) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_158), .A2(n_477), .B(n_485), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_159), .A2(n_328), .B1(n_329), .B2(n_332), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_159), .B(n_262), .Y(n_411) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_177), .Y(n_159) );
AND2x2_ASAP7_75t_L g207 ( .A(n_160), .B(n_193), .Y(n_207) );
AND2x2_ASAP7_75t_L g264 ( .A(n_160), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g269 ( .A(n_160), .Y(n_269) );
INVx3_ASAP7_75t_L g282 ( .A(n_160), .Y(n_282) );
OR2x2_ASAP7_75t_L g302 ( .A(n_160), .B(n_265), .Y(n_302) );
AND2x2_ASAP7_75t_L g321 ( .A(n_160), .B(n_178), .Y(n_321) );
BUFx2_ASAP7_75t_L g353 ( .A(n_160), .Y(n_353) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_174), .Y(n_160) );
INVx4_ASAP7_75t_L g176 ( .A(n_161), .Y(n_176) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_161), .A2(n_530), .B(n_537), .Y(n_529) );
BUFx2_ASAP7_75t_L g250 ( .A(n_163), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_173), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_165), .A2(n_173), .B(n_181), .C(n_182), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_165), .A2(n_173), .B(n_252), .C(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g481 ( .A(n_168), .Y(n_481) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_172), .Y(n_243) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_175), .A2(n_179), .B(n_186), .Y(n_178) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_176), .B(n_223), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_176), .B(n_473), .C(n_510), .Y(n_509) );
AO21x1_ASAP7_75t_L g599 ( .A1(n_176), .A2(n_510), .B(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g268 ( .A(n_177), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
BUFx2_ASAP7_75t_L g191 ( .A(n_178), .Y(n_191) );
INVx2_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
OR2x2_ASAP7_75t_L g284 ( .A(n_178), .B(n_265), .Y(n_284) );
AND2x2_ASAP7_75t_L g314 ( .A(n_178), .B(n_193), .Y(n_314) );
AND2x2_ASAP7_75t_L g331 ( .A(n_178), .B(n_262), .Y(n_331) );
AND2x2_ASAP7_75t_L g371 ( .A(n_178), .B(n_282), .Y(n_371) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_178), .B(n_207), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_183), .A2(n_483), .B(n_484), .Y(n_482) );
O2A1O1Ixp5_ASAP7_75t_L g543 ( .A1(n_183), .A2(n_523), .B(n_544), .C(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp33_ASAP7_75t_SL g188 ( .A(n_189), .B(n_204), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_192), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_190), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
OAI21xp33_ASAP7_75t_L g345 ( .A1(n_191), .A2(n_207), .B(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_191), .B(n_193), .Y(n_401) );
AND2x2_ASAP7_75t_L g337 ( .A(n_192), .B(n_338), .Y(n_337) );
INVx3_ASAP7_75t_L g265 ( .A(n_193), .Y(n_265) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_193), .Y(n_363) );
OAI22xp5_ASAP7_75t_SL g196 ( .A1(n_197), .A2(n_198), .B1(n_199), .B2(n_200), .Y(n_196) );
INVx2_ASAP7_75t_L g199 ( .A(n_197), .Y(n_199) );
INVx4_ASAP7_75t_L g254 ( .A(n_197), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_204), .B(n_262), .Y(n_430) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_205), .A2(n_373), .B1(n_374), .B2(n_379), .Y(n_372) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
AND2x2_ASAP7_75t_L g263 ( .A(n_206), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g301 ( .A(n_206), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g338 ( .A(n_206), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_207), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g392 ( .A(n_207), .Y(n_392) );
CKINVDCx16_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_234), .Y(n_209) );
INVx4_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
AND2x2_ASAP7_75t_L g356 ( .A(n_210), .B(n_323), .Y(n_356) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_224), .Y(n_210) );
INVx3_ASAP7_75t_L g275 ( .A(n_211), .Y(n_275) );
AND2x2_ASAP7_75t_L g289 ( .A(n_211), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g293 ( .A(n_211), .Y(n_293) );
INVx2_ASAP7_75t_L g307 ( .A(n_211), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_211), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g364 ( .A(n_211), .B(n_359), .Y(n_364) );
AND2x2_ASAP7_75t_L g429 ( .A(n_211), .B(n_399), .Y(n_429) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
AOI21xp5_ASAP7_75t_SL g212 ( .A1(n_213), .A2(n_214), .B(n_221), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_218), .A2(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g257 ( .A(n_220), .Y(n_257) );
INVx1_ASAP7_75t_L g231 ( .A(n_221), .Y(n_231) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_221), .A2(n_517), .B(n_527), .Y(n_516) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_221), .A2(n_539), .B(n_546), .Y(n_538) );
AND2x2_ASAP7_75t_L g270 ( .A(n_224), .B(n_248), .Y(n_270) );
INVx2_ASAP7_75t_L g290 ( .A(n_224), .Y(n_290) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_231), .B(n_232), .Y(n_224) );
INVx1_ASAP7_75t_L g295 ( .A(n_234), .Y(n_295) );
AND2x2_ASAP7_75t_L g341 ( .A(n_234), .B(n_289), .Y(n_341) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_247), .Y(n_234) );
INVx2_ASAP7_75t_L g280 ( .A(n_235), .Y(n_280) );
INVx1_ASAP7_75t_L g288 ( .A(n_235), .Y(n_288) );
AND2x2_ASAP7_75t_L g306 ( .A(n_235), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_235), .B(n_290), .Y(n_344) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .Y(n_239) );
AND2x2_ASAP7_75t_L g323 ( .A(n_247), .B(n_280), .Y(n_323) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g276 ( .A(n_248), .Y(n_276) );
AND2x2_ASAP7_75t_L g359 ( .A(n_248), .B(n_290), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_254), .B(n_256), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_254), .A2(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g521 ( .A(n_254), .Y(n_521) );
OAI21xp5_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_266), .B(n_270), .Y(n_259) );
INVx1_ASAP7_75t_SL g304 ( .A(n_260), .Y(n_304) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_261), .B(n_268), .Y(n_361) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g310 ( .A(n_262), .B(n_265), .Y(n_310) );
AND2x2_ASAP7_75t_L g339 ( .A(n_262), .B(n_283), .Y(n_339) );
OR2x2_ASAP7_75t_L g342 ( .A(n_262), .B(n_302), .Y(n_342) );
AOI222xp33_ASAP7_75t_L g406 ( .A1(n_263), .A2(n_355), .B1(n_407), .B2(n_408), .C1(n_410), .C2(n_412), .Y(n_406) );
BUFx2_ASAP7_75t_L g320 ( .A(n_265), .Y(n_320) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g309 ( .A(n_268), .B(n_310), .Y(n_309) );
INVx3_ASAP7_75t_SL g326 ( .A(n_268), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_268), .B(n_320), .Y(n_380) );
AND2x2_ASAP7_75t_L g315 ( .A(n_270), .B(n_275), .Y(n_315) );
INVx1_ASAP7_75t_L g334 ( .A(n_270), .Y(n_334) );
OAI221xp5_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_273), .B1(n_277), .B2(n_281), .C(n_285), .Y(n_271) );
OR2x2_ASAP7_75t_L g343 ( .A(n_273), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g328 ( .A(n_275), .B(n_298), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_275), .B(n_288), .Y(n_368) );
AND2x2_ASAP7_75t_L g373 ( .A(n_275), .B(n_323), .Y(n_373) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_275), .Y(n_383) );
NAND2x1_ASAP7_75t_SL g394 ( .A(n_275), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g279 ( .A(n_276), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_276), .B(n_294), .Y(n_325) );
INVx1_ASAP7_75t_L g391 ( .A(n_276), .Y(n_391) );
INVx1_ASAP7_75t_L g366 ( .A(n_277), .Y(n_366) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g378 ( .A(n_278), .Y(n_378) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_278), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g395 ( .A(n_279), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_279), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g298 ( .A(n_280), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_280), .B(n_290), .Y(n_311) );
INVx1_ASAP7_75t_L g377 ( .A(n_280), .Y(n_377) );
INVx1_ASAP7_75t_L g398 ( .A(n_281), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI21xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_291), .B(n_300), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
AND2x2_ASAP7_75t_L g431 ( .A(n_287), .B(n_364), .Y(n_431) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g399 ( .A(n_288), .B(n_359), .Y(n_399) );
AOI32xp33_ASAP7_75t_L g312 ( .A1(n_289), .A2(n_295), .A3(n_313), .B1(n_315), .B2(n_316), .Y(n_312) );
AOI322xp5_ASAP7_75t_L g414 ( .A1(n_289), .A2(n_321), .A3(n_404), .B1(n_415), .B2(n_416), .C1(n_417), .C2(n_419), .Y(n_414) );
INVx2_ASAP7_75t_L g294 ( .A(n_290), .Y(n_294) );
INVx1_ASAP7_75t_L g404 ( .A(n_290), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B1(n_296), .B2(n_297), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_292), .B(n_298), .Y(n_347) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_293), .B(n_359), .Y(n_409) );
INVx1_ASAP7_75t_L g296 ( .A(n_294), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_294), .B(n_323), .Y(n_413) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_302), .B(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_305), .B1(n_308), .B2(n_311), .C(n_312), .Y(n_303) );
OR2x2_ASAP7_75t_L g324 ( .A(n_305), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g333 ( .A(n_305), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g358 ( .A(n_306), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g362 ( .A(n_316), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B1(n_324), .B2(n_326), .C(n_327), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_320), .A2(n_351), .B1(n_355), .B2(n_356), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_321), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_321), .Y(n_426) );
INVx1_ASAP7_75t_L g420 ( .A(n_323), .Y(n_420) );
INVx1_ASAP7_75t_SL g355 ( .A(n_324), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_326), .B(n_354), .Y(n_416) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_331), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g397 ( .A(n_331), .Y(n_397) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OAI221xp5_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_340), .B1(n_342), .B2(n_343), .C(n_345), .Y(n_335) );
NOR2xp33_ASAP7_75t_SL g336 ( .A(n_337), .B(n_339), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_337), .A2(n_355), .B1(n_401), .B2(n_402), .Y(n_400) );
CKINVDCx14_ASAP7_75t_R g340 ( .A(n_341), .Y(n_340) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_342), .A2(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR3xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_381), .C(n_405), .Y(n_348) );
NAND4xp25_ASAP7_75t_L g349 ( .A(n_350), .B(n_357), .C(n_365), .D(n_372), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g428 ( .A(n_353), .Y(n_428) );
INVx3_ASAP7_75t_SL g422 ( .A(n_354), .Y(n_422) );
OR2x2_ASAP7_75t_L g427 ( .A(n_354), .B(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_362), .B2(n_364), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_359), .B(n_377), .Y(n_418) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI21xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_369), .Y(n_365) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI211xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_384), .B(n_387), .C(n_400), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_392), .B1(n_393), .B2(n_396), .C1(n_398), .C2(n_399), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND4xp25_ASAP7_75t_SL g424 ( .A(n_397), .B(n_425), .C(n_426), .D(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND3xp33_ASAP7_75t_SL g405 ( .A(n_406), .B(n_414), .C(n_423), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_423) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g439 ( .A(n_434), .Y(n_439) );
NOR2x2_ASAP7_75t_L g736 ( .A(n_435), .B(n_726), .Y(n_736) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g725 ( .A(n_436), .B(n_726), .Y(n_725) );
NOR2xp33_ASAP7_75t_SL g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g730 ( .A(n_446), .Y(n_730) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g732 ( .A(n_448), .Y(n_732) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_644), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_593), .C(n_635), .Y(n_449) );
AOI211xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_502), .B(n_547), .C(n_569), .Y(n_450) );
OAI211xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_465), .B(n_486), .C(n_497), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_453), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g656 ( .A(n_453), .B(n_573), .Y(n_656) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g558 ( .A(n_454), .B(n_489), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_454), .B(n_476), .Y(n_675) );
INVx1_ASAP7_75t_L g693 ( .A(n_454), .Y(n_693) );
AND2x2_ASAP7_75t_L g702 ( .A(n_454), .B(n_590), .Y(n_702) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g585 ( .A(n_455), .B(n_476), .Y(n_585) );
AND2x2_ASAP7_75t_L g643 ( .A(n_455), .B(n_590), .Y(n_643) );
INVx1_ASAP7_75t_L g687 ( .A(n_455), .Y(n_687) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g564 ( .A(n_456), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g572 ( .A(n_456), .Y(n_572) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_456), .Y(n_612) );
INVxp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_474), .Y(n_466) );
AND2x2_ASAP7_75t_L g551 ( .A(n_467), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g584 ( .A(n_467), .Y(n_584) );
OR2x2_ASAP7_75t_L g710 ( .A(n_467), .B(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_467), .B(n_476), .Y(n_714) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g489 ( .A(n_468), .Y(n_489) );
INVx1_ASAP7_75t_L g500 ( .A(n_468), .Y(n_500) );
AND2x2_ASAP7_75t_L g573 ( .A(n_468), .B(n_491), .Y(n_573) );
AND2x2_ASAP7_75t_L g613 ( .A(n_468), .B(n_492), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_473), .A2(n_540), .B(n_543), .Y(n_539) );
INVxp67_ASAP7_75t_L g655 ( .A(n_474), .Y(n_655) );
AND2x4_ASAP7_75t_L g680 ( .A(n_474), .B(n_573), .Y(n_680) );
BUFx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_SL g571 ( .A(n_475), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g490 ( .A(n_476), .B(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g559 ( .A(n_476), .B(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g565 ( .A(n_476), .Y(n_565) );
INVx2_ASAP7_75t_L g591 ( .A(n_476), .Y(n_591) );
AND2x2_ASAP7_75t_L g607 ( .A(n_476), .B(n_608), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_487), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
AND2x2_ASAP7_75t_L g670 ( .A(n_489), .B(n_491), .Y(n_670) );
AND2x2_ASAP7_75t_L g587 ( .A(n_490), .B(n_572), .Y(n_587) );
AND2x2_ASAP7_75t_L g686 ( .A(n_490), .B(n_687), .Y(n_686) );
NOR2xp67_ASAP7_75t_L g608 ( .A(n_491), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g711 ( .A(n_491), .B(n_572), .Y(n_711) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g501 ( .A(n_492), .Y(n_501) );
AND2x2_ASAP7_75t_L g590 ( .A(n_492), .B(n_591), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_495), .A2(n_523), .B(n_525), .C(n_526), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_495), .A2(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
AND2x2_ASAP7_75t_L g636 ( .A(n_499), .B(n_571), .Y(n_636) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_500), .B(n_572), .Y(n_621) );
INVx2_ASAP7_75t_L g620 ( .A(n_501), .Y(n_620) );
OAI222xp33_ASAP7_75t_L g624 ( .A1(n_501), .A2(n_564), .B1(n_625), .B2(n_627), .C1(n_628), .C2(n_631), .Y(n_624) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g549 ( .A(n_506), .Y(n_549) );
OR2x2_ASAP7_75t_L g660 ( .A(n_506), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g582 ( .A(n_507), .Y(n_582) );
NOR2x1_ASAP7_75t_L g633 ( .A(n_507), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g639 ( .A(n_507), .B(n_553), .Y(n_639) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g600 ( .A(n_508), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_513), .A2(n_603), .B1(n_642), .B2(n_643), .Y(n_641) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_528), .Y(n_513) );
INVx3_ASAP7_75t_L g575 ( .A(n_514), .Y(n_575) );
OR2x2_ASAP7_75t_L g708 ( .A(n_514), .B(n_584), .Y(n_708) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g581 ( .A(n_515), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g597 ( .A(n_515), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g605 ( .A(n_515), .B(n_553), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_515), .B(n_529), .Y(n_661) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g552 ( .A(n_516), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g556 ( .A(n_516), .B(n_529), .Y(n_556) );
AND2x2_ASAP7_75t_L g632 ( .A(n_516), .B(n_579), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_516), .B(n_538), .Y(n_672) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_528), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g588 ( .A(n_528), .B(n_549), .Y(n_588) );
AND2x2_ASAP7_75t_L g592 ( .A(n_528), .B(n_582), .Y(n_592) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
INVx3_ASAP7_75t_L g553 ( .A(n_529), .Y(n_553) );
AND2x2_ASAP7_75t_L g578 ( .A(n_529), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g713 ( .A(n_529), .B(n_696), .Y(n_713) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_538), .Y(n_567) );
INVx2_ASAP7_75t_L g579 ( .A(n_538), .Y(n_579) );
AND2x2_ASAP7_75t_L g623 ( .A(n_538), .B(n_599), .Y(n_623) );
INVx1_ASAP7_75t_L g666 ( .A(n_538), .Y(n_666) );
OR2x2_ASAP7_75t_L g697 ( .A(n_538), .B(n_599), .Y(n_697) );
AND2x2_ASAP7_75t_L g717 ( .A(n_538), .B(n_553), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_550), .B(n_554), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g555 ( .A(n_549), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_549), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g674 ( .A(n_551), .Y(n_674) );
INVx2_ASAP7_75t_SL g568 ( .A(n_552), .Y(n_568) );
AND2x2_ASAP7_75t_L g688 ( .A(n_552), .B(n_582), .Y(n_688) );
INVx2_ASAP7_75t_L g634 ( .A(n_553), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_553), .B(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_557), .B1(n_560), .B2(n_566), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_556), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g722 ( .A(n_556), .Y(n_722) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g647 ( .A(n_558), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_558), .B(n_590), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_559), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g663 ( .A(n_559), .B(n_612), .Y(n_663) );
INVx2_ASAP7_75t_L g719 ( .A(n_559), .Y(n_719) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g589 ( .A(n_562), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_562), .B(n_607), .Y(n_640) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_564), .B(n_584), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g701 ( .A(n_567), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_SL g651 ( .A1(n_568), .A2(n_652), .B(n_654), .C(n_657), .Y(n_651) );
OR2x2_ASAP7_75t_L g678 ( .A(n_568), .B(n_582), .Y(n_678) );
OAI221xp5_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_574), .B1(n_576), .B2(n_583), .C(n_586), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_571), .B(n_573), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_571), .B(n_620), .Y(n_627) );
AND2x2_ASAP7_75t_L g669 ( .A(n_571), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g705 ( .A(n_571), .Y(n_705) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_572), .Y(n_596) );
INVx1_ASAP7_75t_L g609 ( .A(n_572), .Y(n_609) );
NOR2xp67_ASAP7_75t_L g629 ( .A(n_575), .B(n_630), .Y(n_629) );
INVxp67_ASAP7_75t_L g683 ( .A(n_575), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_575), .B(n_623), .Y(n_699) );
INVx2_ASAP7_75t_L g685 ( .A(n_576), .Y(n_685) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g626 ( .A(n_578), .B(n_597), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_578), .A2(n_594), .B(n_636), .C(n_637), .Y(n_635) );
AND2x2_ASAP7_75t_L g604 ( .A(n_579), .B(n_599), .Y(n_604) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_583), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
OR2x2_ASAP7_75t_L g652 ( .A(n_584), .B(n_653), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_589), .B2(n_592), .Y(n_586) );
INVx1_ASAP7_75t_L g706 ( .A(n_588), .Y(n_706) );
INVx1_ASAP7_75t_L g653 ( .A(n_590), .Y(n_653) );
INVx1_ASAP7_75t_L g704 ( .A(n_592), .Y(n_704) );
AOI211xp5_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_597), .B(n_601), .C(n_624), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g616 ( .A(n_596), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g667 ( .A(n_597), .Y(n_667) );
AND2x2_ASAP7_75t_L g716 ( .A(n_597), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_606), .B(n_614), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx2_ASAP7_75t_L g630 ( .A(n_604), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_604), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g622 ( .A(n_605), .B(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g698 ( .A(n_605), .Y(n_698) );
OAI32xp33_ASAP7_75t_L g709 ( .A1(n_605), .A2(n_657), .A3(n_664), .B1(n_705), .B2(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_SL g606 ( .A(n_607), .B(n_610), .Y(n_606) );
INVx1_ASAP7_75t_SL g677 ( .A(n_607), .Y(n_677) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g617 ( .A(n_613), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .B(n_622), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_616), .A2(n_664), .B1(n_690), .B2(n_692), .Y(n_689) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_620), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g657 ( .A(n_623), .Y(n_657) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2x1p5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g650 ( .A(n_634), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_641), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_643), .A2(n_685), .B1(n_686), .B2(n_688), .C(n_689), .Y(n_684) );
NAND5xp2_ASAP7_75t_L g644 ( .A(n_645), .B(n_668), .C(n_684), .D(n_694), .E(n_712), .Y(n_644) );
AOI211xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_648), .B(n_651), .C(n_658), .Y(n_645) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g715 ( .A(n_652), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_662), .B2(n_664), .Y(n_658) );
INVx1_ASAP7_75t_SL g691 ( .A(n_661), .Y(n_691) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI322xp33_ASAP7_75t_L g673 ( .A1(n_664), .A2(n_674), .A3(n_675), .B1(n_676), .B2(n_677), .C1(n_678), .C2(n_679), .Y(n_673) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g676 ( .A(n_666), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_666), .B(n_691), .Y(n_690) );
AOI211xp5_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_671), .B(n_673), .C(n_681), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_677), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_703) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g720 ( .A(n_687), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_702), .B1(n_703), .B2(n_707), .C(n_709), .Y(n_694) );
OAI211xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_698), .B(n_699), .C(n_700), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g721 ( .A(n_697), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B1(n_715), .B2(n_716), .C(n_718), .Y(n_712) );
AOI21xp33_ASAP7_75t_SL g718 ( .A1(n_719), .A2(n_720), .B(n_721), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_723), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
endmodule