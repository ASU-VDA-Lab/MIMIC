module fake_jpeg_19036_n_298 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_9),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_21),
.B(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_42),
.B(n_25),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_20),
.B(n_16),
.C(n_27),
.Y(n_45)
);

XNOR2x1_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_53),
.Y(n_61)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_31),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_31),
.B1(n_40),
.B2(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_31),
.B1(n_25),
.B2(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_39),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_64),
.C(n_41),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_41),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_47),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_101),
.B(n_102),
.Y(n_116)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_61),
.B1(n_65),
.B2(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_96),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_66),
.A2(n_31),
.B1(n_44),
.B2(n_58),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_44),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_70),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_43),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_33),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_71),
.Y(n_122)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_125),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_85),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_62),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_106),
.B(n_87),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_101),
.B(n_102),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_91),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_62),
.C(n_82),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_138),
.C(n_32),
.Y(n_164)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_28),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_97),
.C(n_87),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_102),
.B1(n_101),
.B2(n_95),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_145),
.B1(n_152),
.B2(n_154),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_146),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_124),
.B1(n_118),
.B2(n_125),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_99),
.Y(n_146)
);

AO22x1_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_76),
.B1(n_79),
.B2(n_99),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_148),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_127),
.B1(n_116),
.B2(n_113),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_78),
.B1(n_81),
.B2(n_90),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_161),
.B1(n_167),
.B2(n_131),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_110),
.B1(n_66),
.B2(n_67),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_19),
.B(n_94),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_157),
.B(n_19),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_88),
.B(n_8),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_88),
.B(n_105),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_134),
.B(n_112),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_84),
.B1(n_67),
.B2(n_72),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_163),
.B1(n_32),
.B2(n_22),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_56),
.C(n_19),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_23),
.B(n_17),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_111),
.B1(n_90),
.B2(n_92),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_92),
.B1(n_94),
.B2(n_33),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_165),
.C(n_28),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_24),
.C(n_28),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_26),
.B1(n_17),
.B2(n_27),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_132),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_175),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_174),
.Y(n_204)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_134),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_177),
.A2(n_178),
.B(n_190),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_112),
.B(n_2),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_184),
.B1(n_165),
.B2(n_166),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_30),
.B1(n_16),
.B2(n_27),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_191),
.B1(n_193),
.B2(n_139),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_162),
.B(n_16),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_181),
.B(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_23),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_17),
.B(n_23),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_185),
.A2(n_0),
.B(n_2),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_32),
.A3(n_22),
.B1(n_28),
.B2(n_24),
.C1(n_30),
.C2(n_7),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_147),
.C(n_163),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_22),
.C(n_2),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_142),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_30),
.B(n_32),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_0),
.B(n_2),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_144),
.B(n_154),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_161),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_195),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_172),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_146),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_208),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_164),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_215),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_213),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_195),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_207),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_140),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_170),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_166),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_217),
.A2(n_185),
.B1(n_179),
.B2(n_178),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_187),
.C(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_216),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_170),
.B1(n_188),
.B2(n_175),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_232),
.B1(n_235),
.B2(n_196),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_204),
.B1(n_201),
.B2(n_217),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_172),
.C(n_177),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_216),
.C(n_215),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_233),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_206),
.A2(n_183),
.B1(n_186),
.B2(n_190),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_229),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_173),
.B1(n_183),
.B2(n_180),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_191),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_209),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_251),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_208),
.C(n_198),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_244),
.C(n_231),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_197),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_248),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_197),
.C(n_205),
.Y(n_244)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_205),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_248),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_250),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_181),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_226),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_259),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_258),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_228),
.B(n_225),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_8),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_235),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_219),
.C(n_224),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_230),
.C(n_182),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_234),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_9),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_223),
.B1(n_241),
.B2(n_243),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_249),
.B(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_268),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_212),
.B(n_194),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_22),
.B1(n_9),
.B2(n_10),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_272),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_15),
.B(n_11),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_262),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_254),
.B(n_263),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_267),
.A2(n_258),
.B1(n_263),
.B2(n_254),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_283),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_11),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_0),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_282),
.B(n_12),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_271),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_277),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_265),
.B1(n_273),
.B2(n_11),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_12),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_285),
.Y(n_293)
);

AOI321xp33_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_276),
.A3(n_292),
.B1(n_284),
.B2(n_290),
.C(n_5),
.Y(n_294)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_285),
.C(n_271),
.Y(n_295)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_295),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_296),
.A2(n_3),
.B(n_4),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_3),
.Y(n_298)
);


endmodule