module fake_jpeg_10727_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_64),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_0),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_57),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_61),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_76),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_59),
.B(n_50),
.C(n_45),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_68),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_47),
.B1(n_52),
.B2(n_61),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_79),
.B1(n_60),
.B2(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_56),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_82),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_47),
.B1(n_52),
.B2(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_46),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_94),
.Y(n_102)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_96),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_54),
.C(n_20),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_16),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_18),
.B1(n_42),
.B2(n_40),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_17),
.B1(n_38),
.B2(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_72),
.B(n_3),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_108),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_90),
.B1(n_93),
.B2(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_105),
.B(n_101),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_121),
.Y(n_131)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_14),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_15),
.B1(n_23),
.B2(n_24),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_101),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_43),
.C(n_27),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_115),
.C(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_136),
.Y(n_139)
);

OAI321xp33_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_120),
.A3(n_122),
.B1(n_121),
.B2(n_130),
.C(n_118),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_110),
.B(n_29),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_138),
.B(n_140),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_134),
.B(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_134),
.Y(n_144)
);

OAI31xp33_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_142),
.A3(n_139),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_127),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_146),
.A2(n_25),
.B(n_30),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_31),
.C(n_36),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);


endmodule