module fake_jpeg_14041_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_9),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_6),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_24),
.Y(n_30)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_18),
.B1(n_16),
.B2(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_20),
.B1(n_28),
.B2(n_23),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_45),
.Y(n_51)
);

AND2x6_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_7),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_25),
.B1(n_28),
.B2(n_15),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_48),
.B1(n_33),
.B2(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_8),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_30),
.A2(n_25),
.B1(n_15),
.B2(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_40),
.B(n_36),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_19),
.C(n_26),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_62),
.C(n_63),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_26),
.C(n_14),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_36),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_14),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_53),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_27),
.C(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_66),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_27),
.C(n_32),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_53),
.B1(n_55),
.B2(n_58),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_31),
.B(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_51),
.B1(n_58),
.B2(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_63),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_52),
.C(n_27),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_78),
.B(n_79),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_31),
.C(n_46),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_73),
.B1(n_70),
.B2(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_82),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_73),
.B1(n_23),
.B2(n_4),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_35),
.B(n_22),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_86),
.C(n_31),
.Y(n_87)
);

AOI21x1_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_31),
.B(n_35),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_35),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_6),
.Y(n_88)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_5),
.B(n_7),
.Y(n_89)
);

AOI21x1_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_90),
.B(n_2),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_4),
.B(n_2),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_3),
.Y(n_93)
);


endmodule