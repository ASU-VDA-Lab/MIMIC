module real_aes_880_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_813, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_812, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_814, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_813;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_812;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_814;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_656;
wire n_532;
wire n_316;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_331;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_397;
wire n_358;
wire n_293;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_762;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_639;
wire n_546;
wire n_587;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_554;
wire n_475;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_0), .A2(n_238), .B1(n_478), .B2(n_609), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_1), .A2(n_115), .B1(n_386), .B2(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_2), .A2(n_251), .B1(n_386), .B2(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_3), .A2(n_132), .B1(n_433), .B2(n_447), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_4), .A2(n_161), .B1(n_525), .B2(n_526), .Y(n_524) );
AOI222xp33_ASAP7_75t_L g495 ( .A1(n_5), .A2(n_99), .B1(n_284), .B2(n_298), .C1(n_314), .C2(n_328), .Y(n_495) );
OA22x2_ASAP7_75t_L g559 ( .A1(n_6), .A2(n_560), .B1(n_561), .B2(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_6), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_7), .A2(n_92), .B1(n_418), .B2(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_8), .A2(n_147), .B1(n_617), .B2(n_650), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_9), .A2(n_182), .B1(n_351), .B2(n_352), .Y(n_490) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_10), .A2(n_210), .B1(n_301), .B2(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g751 ( .A(n_10), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_11), .A2(n_187), .B1(n_348), .B2(n_349), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_12), .A2(n_213), .B1(n_554), .B2(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_13), .A2(n_37), .B1(n_416), .B2(n_423), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_14), .B(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_15), .A2(n_85), .B1(n_523), .B2(n_611), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_16), .A2(n_137), .B1(n_343), .B2(n_345), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_17), .A2(n_209), .B1(n_332), .B2(n_333), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_18), .A2(n_120), .B1(n_390), .B2(n_393), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_19), .A2(n_199), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_20), .A2(n_135), .B1(n_416), .B2(n_514), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g607 ( .A1(n_21), .A2(n_62), .B1(n_245), .B2(n_380), .C1(n_608), .C2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_22), .A2(n_42), .B1(n_318), .B2(n_323), .Y(n_317) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_23), .A2(n_234), .B1(n_638), .B2(n_639), .Y(n_696) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_24), .A2(n_80), .B1(n_301), .B2(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_24), .B(n_750), .Y(n_749) );
OA22x2_ASAP7_75t_L g725 ( .A1(n_25), .A2(n_726), .B1(n_737), .B2(n_738), .Y(n_725) );
INVx1_ASAP7_75t_L g737 ( .A(n_25), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_26), .A2(n_76), .B1(n_433), .B2(n_434), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_27), .A2(n_218), .B1(n_595), .B2(n_596), .Y(n_594) );
AOI22xp5_ASAP7_75t_SL g427 ( .A1(n_28), .A2(n_257), .B1(n_361), .B2(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g604 ( .A(n_29), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_30), .A2(n_285), .B1(n_370), .B2(n_654), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_31), .A2(n_217), .B1(n_653), .B2(n_654), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_32), .A2(n_171), .B1(n_418), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_33), .A2(n_44), .B1(n_340), .B2(n_492), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_34), .A2(n_206), .B1(n_421), .B2(n_551), .Y(n_550) );
OA22x2_ASAP7_75t_L g582 ( .A1(n_35), .A2(n_583), .B1(n_584), .B2(n_600), .Y(n_582) );
INVx1_ASAP7_75t_L g600 ( .A(n_35), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_36), .A2(n_202), .B1(n_399), .B2(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_38), .A2(n_278), .B1(n_549), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_39), .A2(n_194), .B1(n_699), .B2(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_40), .A2(n_134), .B1(n_377), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_41), .A2(n_248), .B1(n_298), .B2(n_314), .Y(n_297) );
OA22x2_ASAP7_75t_L g687 ( .A1(n_43), .A2(n_688), .B1(n_689), .B2(n_705), .Y(n_687) );
INVx1_ASAP7_75t_L g705 ( .A(n_43), .Y(n_705) );
INVx1_ASAP7_75t_L g452 ( .A(n_45), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_45), .A2(n_46), .B(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_45), .A2(n_471), .B1(n_480), .B2(n_814), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_46), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_47), .A2(n_247), .B1(n_332), .B2(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_48), .B(n_426), .Y(n_425) );
AOI222xp33_ASAP7_75t_SL g475 ( .A1(n_49), .A2(n_131), .B1(n_183), .B2(n_476), .C1(n_477), .C2(n_478), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_50), .A2(n_95), .B1(n_416), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_51), .A2(n_203), .B1(n_375), .B2(n_455), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_52), .A2(n_226), .B1(n_433), .B2(n_447), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_53), .A2(n_58), .B1(n_384), .B2(n_386), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_54), .A2(n_190), .B1(n_641), .B2(n_642), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_55), .Y(n_805) );
AOI22xp33_ASAP7_75t_SL g612 ( .A1(n_56), .A2(n_114), .B1(n_386), .B2(n_613), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_57), .A2(n_280), .B1(n_351), .B2(n_352), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_59), .A2(n_258), .B1(n_373), .B2(n_473), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_60), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_61), .A2(n_228), .B1(n_596), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_63), .A2(n_219), .B1(n_590), .B2(n_649), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_64), .A2(n_283), .B1(n_397), .B2(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_65), .A2(n_223), .B1(n_641), .B2(n_642), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_66), .A2(n_195), .B1(n_458), .B2(n_459), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_67), .A2(n_77), .B1(n_543), .B2(n_598), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_68), .A2(n_129), .B1(n_386), .B2(n_543), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_69), .A2(n_276), .B1(n_433), .B2(n_523), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_70), .A2(n_86), .B1(n_638), .B2(n_639), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_71), .A2(n_108), .B1(n_458), .B2(n_459), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_72), .A2(n_764), .B1(n_784), .B2(n_785), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_72), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_73), .A2(n_118), .B1(n_348), .B2(n_349), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_74), .A2(n_139), .B1(n_433), .B2(n_447), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_75), .A2(n_235), .B1(n_617), .B2(n_650), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_78), .A2(n_166), .B1(n_676), .B2(n_678), .Y(n_675) );
AOI222xp33_ASAP7_75t_L g720 ( .A1(n_79), .A2(n_81), .B1(n_277), .B2(n_566), .C1(n_721), .C2(n_722), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_82), .A2(n_121), .B1(n_358), .B2(n_609), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_83), .A2(n_250), .B1(n_649), .B2(n_651), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_84), .A2(n_103), .B1(n_412), .B2(n_413), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_87), .A2(n_205), .B1(n_343), .B2(n_345), .Y(n_493) );
INVx3_ASAP7_75t_L g301 ( .A(n_88), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_89), .A2(n_174), .B1(n_318), .B2(n_323), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_90), .A2(n_155), .B1(n_375), .B2(n_377), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_91), .A2(n_207), .B1(n_390), .B2(n_514), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_93), .A2(n_282), .B1(n_390), .B2(n_460), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_94), .A2(n_262), .B1(n_393), .B2(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_96), .A2(n_173), .B1(n_348), .B2(n_349), .Y(n_347) );
OA22x2_ASAP7_75t_L g708 ( .A1(n_97), .A2(n_709), .B1(n_710), .B2(n_723), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_97), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_98), .B(n_426), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_100), .A2(n_225), .B1(n_449), .B2(n_450), .Y(n_448) );
AO22x2_ASAP7_75t_L g627 ( .A1(n_101), .A2(n_628), .B1(n_629), .B2(n_656), .Y(n_627) );
INVx1_ASAP7_75t_L g656 ( .A(n_101), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_102), .A2(n_214), .B1(n_554), .B2(n_700), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_104), .A2(n_172), .B1(n_421), .B2(n_423), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_105), .A2(n_149), .B1(n_298), .B2(n_526), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_106), .A2(n_136), .B1(n_412), .B2(n_413), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_107), .A2(n_201), .B1(n_412), .B2(n_413), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_109), .A2(n_168), .B1(n_641), .B2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_110), .A2(n_150), .B1(n_458), .B2(n_459), .Y(n_655) );
INVx1_ASAP7_75t_SL g306 ( .A(n_111), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_111), .B(n_146), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_112), .A2(n_232), .B1(n_397), .B2(n_399), .Y(n_396) );
AOI222xp33_ASAP7_75t_L g691 ( .A1(n_113), .A2(n_141), .B1(n_267), .B2(n_635), .C1(n_642), .C2(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g759 ( .A(n_116), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_117), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_119), .A2(n_184), .B1(n_349), .B2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_122), .A2(n_270), .B1(n_339), .B2(n_340), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_123), .A2(n_256), .B1(n_478), .B2(n_635), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_124), .B(n_426), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_125), .A2(n_230), .B1(n_332), .B2(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_126), .A2(n_246), .B1(n_375), .B2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_127), .A2(n_140), .B1(n_596), .B2(n_609), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_128), .A2(n_279), .B1(n_364), .B2(n_366), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_130), .A2(n_181), .B1(n_575), .B2(n_647), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_133), .Y(n_498) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_138), .A2(n_211), .B1(n_318), .B2(n_323), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_142), .A2(n_255), .B1(n_399), .B2(n_421), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_143), .B(n_692), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_144), .A2(n_175), .B1(n_375), .B2(n_460), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_145), .A2(n_185), .B1(n_373), .B2(n_505), .Y(n_734) );
AO22x2_ASAP7_75t_L g300 ( .A1(n_146), .A2(n_220), .B1(n_301), .B2(n_302), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_148), .A2(n_236), .B1(n_384), .B2(n_386), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_151), .B(n_426), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_152), .A2(n_215), .B1(n_680), .B2(n_681), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_153), .A2(n_193), .B1(n_370), .B2(n_373), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_154), .A2(n_204), .B1(n_384), .B2(n_386), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_156), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_157), .A2(n_178), .B1(n_416), .B2(n_460), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_158), .A2(n_196), .B1(n_460), .B2(n_512), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_159), .A2(n_244), .B1(n_433), .B2(n_447), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_160), .A2(n_274), .B1(n_412), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_162), .A2(n_170), .B1(n_400), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_163), .A2(n_269), .B1(n_588), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_164), .A2(n_263), .B1(n_801), .B2(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g307 ( .A(n_165), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_167), .A2(n_197), .B1(n_358), .B2(n_361), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_169), .B(n_569), .Y(n_731) );
AO21x1_ASAP7_75t_SL g753 ( .A1(n_176), .A2(n_754), .B(n_762), .Y(n_753) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_177), .A2(n_242), .B1(n_358), .B2(n_361), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_179), .B(n_328), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_180), .A2(n_281), .B1(n_588), .B2(n_702), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_186), .A2(n_188), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_189), .A2(n_260), .B1(n_339), .B2(n_340), .Y(n_338) );
XNOR2x1_ASAP7_75t_L g354 ( .A(n_191), .B(n_355), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_192), .A2(n_222), .B1(n_416), .B2(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_198), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g660 ( .A(n_200), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_208), .A2(n_221), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_212), .A2(n_231), .B1(n_298), .B2(n_526), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_216), .A2(n_261), .B1(n_370), .B2(n_373), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_224), .A2(n_275), .B1(n_649), .B2(n_651), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_227), .Y(n_436) );
INVx1_ASAP7_75t_L g746 ( .A(n_229), .Y(n_746) );
AND2x4_ASAP7_75t_L g761 ( .A(n_229), .B(n_747), .Y(n_761) );
AO21x1_ASAP7_75t_L g809 ( .A1(n_229), .A2(n_757), .B(n_810), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_233), .A2(n_271), .B1(n_443), .B2(n_446), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_237), .A2(n_266), .B1(n_351), .B2(n_352), .Y(n_576) );
INVx1_ASAP7_75t_L g747 ( .A(n_239), .Y(n_747) );
AND2x2_ASAP7_75t_R g787 ( .A(n_239), .B(n_746), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_240), .A2(n_243), .B1(n_458), .B2(n_459), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_241), .B(n_380), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_249), .A2(n_259), .B1(n_364), .B2(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_252), .A2(n_265), .B1(n_384), .B2(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g758 ( .A(n_253), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_254), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_264), .A2(n_268), .B1(n_433), .B2(n_447), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_272), .B(n_632), .Y(n_631) );
AO22x1_ASAP7_75t_L g539 ( .A1(n_273), .A2(n_540), .B1(n_557), .B2(n_558), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_273), .Y(n_557) );
AOI21xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_742), .B(n_753), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_623), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI21xp33_ASAP7_75t_L g742 ( .A1(n_289), .A2(n_624), .B(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_534), .B1(n_535), .B2(n_622), .Y(n_289) );
INVx1_ASAP7_75t_L g622 ( .A(n_290), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_403), .B(n_531), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_291), .A2(n_405), .B(n_532), .C(n_533), .Y(n_531) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_354), .B1(n_401), .B2(n_402), .Y(n_291) );
OA22x2_ASAP7_75t_L g407 ( .A1(n_292), .A2(n_293), .B1(n_408), .B2(n_437), .Y(n_407) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
XOR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_353), .Y(n_293) );
XOR2x2_ASAP7_75t_L g402 ( .A(n_294), .B(n_353), .Y(n_402) );
NAND2x1_ASAP7_75t_SL g294 ( .A(n_295), .B(n_336), .Y(n_294) );
NOR2x1_ASAP7_75t_L g295 ( .A(n_296), .B(n_326), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_317), .Y(n_296) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_308), .Y(n_298) );
AND2x2_ASAP7_75t_L g339 ( .A(n_299), .B(n_319), .Y(n_339) );
AND2x6_ASAP7_75t_L g348 ( .A(n_299), .B(n_329), .Y(n_348) );
AND2x4_ASAP7_75t_L g362 ( .A(n_299), .B(n_308), .Y(n_362) );
AND2x2_ASAP7_75t_L g372 ( .A(n_299), .B(n_319), .Y(n_372) );
AND2x2_ASAP7_75t_L g398 ( .A(n_299), .B(n_329), .Y(n_398) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_299), .B(n_319), .Y(n_492) );
AND2x2_ASAP7_75t_L g525 ( .A(n_299), .B(n_308), .Y(n_525) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
AND2x2_ASAP7_75t_L g316 ( .A(n_300), .B(n_304), .Y(n_316) );
INVx2_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
BUFx2_ASAP7_75t_L g341 ( .A(n_300), .Y(n_341) );
INVx1_ASAP7_75t_L g302 ( .A(n_301), .Y(n_302) );
OAI22x1_ASAP7_75t_L g304 ( .A1(n_301), .A2(n_305), .B1(n_306), .B2(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_301), .Y(n_305) );
INVx2_ASAP7_75t_L g310 ( .A(n_301), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_301), .Y(n_313) );
AND2x4_ASAP7_75t_L g344 ( .A(n_303), .B(n_322), .Y(n_344) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g321 ( .A(n_304), .B(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
AND2x4_ASAP7_75t_L g332 ( .A(n_308), .B(n_321), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_344), .Y(n_345) );
AND2x2_ASAP7_75t_L g385 ( .A(n_308), .B(n_321), .Y(n_385) );
AND2x4_ASAP7_75t_L g400 ( .A(n_308), .B(n_344), .Y(n_400) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g320 ( .A(n_309), .Y(n_320) );
INVx1_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
AND2x2_ASAP7_75t_L g335 ( .A(n_309), .B(n_312), .Y(n_335) );
INVxp67_ASAP7_75t_L g315 ( .A(n_311), .Y(n_315) );
AND2x4_ASAP7_75t_L g329 ( .A(n_311), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g319 ( .A(n_312), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x4_ASAP7_75t_L g360 ( .A(n_315), .B(n_316), .Y(n_360) );
AND2x2_ASAP7_75t_L g526 ( .A(n_315), .B(n_316), .Y(n_526) );
AND2x2_ASAP7_75t_L g323 ( .A(n_316), .B(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g328 ( .A(n_316), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g367 ( .A(n_316), .B(n_324), .Y(n_367) );
AND2x2_ASAP7_75t_L g382 ( .A(n_316), .B(n_329), .Y(n_382) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
AND2x6_ASAP7_75t_L g349 ( .A(n_319), .B(n_344), .Y(n_349) );
AND2x2_ASAP7_75t_L g365 ( .A(n_319), .B(n_321), .Y(n_365) );
AND2x4_ASAP7_75t_L g395 ( .A(n_319), .B(n_344), .Y(n_395) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_320), .Y(n_325) );
AND2x2_ASAP7_75t_L g351 ( .A(n_321), .B(n_329), .Y(n_351) );
AND2x4_ASAP7_75t_L g376 ( .A(n_321), .B(n_329), .Y(n_376) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_331), .Y(n_326) );
INVx2_ASAP7_75t_SL g518 ( .A(n_328), .Y(n_518) );
BUFx2_ASAP7_75t_L g721 ( .A(n_328), .Y(n_721) );
AND2x2_ASAP7_75t_L g343 ( .A(n_329), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g392 ( .A(n_329), .B(n_344), .Y(n_392) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_332), .Y(n_722) );
AND2x2_ASAP7_75t_SL g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g387 ( .A(n_334), .B(n_335), .Y(n_387) );
AND2x2_ASAP7_75t_SL g566 ( .A(n_334), .B(n_335), .Y(n_566) );
AND2x4_ASAP7_75t_L g340 ( .A(n_335), .B(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g352 ( .A(n_335), .B(n_344), .Y(n_352) );
AND2x4_ASAP7_75t_L g373 ( .A(n_335), .B(n_341), .Y(n_373) );
AND2x4_ASAP7_75t_L g377 ( .A(n_335), .B(n_344), .Y(n_377) );
NOR2x1_ASAP7_75t_L g336 ( .A(n_337), .B(n_346), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_342), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_350), .Y(n_346) );
INVx1_ASAP7_75t_L g509 ( .A(n_348), .Y(n_509) );
INVx2_ASAP7_75t_L g401 ( .A(n_354), .Y(n_401) );
NAND4xp75_ASAP7_75t_L g355 ( .A(n_356), .B(n_368), .C(n_378), .D(n_388), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_363), .Y(n_356) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g428 ( .A(n_359), .Y(n_428) );
INVx2_ASAP7_75t_L g478 ( .A(n_359), .Y(n_478) );
INVx2_ASAP7_75t_L g596 ( .A(n_359), .Y(n_596) );
INVx2_ASAP7_75t_SL g608 ( .A(n_359), .Y(n_608) );
INVx2_ASAP7_75t_L g695 ( .A(n_359), .Y(n_695) );
INVx6_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_362), .Y(n_477) );
BUFx2_ASAP7_75t_L g595 ( .A(n_362), .Y(n_595) );
BUFx3_ASAP7_75t_L g609 ( .A(n_362), .Y(n_609) );
BUFx6f_ASAP7_75t_SL g641 ( .A(n_364), .Y(n_641) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_365), .Y(n_433) );
INVx3_ASAP7_75t_L g445 ( .A(n_365), .Y(n_445) );
BUFx4f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g435 ( .A(n_367), .Y(n_435) );
BUFx3_ASAP7_75t_L g447 ( .A(n_367), .Y(n_447) );
BUFx6f_ASAP7_75t_SL g523 ( .A(n_367), .Y(n_523) );
INVx2_ASAP7_75t_L g644 ( .A(n_367), .Y(n_644) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g474 ( .A(n_371), .Y(n_474) );
INVx1_ASAP7_75t_L g505 ( .A(n_371), .Y(n_505) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_372), .Y(n_412) );
BUFx3_ASAP7_75t_L g700 ( .A(n_372), .Y(n_700) );
INVx5_ASAP7_75t_SL g414 ( .A(n_373), .Y(n_414) );
BUFx2_ASAP7_75t_L g506 ( .A(n_373), .Y(n_506) );
BUFx3_ASAP7_75t_L g554 ( .A(n_373), .Y(n_554) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx6_ASAP7_75t_L g422 ( .A(n_376), .Y(n_422) );
BUFx3_ASAP7_75t_L g512 ( .A(n_376), .Y(n_512) );
BUFx3_ASAP7_75t_L g423 ( .A(n_377), .Y(n_423) );
BUFx3_ASAP7_75t_L g460 ( .A(n_377), .Y(n_460) );
INVx2_ASAP7_75t_L g552 ( .A(n_377), .Y(n_552) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_383), .Y(n_378) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx4_ASAP7_75t_SL g426 ( .A(n_381), .Y(n_426) );
INVx3_ASAP7_75t_L g476 ( .A(n_381), .Y(n_476) );
INVx3_ASAP7_75t_SL g569 ( .A(n_381), .Y(n_569) );
INVx4_ASAP7_75t_SL g633 ( .A(n_381), .Y(n_633) );
BUFx2_ASAP7_75t_L g776 ( .A(n_381), .Y(n_776) );
INVx6_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_384), .Y(n_638) );
BUFx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g463 ( .A(n_385), .Y(n_463) );
BUFx5_ASAP7_75t_L g613 ( .A(n_385), .Y(n_613) );
BUFx3_ASAP7_75t_L g779 ( .A(n_385), .Y(n_779) );
INVx2_ASAP7_75t_L g803 ( .A(n_386), .Y(n_803) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx3_ASAP7_75t_L g431 ( .A(n_387), .Y(n_431) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_396), .Y(n_388) );
INVx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
INVx2_ASAP7_75t_SL g468 ( .A(n_391), .Y(n_468) );
INVx2_ASAP7_75t_L g647 ( .A(n_391), .Y(n_647) );
INVx4_ASAP7_75t_L g677 ( .A(n_391), .Y(n_677) );
INVx3_ASAP7_75t_SL g702 ( .A(n_391), .Y(n_702) );
INVx8_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g449 ( .A(n_394), .Y(n_449) );
INVx2_ASAP7_75t_L g549 ( .A(n_394), .Y(n_549) );
INVx2_ASAP7_75t_SL g590 ( .A(n_394), .Y(n_590) );
INVx2_ASAP7_75t_L g617 ( .A(n_394), .Y(n_617) );
INVx2_ASAP7_75t_L g651 ( .A(n_394), .Y(n_651) );
INVx1_ASAP7_75t_SL g681 ( .A(n_394), .Y(n_681) );
INVx8_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g451 ( .A(n_397), .Y(n_451) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx3_ASAP7_75t_L g419 ( .A(n_398), .Y(n_419) );
BUFx2_ASAP7_75t_L g650 ( .A(n_398), .Y(n_650) );
INVx1_ASAP7_75t_L g666 ( .A(n_399), .Y(n_666) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx3_ASAP7_75t_L g455 ( .A(n_400), .Y(n_455) );
INVx2_ASAP7_75t_L g515 ( .A(n_400), .Y(n_515) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_400), .Y(n_556) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_400), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_438), .B(n_530), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_407), .B(n_438), .Y(n_530) );
INVx1_ASAP7_75t_SL g437 ( .A(n_408), .Y(n_437) );
XNOR2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_436), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_424), .Y(n_409) );
NAND4xp25_ASAP7_75t_L g410 ( .A(n_411), .B(n_415), .C(n_417), .D(n_420), .Y(n_410) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g654 ( .A(n_414), .Y(n_654) );
INVx2_ASAP7_75t_L g795 ( .A(n_414), .Y(n_795) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_SL g680 ( .A(n_419), .Y(n_680) );
INVx3_ASAP7_75t_L g773 ( .A(n_419), .Y(n_773) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g458 ( .A(n_422), .Y(n_458) );
INVx2_ASAP7_75t_L g664 ( .A(n_422), .Y(n_664) );
NAND4xp25_ASAP7_75t_SL g424 ( .A(n_425), .B(n_427), .C(n_429), .D(n_432), .Y(n_424) );
BUFx2_ASAP7_75t_L g639 ( .A(n_430), .Y(n_639) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g598 ( .A(n_431), .Y(n_598) );
INVx3_ASAP7_75t_L g780 ( .A(n_431), .Y(n_780) );
INVx2_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g532 ( .A(n_438), .Y(n_532) );
OA22x2_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_483), .B1(n_484), .B2(n_529), .Y(n_438) );
INVx2_ASAP7_75t_SL g529 ( .A(n_439), .Y(n_529) );
OR2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_464), .Y(n_439) );
OAI222xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_452), .B1(n_453), .B2(n_456), .C1(n_812), .C2(n_813), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_441), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_448), .Y(n_441) );
BUFx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g611 ( .A(n_445), .Y(n_611) );
BUFx6f_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_453), .B(n_456), .C(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_457), .B(n_461), .Y(n_456) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g543 ( .A(n_463), .Y(n_543) );
INVx2_ASAP7_75t_L g801 ( .A(n_463), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_469), .B(n_479), .Y(n_464) );
INVx1_ASAP7_75t_L g482 ( .A(n_467), .Y(n_482) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_499), .B(n_527), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g528 ( .A(n_486), .Y(n_528) );
XNOR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_498), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .C(n_491), .D(n_493), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .C(n_497), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_499), .B(n_528), .Y(n_527) );
XNOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g501 ( .A(n_502), .B(n_516), .Y(n_501) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_505), .Y(n_653) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g588 ( .A(n_515), .Y(n_588) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
OAI21xp5_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_524), .Y(n_521) );
INVx1_ASAP7_75t_L g533 ( .A(n_530), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_602), .B1(n_620), .B2(n_621), .Y(n_535) );
INVx1_ASAP7_75t_L g621 ( .A(n_536), .Y(n_621) );
XNOR2xp5_ASAP7_75t_SL g536 ( .A(n_537), .B(n_579), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AO22x2_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_559), .B1(n_577), .B2(n_578), .Y(n_538) );
INVx1_ASAP7_75t_SL g578 ( .A(n_539), .Y(n_578) );
INVx1_ASAP7_75t_SL g558 ( .A(n_540), .Y(n_558) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_547), .Y(n_540) );
NAND4xp25_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .C(n_545), .D(n_546), .Y(n_541) );
NAND4xp25_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .C(n_553), .D(n_555), .Y(n_547) );
INVx2_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g678 ( .A(n_552), .Y(n_678) );
INVx3_ASAP7_75t_L g577 ( .A(n_559), .Y(n_577) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_563), .B(n_570), .Y(n_562) );
NAND4xp25_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .C(n_567), .D(n_568), .Y(n_563) );
INVx2_ASAP7_75t_L g693 ( .A(n_569), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .C(n_576), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_577), .A2(n_580), .B1(n_581), .B2(n_601), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_577), .Y(n_580) );
BUFx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g601 ( .A(n_582), .Y(n_601) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_592), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .C(n_589), .D(n_591), .Y(n_585) );
NAND4xp25_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .C(n_597), .D(n_599), .Y(n_592) );
INVx1_ASAP7_75t_L g620 ( .A(n_602), .Y(n_620) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
XNOR2x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_614), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .C(n_612), .Y(n_606) );
INVx1_ASAP7_75t_L g636 ( .A(n_609), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .C(n_618), .D(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_684), .B1(n_685), .B2(n_741), .Y(n_624) );
INVx1_ASAP7_75t_L g741 ( .A(n_625), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_657), .B2(n_683), .Y(n_625) );
INVx4_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_645), .Y(n_629) );
NAND4xp25_ASAP7_75t_SL g630 ( .A(n_631), .B(n_634), .C(n_637), .D(n_640), .Y(n_630) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .C(n_652), .D(n_655), .Y(n_645) );
BUFx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g683 ( .A(n_657), .Y(n_683) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_668), .B2(n_682), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_662), .B(n_669), .C(n_674), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_674), .Y(n_668) );
NAND4xp25_ASAP7_75t_SL g669 ( .A(n_670), .B(n_671), .C(n_672), .D(n_673), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .Y(n_674) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AO22x2_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_706), .B1(n_739), .B2(n_740), .Y(n_686) );
INVx1_ASAP7_75t_L g739 ( .A(n_687), .Y(n_739) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_697), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_694), .C(n_696), .Y(n_690) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .C(n_703), .D(n_704), .Y(n_697) );
BUFx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g740 ( .A(n_706), .Y(n_740) );
AO22x1_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_724), .B2(n_725), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g723 ( .A(n_710), .Y(n_723) );
NAND4xp75_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .C(n_717), .D(n_720), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g738 ( .A(n_726), .Y(n_738) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_732), .Y(n_726) );
NAND4xp25_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .C(n_730), .D(n_731), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .C(n_735), .D(n_736), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_748), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_745), .B(n_749), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g810 ( .A(n_747), .Y(n_810) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_760), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVxp67_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI222xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_786), .B1(n_788), .B2(n_805), .C1(n_806), .C2(n_809), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_764), .Y(n_785) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_774), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_781), .Y(n_774) );
OAI21xp5_ASAP7_75t_SL g775 ( .A1(n_776), .A2(n_777), .B(n_778), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
XOR2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_805), .Y(n_789) );
NOR2x1_ASAP7_75t_L g790 ( .A(n_791), .B(n_797), .Y(n_790) );
NAND4xp25_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .C(n_794), .D(n_796), .Y(n_791) );
NAND4xp25_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .C(n_800), .D(n_804), .Y(n_797) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
CKINVDCx6p67_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
endmodule