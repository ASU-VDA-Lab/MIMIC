module fake_netlist_6_3687_n_1652 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1652);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1652;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_78),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_6),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_38),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_87),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_16),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_8),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_108),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_36),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_92),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_35),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_86),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_94),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_141),
.Y(n_172)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_20),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_25),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_76),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_101),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_116),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_44),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_35),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_3),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_109),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_63),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_53),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_23),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_1),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_41),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_80),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_58),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_82),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_26),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_85),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_119),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_61),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_143),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_68),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_47),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_55),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_93),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_120),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_91),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_42),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_149),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_64),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_67),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_25),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_59),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_47),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_56),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_41),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_55),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_42),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_10),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_51),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_44),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_50),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_37),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_45),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_90),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_24),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_71),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_30),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_43),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_11),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_97),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_2),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_62),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_4),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_11),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_32),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_125),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_31),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_112),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_52),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_43),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_13),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_51),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_30),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_17),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_29),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_9),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_28),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_22),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_79),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_81),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_111),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_129),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_113),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_130),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_52),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_84),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_27),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_104),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_83),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_122),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_99),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_48),
.Y(n_275)
);

INVx4_ASAP7_75t_R g276 ( 
.A(n_140),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_32),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_37),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_2),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_121),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_147),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_49),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_22),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_24),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_5),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_49),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_60),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_12),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_20),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_57),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_96),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_146),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_18),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_21),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_33),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_153),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_151),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_204),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_234),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_0),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_206),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_234),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_152),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_158),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_234),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_155),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_180),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_160),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_163),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_234),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_234),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_233),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_170),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_256),
.B(n_294),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_168),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_171),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_240),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_154),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_154),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_246),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_172),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_175),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_287),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_260),
.B(n_3),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_176),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_180),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_181),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_181),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_177),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_198),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_198),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_226),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_162),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_226),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_159),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_239),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_178),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_248),
.B(n_5),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_277),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_277),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_239),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_185),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_186),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_164),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_168),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_187),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_194),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_190),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_197),
.Y(n_360)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_182),
.Y(n_361)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_195),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_199),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_203),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_190),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_192),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_278),
.B(n_6),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_165),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_248),
.B(n_7),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_192),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_205),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_159),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_209),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_218),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_210),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_183),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_218),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_161),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_220),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_296),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_322),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_353),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_332),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_299),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_354),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_299),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_298),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g393 ( 
.A(n_302),
.B(n_196),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

AND3x1_ASAP7_75t_L g395 ( 
.A(n_300),
.B(n_224),
.C(n_222),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_357),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_334),
.B(n_174),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_335),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_358),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_373),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_375),
.Y(n_405)
);

BUFx8_ASAP7_75t_L g406 ( 
.A(n_303),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_355),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_301),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_297),
.B(n_165),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_318),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_346),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_305),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_302),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_372),
.B(n_201),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_304),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_304),
.Y(n_421)
);

AND2x2_ASAP7_75t_SL g422 ( 
.A(n_331),
.B(n_157),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_307),
.B(n_201),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_318),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_307),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_376),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_306),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_308),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_308),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_303),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_311),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_311),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_312),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_313),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_368),
.B(n_294),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_317),
.B(n_211),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_314),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_320),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_315),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_328),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_315),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_321),
.B(n_196),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_336),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_316),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_366),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_329),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_333),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_323),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_370),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_336),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_362),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_157),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_415),
.B(n_337),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_422),
.A2(n_369),
.B1(n_349),
.B2(n_279),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_398),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_420),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_420),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_338),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_R g462 ( 
.A(n_409),
.B(n_361),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_377),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_420),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_422),
.B(n_310),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_348),
.Y(n_468)
);

BUFx10_ASAP7_75t_L g469 ( 
.A(n_427),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_430),
.B(n_166),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_423),
.B(n_360),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_424),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_430),
.B(n_423),
.Y(n_473)
);

BUFx4f_ASAP7_75t_L g474 ( 
.A(n_420),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_429),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_423),
.B(n_431),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_395),
.A2(n_367),
.B1(n_371),
.B2(n_380),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_R g478 ( 
.A(n_409),
.B(n_363),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_436),
.B(n_364),
.Y(n_479)
);

AND2x6_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_166),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_424),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_430),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_393),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_430),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_421),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_421),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_418),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_418),
.Y(n_489)
);

OR2x6_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_319),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_435),
.B(n_337),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_438),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_427),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_430),
.B(n_169),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_388),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_421),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_412),
.B(n_379),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_448),
.B(n_352),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_421),
.B(n_291),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_419),
.B(n_169),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_433),
.B(n_327),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_419),
.B(n_188),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_433),
.B(n_330),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_383),
.B(n_339),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_384),
.B(n_339),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_387),
.B(n_188),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_391),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_417),
.B(n_374),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

BUFx4f_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_442),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_425),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_389),
.A2(n_440),
.B1(n_428),
.B2(n_401),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_428),
.A2(n_251),
.B1(n_232),
.B2(n_245),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_382),
.B(n_378),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_385),
.B(n_340),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_442),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_387),
.B(n_241),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_440),
.B(n_167),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_387),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_444),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_394),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_444),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_387),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_387),
.B(n_241),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_434),
.B(n_213),
.Y(n_529)
);

BUFx4f_ASAP7_75t_L g530 ( 
.A(n_393),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_434),
.B(n_189),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_432),
.B(n_231),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_399),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_399),
.B(n_262),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_399),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_381),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_399),
.Y(n_537)
);

AND2x2_ASAP7_75t_SL g538 ( 
.A(n_447),
.B(n_262),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_444),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_444),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_397),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_399),
.B(n_271),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_402),
.B(n_340),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_403),
.B(n_222),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_432),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_439),
.B(n_191),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_407),
.B(n_271),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_403),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_408),
.A2(n_230),
.B1(n_295),
.B2(n_224),
.Y(n_550)
);

AND3x2_ASAP7_75t_L g551 ( 
.A(n_446),
.B(n_292),
.C(n_173),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_407),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_446),
.B(n_249),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_444),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_392),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_398),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_407),
.B(n_292),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_407),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_439),
.B(n_193),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_407),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_441),
.B(n_196),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_393),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_450),
.B(n_261),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_450),
.B(n_228),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_393),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_452),
.B(n_207),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_393),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_452),
.B(n_179),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_451),
.B(n_208),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_451),
.Y(n_570)
);

OAI21xp33_ASAP7_75t_SL g571 ( 
.A1(n_451),
.A2(n_200),
.B(n_179),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_443),
.Y(n_572)
);

INVx5_ASAP7_75t_L g573 ( 
.A(n_443),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_443),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_443),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_443),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_406),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_406),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_413),
.B(n_200),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_406),
.B(n_266),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_468),
.B(n_386),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_479),
.B(n_202),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_463),
.B(n_202),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_570),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_461),
.B(n_475),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_493),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_541),
.B(n_228),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_481),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_569),
.B(n_214),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_472),
.B(n_214),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_538),
.B(n_386),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_457),
.A2(n_237),
.B(n_244),
.C(n_227),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_466),
.B(n_212),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_L g595 ( 
.A(n_480),
.B(n_270),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_525),
.B(n_237),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_538),
.B(n_390),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_466),
.B(n_216),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_529),
.B(n_219),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_519),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_480),
.A2(n_280),
.B1(n_272),
.B2(n_281),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_570),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_454),
.B(n_221),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_485),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_454),
.B(n_223),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_549),
.B(n_265),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_476),
.A2(n_273),
.B(n_268),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_499),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_507),
.Y(n_609)
);

INVx8_ASAP7_75t_L g610 ( 
.A(n_578),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_507),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_480),
.A2(n_279),
.B1(n_232),
.B2(n_230),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_471),
.B(n_225),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_500),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_508),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_518),
.B(n_390),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_530),
.B(n_196),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_485),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_508),
.Y(n_619)
);

AOI221xp5_ASAP7_75t_L g620 ( 
.A1(n_550),
.A2(n_184),
.B1(n_275),
.B2(n_247),
.C(n_264),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_497),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_530),
.B(n_196),
.Y(n_622)
);

BUFx8_ASAP7_75t_L g623 ( 
.A(n_579),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_541),
.B(n_396),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_558),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_544),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_544),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_456),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_L g629 ( 
.A(n_480),
.B(n_503),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_480),
.B(n_290),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_491),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_491),
.B(n_217),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_510),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_456),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_488),
.B(n_217),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_453),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_490),
.B(n_396),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_512),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_455),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_480),
.A2(n_259),
.B1(n_243),
.B2(n_250),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_515),
.Y(n_642)
);

AOI221xp5_ASAP7_75t_L g643 ( 
.A1(n_531),
.A2(n_253),
.B1(n_250),
.B2(n_251),
.C(n_243),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_553),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_523),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_464),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_489),
.B(n_217),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_492),
.B(n_496),
.Y(n_648)
);

BUFx12f_ASAP7_75t_SL g649 ( 
.A(n_490),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_522),
.B(n_263),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_490),
.B(n_229),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_467),
.B(n_263),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_576),
.B(n_572),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_576),
.B(n_263),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_524),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_502),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_477),
.A2(n_580),
.B1(n_490),
.B2(n_503),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g658 ( 
.A(n_501),
.B(n_400),
.C(n_404),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_576),
.B(n_263),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_580),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_524),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_547),
.B(n_235),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_568),
.B(n_559),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_563),
.B(n_236),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_561),
.B(n_238),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_526),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_526),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_516),
.B(n_242),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_580),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_539),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_511),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_503),
.A2(n_426),
.B1(n_405),
.B2(n_449),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_540),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_540),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_568),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_460),
.B(n_465),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_511),
.B(n_252),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_465),
.B(n_255),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_511),
.B(n_258),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_554),
.Y(n_681)
);

BUFx8_ASAP7_75t_L g682 ( 
.A(n_536),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_511),
.B(n_254),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_545),
.B(n_341),
.Y(n_684)
);

BUFx8_ASAP7_75t_L g685 ( 
.A(n_536),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_SL g686 ( 
.A(n_578),
.B(n_445),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_486),
.B(n_514),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_566),
.B(n_284),
.Y(n_688)
);

BUFx6f_ASAP7_75t_SL g689 ( 
.A(n_469),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_469),
.B(n_289),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_514),
.B(n_293),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_514),
.B(n_341),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_469),
.B(n_161),
.Y(n_693)
);

NAND2x1p5_ASAP7_75t_L g694 ( 
.A(n_562),
.B(n_254),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_554),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_505),
.B(n_161),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_505),
.B(n_161),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_455),
.A2(n_286),
.B1(n_259),
.B2(n_267),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_581),
.B(n_269),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_527),
.Y(n_700)
);

AOI221xp5_ASAP7_75t_L g701 ( 
.A1(n_517),
.A2(n_286),
.B1(n_267),
.B2(n_282),
.C(n_285),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_545),
.B(n_564),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_494),
.B(n_269),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_545),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_473),
.A2(n_288),
.B1(n_282),
.B2(n_285),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_523),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_455),
.A2(n_295),
.B1(n_288),
.B2(n_257),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_572),
.B(n_269),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_533),
.B(n_351),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_494),
.B(n_545),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_527),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_527),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_503),
.B(n_257),
.Y(n_713)
);

AOI22x1_ASAP7_75t_L g714 ( 
.A1(n_575),
.A2(n_351),
.B1(n_350),
.B2(n_345),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_535),
.B(n_350),
.Y(n_715)
);

INVx11_ASAP7_75t_L g716 ( 
.A(n_682),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_682),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_688),
.A2(n_599),
.B(n_583),
.C(n_662),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_629),
.A2(n_513),
.B(n_474),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_644),
.B(n_504),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_608),
.B(n_506),
.Y(n_721)
);

AO21x1_ASAP7_75t_L g722 ( 
.A1(n_590),
.A2(n_495),
.B(n_470),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_640),
.A2(n_474),
.B(n_513),
.Y(n_723)
);

CKINVDCx6p67_ASAP7_75t_R g724 ( 
.A(n_689),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_599),
.B(n_482),
.Y(n_725)
);

INVx3_ASAP7_75t_SL g726 ( 
.A(n_683),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_640),
.A2(n_498),
.B(n_459),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_636),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_586),
.B(n_484),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_593),
.A2(n_571),
.B(n_564),
.C(n_542),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_688),
.B(n_503),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_685),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_663),
.A2(n_577),
.B1(n_574),
.B2(n_564),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_663),
.A2(n_455),
.B1(n_503),
.B2(n_478),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_657),
.A2(n_577),
.B1(n_574),
.B2(n_564),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_631),
.B(n_662),
.Y(n_736)
);

O2A1O1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_584),
.A2(n_542),
.B(n_521),
.C(n_557),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_600),
.B(n_483),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_612),
.A2(n_556),
.B1(n_458),
.B2(n_495),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_613),
.A2(n_455),
.B1(n_470),
.B2(n_462),
.Y(n_740)
);

CKINVDCx8_ASAP7_75t_R g741 ( 
.A(n_683),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_624),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_603),
.B(n_455),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_640),
.A2(n_498),
.B(n_459),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_656),
.A2(n_520),
.B(n_487),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_587),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_628),
.A2(n_509),
.B(n_521),
.C(n_557),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_645),
.A2(n_520),
.B(n_487),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_603),
.B(n_537),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_602),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_589),
.B(n_551),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_616),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_704),
.B(n_562),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_645),
.A2(n_487),
.B(n_560),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_653),
.A2(n_632),
.B(n_634),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_708),
.A2(n_548),
.B(n_534),
.C(n_509),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_685),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_602),
.Y(n_758)
);

O2A1O1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_708),
.A2(n_548),
.B(n_534),
.C(n_528),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_706),
.A2(n_487),
.B(n_560),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_676),
.A2(n_567),
.B1(n_565),
.B2(n_562),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_684),
.B(n_565),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_706),
.A2(n_558),
.B(n_560),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_612),
.A2(n_641),
.B1(n_643),
.B2(n_698),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_677),
.A2(n_687),
.B(n_713),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_605),
.B(n_555),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_625),
.A2(n_558),
.B(n_560),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_604),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_625),
.A2(n_558),
.B(n_532),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_692),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_605),
.B(n_537),
.Y(n_771)
);

NAND2x1p5_ASAP7_75t_L g772 ( 
.A(n_636),
.B(n_567),
.Y(n_772)
);

NOR2x1_ASAP7_75t_L g773 ( 
.A(n_592),
.B(n_537),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_595),
.A2(n_573),
.B(n_483),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_641),
.A2(n_567),
.B1(n_565),
.B2(n_343),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_587),
.B(n_573),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_613),
.B(n_626),
.Y(n_777)
);

CKINVDCx10_ASAP7_75t_R g778 ( 
.A(n_689),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_698),
.A2(n_565),
.B1(n_343),
.B2(n_344),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_594),
.A2(n_552),
.B1(n_528),
.B2(n_573),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_594),
.A2(n_552),
.B1(n_573),
.B2(n_483),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_642),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_598),
.A2(n_483),
.B1(n_345),
.B2(n_344),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_642),
.Y(n_784)
);

NOR3xp33_ASAP7_75t_L g785 ( 
.A(n_620),
.B(n_276),
.C(n_546),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_598),
.B(n_7),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_665),
.B(n_483),
.C(n_546),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_604),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_597),
.B(n_9),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_627),
.B(n_546),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_623),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_702),
.A2(n_543),
.B1(n_65),
.B2(n_69),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_654),
.A2(n_543),
.B(n_150),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_618),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_587),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_654),
.A2(n_543),
.B(n_144),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_582),
.Y(n_797)
);

NOR2xp67_ASAP7_75t_L g798 ( 
.A(n_673),
.B(n_142),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_630),
.A2(n_139),
.B(n_135),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_614),
.B(n_591),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_665),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_801)
);

AOI21xp33_ASAP7_75t_L g802 ( 
.A1(n_699),
.A2(n_697),
.B(n_696),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_648),
.A2(n_134),
.B(n_131),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_614),
.B(n_14),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_696),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_649),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_702),
.A2(n_127),
.B1(n_126),
.B2(n_123),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_636),
.B(n_106),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_617),
.A2(n_103),
.B(n_100),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_SL g810 ( 
.A(n_686),
.B(n_15),
.Y(n_810)
);

CKINVDCx10_ASAP7_75t_R g811 ( 
.A(n_683),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_609),
.B(n_19),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_651),
.B(n_19),
.Y(n_813)
);

AO32x1_ASAP7_75t_L g814 ( 
.A1(n_705),
.A2(n_695),
.A3(n_667),
.B1(n_671),
.B2(n_674),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_622),
.A2(n_98),
.B(n_89),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_638),
.Y(n_816)
);

AND2x2_ASAP7_75t_SL g817 ( 
.A(n_658),
.B(n_21),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_636),
.Y(n_818)
);

NAND2x1p5_ASAP7_75t_L g819 ( 
.A(n_587),
.B(n_72),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_679),
.A2(n_70),
.B(n_28),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_697),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_707),
.A2(n_56),
.B1(n_34),
.B2(n_36),
.Y(n_822)
);

AO22x1_ASAP7_75t_L g823 ( 
.A1(n_678),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_621),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_659),
.A2(n_611),
.B(n_615),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_619),
.B(n_40),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_655),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_651),
.B(n_46),
.Y(n_828)
);

OR2x6_ASAP7_75t_SL g829 ( 
.A(n_668),
.B(n_48),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_664),
.A2(n_54),
.B1(n_637),
.B2(n_646),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_684),
.B(n_670),
.Y(n_831)
);

OAI21xp33_ASAP7_75t_L g832 ( 
.A1(n_699),
.A2(n_680),
.B(n_678),
.Y(n_832)
);

AOI21x1_ASAP7_75t_L g833 ( 
.A1(n_659),
.A2(n_650),
.B(n_635),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_SL g834 ( 
.A(n_610),
.B(n_672),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_691),
.A2(n_709),
.B(n_715),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_655),
.Y(n_836)
);

OAI21xp5_ASAP7_75t_L g837 ( 
.A1(n_607),
.A2(n_633),
.B(n_639),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_700),
.A2(n_711),
.B(n_712),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_660),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_596),
.B(n_606),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_707),
.B(n_680),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_601),
.A2(n_674),
.B1(n_695),
.B2(n_669),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_647),
.A2(n_652),
.B(n_681),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_661),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_666),
.A2(n_681),
.B(n_667),
.C(n_669),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_666),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_675),
.B(n_694),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_690),
.B(n_703),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_588),
.B(n_693),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_694),
.B(n_588),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_610),
.A2(n_714),
.B(n_588),
.Y(n_851)
);

CKINVDCx10_ASAP7_75t_R g852 ( 
.A(n_623),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_701),
.B(n_610),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_612),
.A2(n_457),
.B1(n_641),
.B2(n_663),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_644),
.B(n_468),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_629),
.A2(n_513),
.B(n_474),
.Y(n_856)
);

AO22x1_ASAP7_75t_L g857 ( 
.A1(n_599),
.A2(n_662),
.B1(n_529),
.B2(n_598),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_663),
.B(n_538),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_631),
.B(n_481),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_583),
.A2(n_422),
.B1(n_688),
.B2(n_599),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_629),
.A2(n_513),
.B(n_474),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_670),
.B(n_624),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_663),
.B(n_538),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_629),
.A2(n_513),
.B(n_474),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_644),
.B(n_468),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_583),
.B(n_599),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_583),
.B(n_599),
.Y(n_867)
);

BUFx4f_ASAP7_75t_L g868 ( 
.A(n_710),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_585),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_636),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_653),
.A2(n_593),
.B(n_461),
.Y(n_871)
);

OAI21xp33_ASAP7_75t_L g872 ( 
.A1(n_599),
.A2(n_643),
.B(n_605),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_653),
.A2(n_593),
.B(n_461),
.Y(n_873)
);

AO31x2_ASAP7_75t_L g874 ( 
.A1(n_722),
.A2(n_718),
.A3(n_786),
.B(n_842),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_794),
.Y(n_875)
);

BUFx6f_ASAP7_75t_SL g876 ( 
.A(n_717),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_866),
.B(n_867),
.Y(n_877)
);

AO31x2_ASAP7_75t_L g878 ( 
.A1(n_735),
.A2(n_854),
.A3(n_733),
.B(n_845),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_765),
.A2(n_864),
.B(n_861),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_728),
.Y(n_880)
);

NAND2x1_ASAP7_75t_L g881 ( 
.A(n_728),
.B(n_818),
.Y(n_881)
);

AOI21x1_ASAP7_75t_L g882 ( 
.A1(n_749),
.A2(n_771),
.B(n_833),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_838),
.A2(n_769),
.B(n_837),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_742),
.B(n_797),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_743),
.A2(n_835),
.B(n_723),
.Y(n_885)
);

BUFx12f_ASAP7_75t_L g886 ( 
.A(n_806),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_800),
.A2(n_774),
.B(n_840),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_860),
.A2(n_854),
.B1(n_764),
.B2(n_872),
.Y(n_888)
);

NAND3xp33_ASAP7_75t_L g889 ( 
.A(n_802),
.B(n_857),
.C(n_828),
.Y(n_889)
);

OAI21x1_ASAP7_75t_L g890 ( 
.A1(n_754),
.A2(n_763),
.B(n_760),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_SL g891 ( 
.A1(n_734),
.A2(n_764),
.B(n_858),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_777),
.B(n_770),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_716),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_727),
.A2(n_744),
.B(n_847),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_729),
.B(n_725),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_750),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_752),
.Y(n_897)
);

BUFx12f_ASAP7_75t_L g898 ( 
.A(n_791),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_745),
.A2(n_748),
.B(n_755),
.Y(n_899)
);

INVx4_ASAP7_75t_L g900 ( 
.A(n_728),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_813),
.A2(n_863),
.B(n_841),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_873),
.A2(n_871),
.B(n_755),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_797),
.B(n_742),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_818),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_721),
.B(n_736),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_873),
.A2(n_825),
.B(n_730),
.Y(n_906)
);

AO21x2_ASAP7_75t_L g907 ( 
.A1(n_825),
.A2(n_740),
.B(n_851),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_832),
.B(n_855),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_859),
.B(n_831),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_805),
.A2(n_789),
.B1(n_830),
.B2(n_821),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_812),
.A2(n_826),
.B1(n_822),
.B2(n_853),
.Y(n_911)
);

INVx8_ASAP7_75t_L g912 ( 
.A(n_862),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_720),
.B(n_848),
.Y(n_913)
);

OR2x2_ASAP7_75t_L g914 ( 
.A(n_816),
.B(n_839),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_870),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_782),
.B(n_784),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_870),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_767),
.A2(n_747),
.B(n_759),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_758),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_737),
.A2(n_756),
.B(n_785),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_768),
.B(n_788),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_844),
.A2(n_846),
.B(n_804),
.Y(n_922)
);

OAI21x1_ASAP7_75t_L g923 ( 
.A1(n_827),
.A2(n_836),
.B(n_869),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_818),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_816),
.B(n_839),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_793),
.A2(n_796),
.B(n_824),
.Y(n_926)
);

OAI21x1_ASAP7_75t_SL g927 ( 
.A1(n_793),
.A2(n_796),
.B(n_799),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_781),
.A2(n_780),
.B(n_787),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_827),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_761),
.A2(n_790),
.B(n_762),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_865),
.B(n_766),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_836),
.A2(n_772),
.B(n_773),
.Y(n_932)
);

AOI21x1_ASAP7_75t_SL g933 ( 
.A1(n_850),
.A2(n_753),
.B(n_849),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_868),
.A2(n_798),
.B1(n_801),
.B2(n_817),
.Y(n_934)
);

NAND2x1p5_ASAP7_75t_L g935 ( 
.A(n_870),
.B(n_762),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_772),
.A2(n_776),
.B(n_795),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_SL g937 ( 
.A1(n_775),
.A2(n_819),
.B(n_792),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_859),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_738),
.A2(n_795),
.B(n_746),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_753),
.B(n_831),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_862),
.Y(n_941)
);

AOI21xp33_ASAP7_75t_L g942 ( 
.A1(n_810),
.A2(n_739),
.B(n_862),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_868),
.B(n_751),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_808),
.A2(n_775),
.B(n_809),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_815),
.A2(n_783),
.B(n_803),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_834),
.A2(n_814),
.B(n_779),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_726),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_819),
.A2(n_820),
.B(n_807),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_779),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_732),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_739),
.A2(n_810),
.B(n_834),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_814),
.A2(n_751),
.B(n_823),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_814),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_741),
.B(n_757),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_829),
.A2(n_811),
.B(n_724),
.C(n_778),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_852),
.B(n_866),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_866),
.B(n_867),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_721),
.B(n_872),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_742),
.B(n_797),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_960)
);

AO31x2_ASAP7_75t_L g961 ( 
.A1(n_722),
.A2(n_718),
.A3(n_786),
.B(n_842),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_872),
.A2(n_718),
.B(n_802),
.C(n_786),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_742),
.B(n_797),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_794),
.Y(n_965)
);

OAI21x1_ASAP7_75t_SL g966 ( 
.A1(n_825),
.A2(n_871),
.B(n_873),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_866),
.B(n_867),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_728),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_794),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_718),
.A2(n_872),
.B(n_871),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_728),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_794),
.Y(n_972)
);

AOI21x1_ASAP7_75t_L g973 ( 
.A1(n_749),
.A2(n_771),
.B(n_843),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_859),
.B(n_831),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_866),
.B(n_867),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_860),
.A2(n_854),
.B1(n_764),
.B2(n_718),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_872),
.A2(n_718),
.B(n_802),
.C(n_786),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_718),
.A2(n_872),
.B(n_871),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_872),
.A2(n_718),
.B(n_802),
.C(n_786),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_718),
.A2(n_872),
.B(n_871),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_866),
.B(n_867),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_718),
.A2(n_872),
.B(n_871),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_731),
.A2(n_640),
.B(n_629),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_L g991 ( 
.A(n_718),
.B(n_860),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_862),
.B(n_717),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_742),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_731),
.A2(n_640),
.B(n_629),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_866),
.B(n_867),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_716),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_718),
.A2(n_872),
.B(n_871),
.Y(n_998)
);

OAI21x1_ASAP7_75t_SL g999 ( 
.A1(n_825),
.A2(n_871),
.B(n_873),
.Y(n_999)
);

AO31x2_ASAP7_75t_L g1000 ( 
.A1(n_722),
.A2(n_718),
.A3(n_786),
.B(n_842),
.Y(n_1000)
);

AO31x2_ASAP7_75t_L g1001 ( 
.A1(n_722),
.A2(n_718),
.A3(n_786),
.B(n_842),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_L g1002 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_1002)
);

NAND2x1_ASAP7_75t_L g1003 ( 
.A(n_728),
.B(n_636),
.Y(n_1003)
);

AOI21x1_ASAP7_75t_L g1004 ( 
.A1(n_749),
.A2(n_771),
.B(n_843),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_765),
.A2(n_856),
.B(n_719),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_SL g1006 ( 
.A1(n_825),
.A2(n_871),
.B(n_873),
.Y(n_1006)
);

BUFx12f_ASAP7_75t_L g1007 ( 
.A(n_806),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_866),
.B(n_867),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_915),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_884),
.Y(n_1010)
);

AO32x2_ASAP7_75t_L g1011 ( 
.A1(n_978),
.A2(n_888),
.A3(n_910),
.B1(n_911),
.B2(n_934),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_887),
.A2(n_991),
.B(n_885),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_875),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_935),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_958),
.B(n_967),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_915),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_959),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_903),
.B(n_877),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_909),
.B(n_974),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_898),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_993),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_877),
.B(n_957),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_963),
.B(n_931),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_957),
.B(n_975),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_975),
.B(n_1008),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_909),
.B(n_974),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_914),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_L g1028 ( 
.A(n_962),
.B(n_980),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1008),
.B(n_925),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_920),
.A2(n_995),
.B(n_988),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_896),
.Y(n_1031)
);

AO21x1_ASAP7_75t_L g1032 ( 
.A1(n_978),
.A2(n_888),
.B(n_982),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_892),
.B(n_895),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_993),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_912),
.B(n_992),
.Y(n_1035)
);

OR2x6_ASAP7_75t_L g1036 ( 
.A(n_912),
.B(n_992),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_943),
.B(n_938),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_892),
.B(n_895),
.Y(n_1038)
);

BUFx2_ASAP7_75t_SL g1039 ( 
.A(n_876),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_983),
.A2(n_889),
.B(n_989),
.C(n_982),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_970),
.A2(n_998),
.B(n_986),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_924),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_919),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_905),
.B(n_970),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_986),
.A2(n_998),
.B(n_989),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_951),
.A2(n_910),
.B1(n_949),
.B2(n_906),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_911),
.B(n_908),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_SL g1048 ( 
.A(n_951),
.B(n_942),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_901),
.B(n_916),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_965),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_897),
.B(n_956),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_916),
.B(n_969),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_942),
.A2(n_934),
.B1(n_913),
.B2(n_912),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_SL g1054 ( 
.A1(n_927),
.A2(n_941),
.B1(n_947),
.B2(n_876),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_940),
.B(n_941),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_972),
.B(n_891),
.Y(n_1056)
);

INVx5_ASAP7_75t_L g1057 ( 
.A(n_915),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_917),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_947),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_941),
.B(n_992),
.Y(n_1060)
);

AOI21xp33_ASAP7_75t_SL g1061 ( 
.A1(n_954),
.A2(n_955),
.B(n_940),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_906),
.A2(n_966),
.B1(n_999),
.B2(n_1006),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_917),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_929),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_937),
.A2(n_902),
.B1(n_926),
.B2(n_944),
.Y(n_1065)
);

CKINVDCx8_ASAP7_75t_R g1066 ( 
.A(n_893),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_886),
.Y(n_1067)
);

BUFx12f_ASAP7_75t_L g1068 ( 
.A(n_996),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_878),
.B(n_921),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_968),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_1007),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_950),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_935),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_946),
.A2(n_918),
.B(n_928),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_SL g1075 ( 
.A1(n_928),
.A2(n_945),
.B(n_930),
.C(n_894),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_948),
.A2(n_899),
.B(n_990),
.C(n_994),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_924),
.B(n_900),
.Y(n_1077)
);

CKINVDCx6p67_ASAP7_75t_R g1078 ( 
.A(n_924),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_968),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_879),
.A2(n_960),
.B(n_1002),
.Y(n_1080)
);

OAI21xp33_ASAP7_75t_SL g1081 ( 
.A1(n_923),
.A2(n_932),
.B(n_936),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_971),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_880),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_924),
.B(n_900),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_880),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_904),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_881),
.B(n_1003),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_904),
.B(n_874),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_907),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_L g1090 ( 
.A(n_939),
.B(n_933),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_878),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_874),
.B(n_1000),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_878),
.B(n_874),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_953),
.Y(n_1094)
);

CKINVDCx6p67_ASAP7_75t_R g1095 ( 
.A(n_922),
.Y(n_1095)
);

AOI21x1_ASAP7_75t_L g1096 ( 
.A1(n_973),
.A2(n_1004),
.B(n_882),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_883),
.B(n_979),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_964),
.A2(n_981),
.B(n_997),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_961),
.B(n_1001),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_961),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1000),
.B(n_1001),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1000),
.B(n_1001),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_890),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_976),
.B(n_977),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_984),
.B(n_985),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_987),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_1005),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_897),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_877),
.B(n_957),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_962),
.A2(n_802),
.B(n_872),
.C(n_718),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_950),
.Y(n_1111)
);

BUFx12f_ASAP7_75t_L g1112 ( 
.A(n_898),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_915),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_886),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_877),
.A2(n_975),
.B1(n_1008),
.B2(n_957),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_875),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_931),
.B(n_797),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_931),
.B(n_797),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_993),
.Y(n_1119)
);

INVxp67_ASAP7_75t_L g1120 ( 
.A(n_897),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_909),
.B(n_974),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_886),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_875),
.Y(n_1123)
);

AOI222xp33_ASAP7_75t_L g1124 ( 
.A1(n_888),
.A2(n_643),
.B1(n_872),
.B2(n_958),
.C1(n_978),
.C2(n_764),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_915),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_877),
.B(n_957),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_914),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_935),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_935),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_SL g1130 ( 
.A1(n_958),
.A2(n_817),
.B1(n_398),
.B2(n_536),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_884),
.B(n_959),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_884),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_884),
.B(n_959),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_877),
.B(n_957),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_884),
.Y(n_1135)
);

OAI21xp33_ASAP7_75t_L g1136 ( 
.A1(n_958),
.A2(n_872),
.B(n_599),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_958),
.A2(n_872),
.B(n_802),
.C(n_718),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_912),
.B(n_992),
.Y(n_1138)
);

NOR2x1_ASAP7_75t_SL g1139 ( 
.A(n_924),
.B(n_728),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_909),
.B(n_974),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_875),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_903),
.B(n_797),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_914),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_877),
.A2(n_975),
.B1(n_1008),
.B2(n_957),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_903),
.B(n_797),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_875),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1015),
.A2(n_1109),
.B1(n_1134),
.B2(n_1022),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1019),
.B(n_1026),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1034),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1130),
.A2(n_1136),
.B1(n_1124),
.B2(n_1048),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1013),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1057),
.Y(n_1152)
);

BUFx2_ASAP7_75t_R g1153 ( 
.A(n_1066),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1031),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1043),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1124),
.A2(n_1028),
.B1(n_1032),
.B2(n_1046),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_1027),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1017),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1046),
.A2(n_1048),
.B1(n_1047),
.B2(n_1065),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1022),
.A2(n_1134),
.B1(n_1126),
.B2(n_1025),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_1042),
.B(n_1070),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1050),
.Y(n_1162)
);

NAND2x1p5_ASAP7_75t_L g1163 ( 
.A(n_1042),
.B(n_1070),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_SL g1164 ( 
.A1(n_1065),
.A2(n_1023),
.B1(n_1033),
.B2(n_1038),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_1072),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1047),
.A2(n_1115),
.B1(n_1144),
.B2(n_1030),
.Y(n_1166)
);

CKINVDCx11_ASAP7_75t_R g1167 ( 
.A(n_1111),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1077),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1116),
.Y(n_1169)
);

OAI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_1033),
.A2(n_1038),
.B1(n_1024),
.B2(n_1025),
.Y(n_1170)
);

CKINVDCx12_ASAP7_75t_R g1171 ( 
.A(n_1035),
.Y(n_1171)
);

AOI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1096),
.A2(n_1097),
.B(n_1045),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1059),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1115),
.A2(n_1144),
.B1(n_1041),
.B2(n_1109),
.Y(n_1174)
);

INVx2_ASAP7_75t_SL g1175 ( 
.A(n_1127),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1123),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1019),
.B(n_1026),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1117),
.A2(n_1118),
.B1(n_1053),
.B2(n_1037),
.Y(n_1178)
);

AND2x6_ASAP7_75t_L g1179 ( 
.A(n_1088),
.B(n_1056),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_SL g1180 ( 
.A1(n_1024),
.A2(n_1126),
.B1(n_1132),
.B2(n_1135),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1094),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1141),
.Y(n_1182)
);

AO21x1_ASAP7_75t_L g1183 ( 
.A1(n_1110),
.A2(n_1049),
.B(n_1056),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1146),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1062),
.A2(n_1044),
.B1(n_1010),
.B2(n_1133),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1137),
.A2(n_1029),
.B1(n_1018),
.B2(n_1108),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1071),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1131),
.B(n_1142),
.Y(n_1188)
);

CKINVDCx11_ASAP7_75t_R g1189 ( 
.A(n_1020),
.Y(n_1189)
);

AO21x2_ASAP7_75t_L g1190 ( 
.A1(n_1080),
.A2(n_1098),
.B(n_1012),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_1143),
.Y(n_1191)
);

BUFx12f_ASAP7_75t_L g1192 ( 
.A(n_1112),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_SL g1193 ( 
.A1(n_1039),
.A2(n_1037),
.B1(n_1060),
.B2(n_1119),
.Y(n_1193)
);

INVx6_ASAP7_75t_SL g1194 ( 
.A(n_1035),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1120),
.Y(n_1195)
);

CKINVDCx11_ASAP7_75t_R g1196 ( 
.A(n_1068),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_1070),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1040),
.A2(n_1052),
.B1(n_1119),
.B2(n_1021),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1052),
.A2(n_1021),
.B1(n_1051),
.B2(n_1145),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1094),
.Y(n_1200)
);

INVx11_ASAP7_75t_L g1201 ( 
.A(n_1107),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1044),
.A2(n_1054),
.B1(n_1035),
.B2(n_1138),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_L g1203 ( 
.A(n_1067),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1121),
.B(n_1140),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1060),
.A2(n_1055),
.B1(n_1138),
.B2(n_1036),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_1114),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1091),
.A2(n_1049),
.B1(n_1074),
.B2(n_1011),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1011),
.A2(n_1036),
.B1(n_1138),
.B2(n_1074),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1064),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1083),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1069),
.Y(n_1211)
);

INVx2_ASAP7_75t_SL g1212 ( 
.A(n_1122),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1085),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1036),
.A2(n_1061),
.B1(n_1095),
.B2(n_1069),
.Y(n_1214)
);

BUFx4f_ASAP7_75t_SL g1215 ( 
.A(n_1078),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1113),
.Y(n_1216)
);

AO21x1_ASAP7_75t_SL g1217 ( 
.A1(n_1100),
.A2(n_1093),
.B(n_1099),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1063),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1077),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1075),
.A2(n_1105),
.B(n_1104),
.Y(n_1220)
);

INVx6_ASAP7_75t_L g1221 ( 
.A(n_1084),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1014),
.B(n_1128),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1011),
.Y(n_1223)
);

BUFx8_ASAP7_75t_SL g1224 ( 
.A(n_1009),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1092),
.A2(n_1101),
.B(n_1102),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1014),
.B(n_1129),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1103),
.A2(n_1139),
.B1(n_1129),
.B2(n_1128),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1073),
.A2(n_1090),
.B1(n_1106),
.B2(n_1082),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1079),
.A2(n_1073),
.B1(n_1089),
.B2(n_1086),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1087),
.A2(n_1009),
.B1(n_1016),
.B2(n_1058),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1009),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1016),
.B(n_1058),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1125),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1087),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1076),
.A2(n_1081),
.B(n_1125),
.Y(n_1235)
);

CKINVDCx11_ASAP7_75t_R g1236 ( 
.A(n_1072),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1057),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1130),
.A2(n_817),
.B1(n_958),
.B2(n_398),
.Y(n_1238)
);

BUFx2_ASAP7_75t_R g1239 ( 
.A(n_1066),
.Y(n_1239)
);

INVx5_ASAP7_75t_L g1240 ( 
.A(n_1042),
.Y(n_1240)
);

CKINVDCx11_ASAP7_75t_R g1241 ( 
.A(n_1072),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1124),
.A2(n_872),
.B1(n_958),
.B2(n_1136),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1023),
.B(n_1131),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1057),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1124),
.A2(n_872),
.B1(n_958),
.B2(n_1136),
.Y(n_1245)
);

AND2x2_ASAP7_75t_SL g1246 ( 
.A(n_1028),
.B(n_991),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1023),
.B(n_1131),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1015),
.B(n_967),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1124),
.A2(n_872),
.B1(n_958),
.B2(n_1136),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1023),
.B(n_1131),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1034),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1130),
.A2(n_872),
.B1(n_390),
.B2(n_396),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1034),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1137),
.A2(n_718),
.B(n_802),
.Y(n_1254)
);

INVx8_ASAP7_75t_L g1255 ( 
.A(n_1057),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_SL g1256 ( 
.A1(n_1053),
.A2(n_951),
.B(n_952),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1225),
.B(n_1211),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1211),
.B(n_1208),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1147),
.B(n_1160),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1223),
.B(n_1207),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1149),
.Y(n_1261)
);

INVx11_ASAP7_75t_L g1262 ( 
.A(n_1206),
.Y(n_1262)
);

HB1xp67_ASAP7_75t_L g1263 ( 
.A(n_1149),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1223),
.B(n_1207),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1251),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1170),
.B(n_1174),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1235),
.Y(n_1267)
);

NOR2x1_ASAP7_75t_SL g1268 ( 
.A(n_1217),
.B(n_1214),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1235),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1183),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1181),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1251),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1220),
.A2(n_1254),
.B(n_1166),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1235),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1234),
.B(n_1205),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1238),
.A2(n_1246),
.B1(n_1256),
.B2(n_1202),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1181),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1248),
.B(n_1243),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1172),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1166),
.A2(n_1159),
.B(n_1174),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1190),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1159),
.B(n_1200),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1200),
.B(n_1186),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1253),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1156),
.A2(n_1185),
.B(n_1242),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1198),
.B(n_1185),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1234),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1164),
.B(n_1156),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1247),
.B(n_1250),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1150),
.A2(n_1229),
.B(n_1176),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1179),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1158),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1242),
.A2(n_1249),
.B1(n_1245),
.B2(n_1246),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1245),
.A2(n_1249),
.B(n_1155),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1199),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1151),
.A2(n_1162),
.B(n_1154),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_1195),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1169),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1182),
.B(n_1184),
.Y(n_1299)
);

AO21x2_ASAP7_75t_L g1300 ( 
.A1(n_1178),
.A2(n_1213),
.B(n_1210),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1179),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1179),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1173),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1188),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1252),
.A2(n_1180),
.B1(n_1194),
.B2(n_1193),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1167),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1157),
.Y(n_1307)
);

INVx5_ASAP7_75t_SL g1308 ( 
.A(n_1201),
.Y(n_1308)
);

NOR2x1_ASAP7_75t_SL g1309 ( 
.A(n_1240),
.B(n_1244),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1255),
.Y(n_1310)
);

AO21x2_ASAP7_75t_L g1311 ( 
.A1(n_1222),
.A2(n_1226),
.B(n_1209),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1171),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1168),
.B(n_1219),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1255),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1230),
.A2(n_1161),
.B(n_1163),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1175),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1194),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1194),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1228),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1191),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1167),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1227),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1148),
.B(n_1177),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1152),
.A2(n_1216),
.B(n_1237),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1218),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1232),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1260),
.B(n_1231),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1311),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1257),
.B(n_1231),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1259),
.B(n_1231),
.Y(n_1330)
);

AOI222xp33_ASAP7_75t_L g1331 ( 
.A1(n_1288),
.A2(n_1189),
.B1(n_1241),
.B2(n_1236),
.C1(n_1192),
.C2(n_1196),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1259),
.B(n_1197),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1271),
.B(n_1216),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1271),
.B(n_1197),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1293),
.A2(n_1241),
.B1(n_1236),
.B2(n_1204),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1296),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1296),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1291),
.B(n_1233),
.Y(n_1338)
);

INVx5_ASAP7_75t_L g1339 ( 
.A(n_1279),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1301),
.B(n_1302),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1311),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1315),
.Y(n_1342)
);

NAND4xp25_ASAP7_75t_L g1343 ( 
.A(n_1293),
.B(n_1153),
.C(n_1239),
.D(n_1189),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1311),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1296),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1315),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1287),
.B(n_1212),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1298),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1267),
.B(n_1221),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1269),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1281),
.A2(n_1165),
.B(n_1224),
.Y(n_1351)
);

AND2x4_ASAP7_75t_SL g1352 ( 
.A(n_1275),
.B(n_1187),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1260),
.B(n_1203),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1277),
.B(n_1215),
.Y(n_1354)
);

AND2x4_ASAP7_75t_SL g1355 ( 
.A(n_1275),
.B(n_1196),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1274),
.B(n_1206),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1300),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1300),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1264),
.B(n_1258),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1264),
.B(n_1258),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1300),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1295),
.B(n_1270),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1335),
.A2(n_1276),
.B1(n_1286),
.B2(n_1288),
.Y(n_1363)
);

OAI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1335),
.A2(n_1343),
.B1(n_1331),
.B2(n_1305),
.C(n_1266),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1359),
.B(n_1304),
.Y(n_1365)
);

NAND2xp33_ASAP7_75t_SL g1366 ( 
.A(n_1338),
.B(n_1306),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1343),
.B(n_1278),
.Y(n_1367)
);

AOI221xp5_ASAP7_75t_L g1368 ( 
.A1(n_1332),
.A2(n_1266),
.B1(n_1362),
.B2(n_1304),
.C(n_1322),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1360),
.B(n_1261),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1360),
.B(n_1263),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1348),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_R g1372 ( 
.A(n_1353),
.B(n_1321),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1332),
.A2(n_1286),
.B1(n_1322),
.B2(n_1285),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1331),
.B(n_1313),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1362),
.B(n_1265),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1355),
.A2(n_1319),
.B(n_1352),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1330),
.B(n_1272),
.Y(n_1377)
);

AOI221xp5_ASAP7_75t_L g1378 ( 
.A1(n_1357),
.A2(n_1297),
.B1(n_1319),
.B2(n_1284),
.C(n_1307),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1353),
.A2(n_1285),
.B1(n_1280),
.B2(n_1283),
.Y(n_1379)
);

OAI221xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1353),
.A2(n_1283),
.B1(n_1282),
.B2(n_1324),
.C(n_1312),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1329),
.B(n_1273),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1355),
.A2(n_1282),
.B(n_1323),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1357),
.B(n_1285),
.C(n_1280),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1329),
.B(n_1268),
.Y(n_1384)
);

NAND3xp33_ASAP7_75t_L g1385 ( 
.A(n_1358),
.B(n_1285),
.C(n_1280),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1354),
.A2(n_1280),
.B1(n_1292),
.B2(n_1275),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1356),
.B(n_1326),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1356),
.B(n_1326),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1356),
.B(n_1300),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1333),
.B(n_1290),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1333),
.B(n_1290),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1334),
.B(n_1290),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_1355),
.B(n_1313),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1354),
.B(n_1289),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1358),
.B(n_1325),
.C(n_1361),
.Y(n_1395)
);

OAI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1342),
.A2(n_1318),
.B1(n_1317),
.B2(n_1324),
.C(n_1292),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1334),
.B(n_1290),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1340),
.B(n_1279),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1352),
.A2(n_1292),
.B1(n_1308),
.B2(n_1294),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1340),
.B(n_1299),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1352),
.A2(n_1308),
.B1(n_1294),
.B2(n_1317),
.Y(n_1401)
);

OAI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1342),
.A2(n_1317),
.B1(n_1318),
.B2(n_1303),
.C(n_1316),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_SL g1403 ( 
.A1(n_1351),
.A2(n_1309),
.B(n_1294),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1349),
.B(n_1299),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1398),
.B(n_1346),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1390),
.B(n_1336),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1371),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1391),
.B(n_1336),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1371),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1398),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1381),
.B(n_1346),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1392),
.B(n_1328),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1400),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1381),
.B(n_1346),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1397),
.B(n_1328),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1375),
.B(n_1341),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1404),
.Y(n_1417)
);

INVx5_ASAP7_75t_L g1418 ( 
.A(n_1384),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1395),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1384),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1365),
.B(n_1341),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1395),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1367),
.B(n_1347),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1389),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1369),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1370),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1383),
.B(n_1339),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1386),
.B(n_1350),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1377),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1364),
.A2(n_1294),
.B1(n_1327),
.B2(n_1351),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1373),
.B(n_1344),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1409),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1412),
.B(n_1387),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1406),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1410),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1418),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1412),
.B(n_1388),
.Y(n_1437)
);

AND2x4_ASAP7_75t_SL g1438 ( 
.A(n_1427),
.B(n_1338),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1410),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1410),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1406),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1418),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1418),
.B(n_1394),
.Y(n_1443)
);

OAI21xp33_ASAP7_75t_L g1444 ( 
.A1(n_1431),
.A2(n_1363),
.B(n_1368),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1427),
.B(n_1403),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1409),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1418),
.B(n_1351),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1418),
.B(n_1393),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1410),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1418),
.B(n_1337),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1407),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1423),
.B(n_1374),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1419),
.B(n_1422),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1407),
.Y(n_1454)
);

NOR2x1p5_ASAP7_75t_SL g1455 ( 
.A(n_1419),
.B(n_1345),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1418),
.B(n_1351),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1422),
.B(n_1378),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1418),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1429),
.B(n_1425),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1427),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1420),
.B(n_1351),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1413),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1415),
.B(n_1383),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1417),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1415),
.B(n_1385),
.Y(n_1465)
);

OAI21xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1420),
.A2(n_1403),
.B(n_1402),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1427),
.B(n_1345),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1431),
.B(n_1385),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1417),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1429),
.B(n_1344),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1451),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1458),
.B(n_1427),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1451),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1435),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1444),
.B(n_1423),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1444),
.B(n_1425),
.Y(n_1476)
);

AOI32xp33_ASAP7_75t_L g1477 ( 
.A1(n_1457),
.A2(n_1363),
.A3(n_1430),
.B1(n_1428),
.B2(n_1366),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1457),
.B(n_1426),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1453),
.B(n_1426),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1453),
.B(n_1406),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1452),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1451),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1438),
.B(n_1424),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1454),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1466),
.A2(n_1430),
.B1(n_1382),
.B2(n_1376),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1459),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1438),
.B(n_1424),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1454),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1468),
.B(n_1424),
.Y(n_1489)
);

AO221x1_ASAP7_75t_L g1490 ( 
.A1(n_1442),
.A2(n_1399),
.B1(n_1401),
.B2(n_1424),
.C(n_1379),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1438),
.B(n_1443),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1454),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1433),
.B(n_1262),
.Y(n_1493)
);

OAI311xp33_ASAP7_75t_L g1494 ( 
.A1(n_1466),
.A2(n_1396),
.A3(n_1376),
.B1(n_1382),
.C1(n_1408),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1432),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1443),
.B(n_1424),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1460),
.B(n_1411),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1468),
.B(n_1416),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1432),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1460),
.B(n_1411),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1446),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1458),
.B(n_1405),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1435),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1460),
.B(n_1411),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1458),
.B(n_1405),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1435),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1446),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1448),
.B(n_1414),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1433),
.B(n_1416),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1437),
.B(n_1421),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1459),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1439),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1462),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1474),
.Y(n_1514)
);

NOR2x1_ASAP7_75t_L g1515 ( 
.A(n_1476),
.B(n_1458),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1481),
.B(n_1437),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1475),
.B(n_1463),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1491),
.B(n_1442),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1474),
.A2(n_1456),
.B(n_1447),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1478),
.B(n_1463),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1477),
.B(n_1465),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1491),
.B(n_1436),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1493),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1495),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1472),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1498),
.B(n_1262),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1490),
.A2(n_1372),
.B1(n_1428),
.B2(n_1448),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1508),
.B(n_1436),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1508),
.B(n_1436),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1477),
.B(n_1448),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1485),
.A2(n_1380),
.B1(n_1448),
.B2(n_1445),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1490),
.A2(n_1428),
.B1(n_1465),
.B2(n_1338),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1499),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1486),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1513),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1511),
.B(n_1434),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1509),
.A2(n_1445),
.B1(n_1417),
.B2(n_1461),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1497),
.B(n_1445),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1502),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1494),
.A2(n_1445),
.B1(n_1456),
.B2(n_1447),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1513),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1497),
.B(n_1500),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1479),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1501),
.Y(n_1545)
);

INVx1_ASAP7_75t_SL g1546 ( 
.A(n_1500),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1501),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1480),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1507),
.Y(n_1549)
);

OAI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1541),
.A2(n_1445),
.B1(n_1489),
.B2(n_1480),
.C(n_1507),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1535),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1543),
.B(n_1504),
.Y(n_1552)
);

OAI32xp33_ASAP7_75t_L g1553 ( 
.A1(n_1521),
.A2(n_1533),
.A3(n_1530),
.B1(n_1517),
.B2(n_1534),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1524),
.B(n_1510),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1546),
.B(n_1504),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1516),
.B(n_1434),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1533),
.B(n_1441),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1535),
.Y(n_1558)
);

AOI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1527),
.A2(n_1472),
.B1(n_1441),
.B2(n_1502),
.C(n_1505),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1543),
.B(n_1502),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1532),
.A2(n_1445),
.B1(n_1502),
.B2(n_1505),
.Y(n_1561)
);

NAND2x1_ASAP7_75t_SL g1562 ( 
.A(n_1515),
.B(n_1532),
.Y(n_1562)
);

OAI32xp33_ASAP7_75t_L g1563 ( 
.A1(n_1531),
.A2(n_1483),
.A3(n_1487),
.B1(n_1496),
.B2(n_1461),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1542),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1548),
.B(n_1496),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1544),
.B(n_1462),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1542),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1545),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1540),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1525),
.Y(n_1570)
);

NOR4xp25_ASAP7_75t_SL g1571 ( 
.A(n_1540),
.B(n_1484),
.C(n_1488),
.D(n_1471),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1518),
.B(n_1505),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1520),
.B(n_1483),
.Y(n_1573)
);

OAI31xp33_ASAP7_75t_L g1574 ( 
.A1(n_1537),
.A2(n_1472),
.A3(n_1505),
.B(n_1487),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1528),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1559),
.B(n_1570),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1555),
.B(n_1536),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1569),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1572),
.B(n_1552),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1565),
.B(n_1549),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1552),
.B(n_1523),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1569),
.B(n_1549),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1557),
.B(n_1518),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1558),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1558),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1567),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1567),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1575),
.B(n_1526),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1551),
.Y(n_1589)
);

CKINVDCx16_ASAP7_75t_R g1590 ( 
.A(n_1572),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1560),
.B(n_1528),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1553),
.A2(n_1525),
.B1(n_1538),
.B2(n_1529),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1560),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1575),
.B(n_1529),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1553),
.B(n_1515),
.Y(n_1595)
);

OAI21xp33_ASAP7_75t_L g1596 ( 
.A1(n_1592),
.A2(n_1595),
.B(n_1579),
.Y(n_1596)
);

AOI211xp5_ASAP7_75t_L g1597 ( 
.A1(n_1595),
.A2(n_1550),
.B(n_1563),
.C(n_1561),
.Y(n_1597)
);

OAI21xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1576),
.A2(n_1562),
.B(n_1574),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1592),
.B(n_1571),
.C(n_1570),
.Y(n_1599)
);

NAND4xp25_ASAP7_75t_L g1600 ( 
.A(n_1581),
.B(n_1570),
.C(n_1563),
.D(n_1554),
.Y(n_1600)
);

OAI21xp33_ASAP7_75t_L g1601 ( 
.A1(n_1576),
.A2(n_1562),
.B(n_1556),
.Y(n_1601)
);

AOI21xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1590),
.A2(n_1573),
.B(n_1568),
.Y(n_1602)
);

AOI211xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1582),
.A2(n_1564),
.B(n_1538),
.C(n_1566),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1583),
.B(n_1522),
.Y(n_1604)
);

AOI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1591),
.A2(n_1522),
.B1(n_1472),
.B2(n_1547),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1588),
.A2(n_1547),
.B(n_1545),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1593),
.A2(n_1522),
.B1(n_1514),
.B2(n_1539),
.Y(n_1607)
);

OAI211xp5_ASAP7_75t_L g1608 ( 
.A1(n_1598),
.A2(n_1578),
.B(n_1580),
.C(n_1593),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1604),
.Y(n_1609)
);

NOR3x1_ASAP7_75t_L g1610 ( 
.A(n_1600),
.B(n_1578),
.C(n_1594),
.Y(n_1610)
);

NOR3x1_ASAP7_75t_L g1611 ( 
.A(n_1599),
.B(n_1577),
.C(n_1589),
.Y(n_1611)
);

NAND4xp25_ASAP7_75t_L g1612 ( 
.A(n_1596),
.B(n_1587),
.C(n_1586),
.D(n_1585),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1606),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1601),
.B(n_1584),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1602),
.B(n_1522),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1605),
.Y(n_1616)
);

AO22x2_ASAP7_75t_L g1617 ( 
.A1(n_1597),
.A2(n_1539),
.B1(n_1514),
.B2(n_1482),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_SL g1618 ( 
.A(n_1603),
.B(n_1473),
.C(n_1471),
.Y(n_1618)
);

NOR2x1_ASAP7_75t_L g1619 ( 
.A(n_1607),
.B(n_1473),
.Y(n_1619)
);

AOI211xp5_ASAP7_75t_L g1620 ( 
.A1(n_1608),
.A2(n_1519),
.B(n_1320),
.C(n_1488),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1614),
.B(n_1519),
.Y(n_1621)
);

NOR3xp33_ASAP7_75t_L g1622 ( 
.A(n_1609),
.B(n_1318),
.C(n_1317),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1619),
.Y(n_1623)
);

NOR4xp25_ASAP7_75t_L g1624 ( 
.A(n_1612),
.B(n_1492),
.C(n_1484),
.D(n_1482),
.Y(n_1624)
);

NAND4xp25_ASAP7_75t_SL g1625 ( 
.A(n_1616),
.B(n_1492),
.C(n_1506),
.D(n_1503),
.Y(n_1625)
);

OAI211xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1613),
.A2(n_1615),
.B(n_1611),
.C(n_1610),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1623),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1624),
.B(n_1617),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1621),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1625),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1626),
.A2(n_1618),
.B1(n_1467),
.B2(n_1506),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1622),
.Y(n_1632)
);

NAND4xp75_ASAP7_75t_L g1633 ( 
.A(n_1630),
.B(n_1620),
.C(n_1455),
.D(n_1512),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1627),
.B(n_1464),
.Y(n_1634)
);

AOI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1628),
.A2(n_1512),
.B1(n_1467),
.B2(n_1470),
.C(n_1450),
.Y(n_1635)
);

NOR3xp33_ASAP7_75t_L g1636 ( 
.A(n_1629),
.B(n_1632),
.C(n_1628),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_L g1637 ( 
.A(n_1631),
.B(n_1470),
.C(n_1467),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1636),
.B(n_1464),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1634),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1633),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1638),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_L g1642 ( 
.A(n_1641),
.B(n_1640),
.C(n_1639),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1642),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1642),
.Y(n_1644)
);

NOR2xp67_ASAP7_75t_L g1645 ( 
.A(n_1643),
.B(n_1637),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1644),
.A2(n_1635),
.B(n_1469),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1645),
.A2(n_1439),
.B1(n_1440),
.B2(n_1449),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1646),
.B(n_1467),
.C(n_1440),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1648),
.Y(n_1649)
);

AOI322xp5_ASAP7_75t_L g1650 ( 
.A1(n_1649),
.A2(n_1647),
.A3(n_1450),
.B1(n_1464),
.B2(n_1469),
.C1(n_1439),
.C2(n_1449),
.Y(n_1650)
);

AOI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1440),
.B1(n_1449),
.B2(n_1469),
.C(n_1450),
.Y(n_1651)
);

AOI211xp5_ASAP7_75t_L g1652 ( 
.A1(n_1651),
.A2(n_1314),
.B(n_1310),
.C(n_1308),
.Y(n_1652)
);


endmodule