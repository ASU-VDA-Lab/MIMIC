module real_jpeg_10363_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_325, n_11, n_14, n_7, n_3, n_5, n_4, n_324, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_325;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_324;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_1),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_23),
.B1(n_60),
.B2(n_61),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_1),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_2),
.A2(n_11),
.B(n_32),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_3),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_140),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_140),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_140),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_6),
.A2(n_34),
.B1(n_60),
.B2(n_61),
.Y(n_218)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_45),
.B(n_58),
.C(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_9),
.B(n_45),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_10),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_53),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_11),
.A2(n_45),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_11),
.B(n_45),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_11),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_11),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_11),
.A2(n_31),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_11),
.B(n_31),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_11),
.B(n_35),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_106),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_12),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_93),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_93),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_14),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_55),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_15),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_15),
.A2(n_45),
.B1(n_46),
.B2(n_86),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_86),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_86),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_16),
.A2(n_60),
.B1(n_61),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_16),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_122),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_122),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_16),
.A2(n_24),
.B1(n_25),
.B2(n_122),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_17),
.A2(n_60),
.B1(n_61),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_17),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_81),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_81),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_17),
.A2(n_24),
.B1(n_25),
.B2(n_81),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_316),
.B(n_319),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_68),
.B(n_315),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_21),
.B(n_36),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_21),
.B(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_21),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_22),
.A2(n_26),
.B1(n_35),
.B2(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_24),
.A2(n_28),
.B(n_106),
.C(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_26),
.A2(n_35),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_26),
.A2(n_33),
.B(n_35),
.Y(n_318)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_27),
.A2(n_30),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_27),
.A2(n_30),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_27),
.A2(n_30),
.B1(n_203),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_27),
.A2(n_30),
.B1(n_228),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_27),
.A2(n_30),
.B1(n_246),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_27),
.A2(n_30),
.B1(n_52),
.B2(n_267),
.Y(n_289)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_42),
.Y(n_43)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_64),
.C(n_66),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_37),
.A2(n_38),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_50),
.C(n_56),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_39),
.A2(n_40),
.B1(n_56),
.B2(n_293),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_44),
.B(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_41),
.A2(n_44),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_41),
.A2(n_44),
.B1(n_131),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_41),
.A2(n_44),
.B1(n_148),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_41),
.A2(n_44),
.B1(n_188),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_41),
.A2(n_44),
.B1(n_199),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_41),
.A2(n_44),
.B1(n_225),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_41),
.A2(n_44),
.B1(n_243),
.B2(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_41),
.A2(n_44),
.B1(n_48),
.B2(n_260),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_44),
.B(n_106),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_45),
.B(n_47),
.Y(n_135)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_46),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_50),
.A2(n_51),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_56),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_56),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_59),
.B(n_63),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_59),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_57),
.A2(n_59),
.B1(n_92),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_57),
.A2(n_59),
.B1(n_119),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_57),
.A2(n_59),
.B1(n_127),
.B2(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_57),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_57),
.A2(n_59),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_57),
.A2(n_59),
.B1(n_211),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_57),
.A2(n_59),
.B1(n_220),
.B2(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_57),
.A2(n_59),
.B1(n_63),
.B2(n_252),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_59),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_59),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_60),
.B(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_60),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_61),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_64),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_308),
.B(n_314),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_285),
.A3(n_303),
.B1(n_306),
.B2(n_307),
.C(n_324),
.Y(n_69)
);

AOI321xp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_236),
.A3(n_273),
.B1(n_279),
.B2(n_284),
.C(n_325),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_193),
.C(n_232),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_163),
.B(n_192),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_142),
.B(n_162),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_124),
.B(n_141),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_113),
.B(n_123),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_99),
.B(n_112),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_82),
.A2(n_83),
.B1(n_139),
.B2(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_103),
.B1(n_104),
.B2(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_94),
.B2(n_98),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_98),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_107),
.B(n_111),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_104),
.B1(n_121),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_103),
.A2(n_104),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_103),
.A2(n_104),
.B1(n_174),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_103),
.A2(n_104),
.B1(n_208),
.B2(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_103),
.A2(n_104),
.B(n_218),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_115),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_125),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.CI(n_120),
.CON(n_116),
.SN(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_128),
.CI(n_132),
.CON(n_125),
.SN(n_125)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_143),
.B(n_144),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_155),
.B2(n_156),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_158),
.C(n_160),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_149),
.B1(n_150),
.B2(n_154),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_147),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_152),
.C(n_154),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_164),
.B(n_165),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_178),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_167),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_167),
.B(n_177),
.C(n_178),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_172),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_189),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_186),
.B2(n_187),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_186),
.C(n_189),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_194),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_213),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_195),
.B(n_213),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.C(n_212),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_205),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_204),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_198),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_SL g230 ( 
.A(n_200),
.B(n_204),
.C(n_205),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_212),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_209),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_230),
.B2(n_231),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_221),
.C(n_231),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_219),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_226),
.C(n_229),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_226),
.B1(n_227),
.B2(n_229),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_224),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_230),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_234),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_255),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_237),
.B(n_255),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_248),
.C(n_254),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_238),
.A2(n_239),
.B1(n_248),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_244),
.C(n_247),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_242),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_248),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_249),
.A2(n_250),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_249),
.A2(n_266),
.B(n_269),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_251),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_251),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_271),
.B2(n_272),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_263),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_263),
.C(n_272),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_261),
.B(n_262),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_261),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_287),
.C(n_295),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_262),
.B(n_287),
.CI(n_295),
.CON(n_305),
.SN(n_305)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_269),
.B2(n_270),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_271),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_280),
.B(n_283),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_296),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_296),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_289),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_293),
.C(n_294),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_298),
.C(n_302),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_305),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_313),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_310),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_321),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);


endmodule