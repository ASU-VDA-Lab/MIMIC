module fake_jpeg_27055_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_15),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_64),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_36),
.B1(n_22),
.B2(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_55),
.A2(n_59),
.B1(n_70),
.B2(n_17),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_36),
.B1(n_35),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_80),
.B1(n_19),
.B2(n_17),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_57),
.B(n_63),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_72),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_28),
.B1(n_33),
.B2(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_71),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_27),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_27),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_47),
.Y(n_94)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_21),
.B1(n_26),
.B2(n_31),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_38),
.A2(n_21),
.B1(n_26),
.B2(n_23),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_39),
.B1(n_37),
.B2(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_37),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_43),
.B(n_2),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_84),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_85),
.B(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_87),
.B(n_92),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_88),
.B(n_53),
.Y(n_154)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_90),
.Y(n_126)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_98),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_118),
.B1(n_19),
.B2(n_25),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_34),
.B(n_29),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_111),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_1),
.B(n_2),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_104),
.Y(n_131)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_106),
.Y(n_132)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_65),
.B1(n_38),
.B2(n_25),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_54),
.A2(n_41),
.B(n_40),
.C(n_39),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_110),
.A2(n_51),
.B1(n_73),
.B2(n_78),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_37),
.C(n_47),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_31),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_120),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_63),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_38),
.B1(n_54),
.B2(n_65),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_82),
.Y(n_142)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_51),
.A2(n_29),
.B1(n_41),
.B2(n_32),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_61),
.B(n_29),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_32),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_25),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_55),
.B(n_37),
.C(n_47),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_139),
.B1(n_148),
.B2(n_151),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_109),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_146),
.B1(n_113),
.B2(n_99),
.Y(n_159)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_140),
.Y(n_155)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_147),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_87),
.B1(n_103),
.B2(n_92),
.Y(n_148)
);

INVx5_ASAP7_75t_SL g149 ( 
.A(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_122),
.A2(n_46),
.B1(n_83),
.B2(n_71),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_94),
.A2(n_58),
.B1(n_32),
.B2(n_37),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_154),
.B1(n_53),
.B2(n_20),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_101),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_14),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_97),
.B(n_84),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_1),
.B(n_2),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_169),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_91),
.B(n_121),
.C(n_108),
.D(n_98),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_175),
.C(n_144),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_91),
.A3(n_113),
.B1(n_100),
.B2(n_114),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_14),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_111),
.B1(n_88),
.B2(n_100),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_106),
.B1(n_109),
.B2(n_85),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_170),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_172),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_176),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_95),
.B1(n_86),
.B2(n_90),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_86),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_149),
.A2(n_89),
.B1(n_58),
.B2(n_119),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_174),
.B1(n_179),
.B2(n_186),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_149),
.A2(n_119),
.B1(n_107),
.B2(n_112),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_95),
.C(n_53),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_93),
.C(n_116),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_102),
.C(n_47),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_183),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_2),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_102),
.B1(n_20),
.B2(n_39),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_124),
.B1(n_137),
.B2(n_154),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_148),
.A2(n_20),
.B1(n_8),
.B2(n_14),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_53),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_182),
.B(n_184),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_1),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_128),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_187),
.B(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g242 ( 
.A1(n_190),
.A2(n_202),
.B(n_7),
.Y(n_242)
);

INVxp33_ASAP7_75t_SL g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_124),
.B1(n_154),
.B2(n_145),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_162),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_137),
.B1(n_151),
.B2(n_143),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_138),
.B1(n_125),
.B2(n_140),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_197),
.A2(n_199),
.B(n_200),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_203),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_147),
.B(n_125),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_201),
.B(n_8),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_217),
.Y(n_225)
);

NAND2x1p5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_1),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_206),
.A2(n_212),
.B(n_214),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_13),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_215),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_211),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_13),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_216),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_3),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_4),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_156),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_242),
.B1(n_203),
.B2(n_196),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_176),
.C(n_170),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_232),
.C(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_173),
.B1(n_180),
.B2(n_172),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_230),
.B1(n_244),
.B2(n_196),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_233),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_184),
.B1(n_160),
.B2(n_177),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_182),
.C(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_175),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_238),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_192),
.C(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_243),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_190),
.A2(n_9),
.A3(n_12),
.B1(n_6),
.B2(n_7),
.C1(n_4),
.C2(n_5),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_200),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_192),
.B(n_9),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_4),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_251),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_249),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_216),
.B1(n_206),
.B2(n_212),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_250),
.B1(n_243),
.B2(n_231),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_194),
.B1(n_222),
.B2(n_220),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_209),
.B(n_214),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_259),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_209),
.B1(n_211),
.B2(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_262),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_214),
.B(n_218),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_217),
.B(n_5),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_244),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_222),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_6),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_6),
.C(n_235),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_224),
.C(n_232),
.Y(n_268)
);

XOR2x2_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_234),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_269),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_278),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_230),
.C(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_225),
.C(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_266),
.C(n_260),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

OAI211xp5_ASAP7_75t_SL g276 ( 
.A1(n_253),
.A2(n_225),
.B(n_236),
.C(n_228),
.Y(n_276)
);

OAI31xp33_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_256),
.A3(n_261),
.B(n_251),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_256),
.B(n_229),
.CI(n_233),
.CON(n_277),
.SN(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_281),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_259),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_250),
.B(n_263),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_286),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_267),
.A2(n_249),
.B1(n_254),
.B2(n_255),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_286),
.A2(n_280),
.B1(n_279),
.B2(n_276),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_295),
.C(n_296),
.Y(n_305)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_260),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_272),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_297),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_247),
.C(n_258),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_252),
.C(n_270),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_291),
.A2(n_274),
.B(n_283),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_301),
.A2(n_292),
.B(n_287),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_306),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_304),
.A2(n_303),
.B1(n_307),
.B2(n_306),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_279),
.B(n_280),
.C(n_296),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_295),
.B(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_292),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_312),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_306),
.B(n_305),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_305),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_320),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_315),
.B(n_321),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_306),
.B1(n_302),
.B2(n_293),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_322),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_309),
.Y(n_322)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_319),
.B(n_324),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_326),
.Y(n_329)
);


endmodule