module fake_jpeg_28412_n_197 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_197);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_25),
.Y(n_54)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_40),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_31),
.B1(n_32),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_56),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_31),
.B1(n_18),
.B2(n_32),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_41),
.B1(n_35),
.B2(n_42),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_21),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_32),
.B1(n_31),
.B2(n_18),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_37),
.B1(n_25),
.B2(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_64),
.B(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_72),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_17),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_70),
.Y(n_92)
);

NOR2x1_ASAP7_75t_R g96 ( 
.A(n_69),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_30),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_55),
.B1(n_53),
.B2(n_44),
.Y(n_105)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_19),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_22),
.B(n_20),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_29),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_20),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_84),
.B(n_29),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_96),
.B1(n_105),
.B2(n_65),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_91),
.Y(n_110)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_51),
.A3(n_19),
.B1(n_39),
.B2(n_26),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_67),
.B(n_76),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_60),
.B1(n_58),
.B2(n_51),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_46),
.B1(n_63),
.B2(n_39),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_26),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_75),
.B(n_72),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_58),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_67),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_104),
.B(n_64),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_63),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_73),
.B1(n_82),
.B2(n_67),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_124),
.B1(n_85),
.B2(n_101),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_116),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_87),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_67),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_123),
.C(n_95),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_65),
.B1(n_83),
.B2(n_46),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_120),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_89),
.B1(n_96),
.B2(n_93),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_53),
.C(n_44),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_129),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_135),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_100),
.B(n_98),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_137),
.B(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_114),
.B1(n_109),
.B2(n_120),
.C(n_108),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_100),
.B(n_92),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_92),
.B1(n_85),
.B2(n_94),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_140),
.B1(n_141),
.B2(n_27),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_94),
.B1(n_106),
.B2(n_27),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_145),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g145 ( 
.A(n_143),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_118),
.C(n_123),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_134),
.C(n_137),
.Y(n_159)
);

OAI211xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_158),
.B(n_142),
.C(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_129),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_122),
.B1(n_106),
.B2(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_135),
.Y(n_163)
);

AO221x1_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_166),
.C(n_150),
.Y(n_175)
);

NOR4xp25_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_167),
.C(n_156),
.D(n_10),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_157),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_150),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_142),
.C(n_136),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_139),
.A3(n_132),
.B1(n_140),
.B2(n_11),
.C1(n_14),
.C2(n_15),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_24),
.B1(n_12),
.B2(n_11),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_169),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_176),
.B1(n_168),
.B2(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_1),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_159),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_175),
.C(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_146),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

AOI321xp33_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_154),
.A3(n_153),
.B1(n_12),
.B2(n_4),
.C(n_5),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_2),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_153),
.B(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_4),
.C(n_6),
.Y(n_189)
);

OAI31xp33_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_154),
.A3(n_161),
.B(n_3),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_3),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_173),
.B1(n_175),
.B2(n_6),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_189),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_190),
.A2(n_191),
.B(n_193),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_181),
.B1(n_182),
.B2(n_8),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_8),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_192),
.A2(n_189),
.B(n_8),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_195),
.B(n_191),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_194),
.Y(n_197)
);


endmodule