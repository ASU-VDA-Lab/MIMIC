module fake_jpeg_29334_n_488 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_488);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_488;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_8),
.B(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_38),
.C(n_28),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_54),
.A2(n_22),
.B(n_49),
.Y(n_134)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_57),
.Y(n_159)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_58),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_35),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_59),
.B(n_22),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_72),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_27),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_75),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_16),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_84),
.Y(n_138)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_33),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_14),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_87),
.B(n_90),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_21),
.B(n_14),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_24),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_49),
.Y(n_137)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_116),
.B(n_100),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_22),
.B1(n_47),
.B2(n_26),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_45),
.B1(n_34),
.B2(n_31),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_45),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_39),
.Y(n_175)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_68),
.Y(n_141)
);

NAND2x1_ASAP7_75t_SL g212 ( 
.A(n_141),
.B(n_150),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_53),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_45),
.Y(n_183)
);

INVx6_ASAP7_75t_SL g150 ( 
.A(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_76),
.Y(n_156)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_160),
.Y(n_240)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_163),
.A2(n_26),
.B(n_47),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_51),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_169),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_102),
.A2(n_54),
.B(n_42),
.C(n_44),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_167),
.B(n_213),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_46),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_23),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_170),
.B(n_172),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_102),
.B(n_46),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_175),
.B(n_188),
.Y(n_255)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_178),
.Y(n_257)
);

OR2x4_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_47),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_179),
.A2(n_44),
.B(n_42),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_108),
.A2(n_86),
.B1(n_82),
.B2(n_67),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_197),
.B1(n_92),
.B2(n_118),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_101),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_181),
.B(n_201),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_183),
.B(n_184),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_105),
.B(n_39),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_190),
.Y(n_238)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_128),
.Y(n_187)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_105),
.B(n_72),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_114),
.A2(n_60),
.B1(n_64),
.B2(n_74),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_189),
.A2(n_57),
.B1(n_159),
.B2(n_91),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_23),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_138),
.B(n_21),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_196),
.Y(n_252)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_109),
.Y(n_194)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_117),
.B(n_44),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_125),
.A2(n_66),
.B1(n_56),
.B2(n_80),
.Y(n_197)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_136),
.B(n_31),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_207),
.Y(n_254)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_112),
.B(n_95),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_144),
.B(n_81),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_104),
.C(n_115),
.Y(n_245)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_110),
.Y(n_210)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_103),
.A2(n_89),
.B1(n_88),
.B2(n_85),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_211),
.A2(n_113),
.B1(n_145),
.B2(n_121),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_127),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_119),
.Y(n_214)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_SL g286 ( 
.A(n_219),
.B(n_246),
.C(n_70),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_220),
.B(n_245),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_115),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_226),
.B(n_248),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_164),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_235),
.A2(n_241),
.B1(n_208),
.B2(n_42),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_179),
.A2(n_124),
.B1(n_155),
.B2(n_120),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_249),
.B1(n_189),
.B2(n_194),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_183),
.B(n_135),
.C(n_26),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_167),
.B(n_157),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_180),
.A2(n_145),
.B1(n_132),
.B2(n_121),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_198),
.B1(n_159),
.B2(n_195),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_174),
.B(n_131),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_212),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_214),
.Y(n_277)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_263),
.A2(n_283),
.B1(n_240),
.B2(n_228),
.Y(n_316)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_264),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_265),
.B(n_275),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_182),
.B(n_192),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_266),
.A2(n_296),
.B(n_277),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_268),
.A2(n_269),
.B1(n_274),
.B2(n_278),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_220),
.A2(n_206),
.B1(n_129),
.B2(n_132),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_208),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_270),
.A2(n_286),
.B(n_257),
.Y(n_315)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_273),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_277),
.B(n_287),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_241),
.B1(n_229),
.B2(n_233),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_162),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_280),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_171),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_282),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_129),
.B1(n_79),
.B2(n_193),
.Y(n_283)
);

INVx13_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_290),
.Y(n_309)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_285),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_218),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_216),
.A2(n_178),
.B1(n_168),
.B2(n_206),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_288),
.A2(n_292),
.B1(n_297),
.B2(n_228),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_289),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_218),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_243),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_293),
.Y(n_308)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_227),
.B(n_252),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_294),
.B(n_295),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_165),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_244),
.A2(n_235),
.B(n_219),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_216),
.A2(n_160),
.B1(n_205),
.B2(n_210),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_299),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_221),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_248),
.A3(n_246),
.B1(n_231),
.B2(n_244),
.Y(n_300)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_226),
.B(n_244),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_301),
.A2(n_317),
.B(n_272),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_302),
.A2(n_321),
.B(n_272),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_274),
.A2(n_161),
.B1(n_203),
.B2(n_173),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_322),
.B1(n_287),
.B2(n_290),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_240),
.C(n_257),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_323),
.C(n_325),
.Y(n_337)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_261),
.A2(n_234),
.A3(n_222),
.B1(n_217),
.B2(n_256),
.Y(n_311)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_318),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_316),
.A2(n_319),
.B1(n_324),
.B2(n_292),
.Y(n_357)
);

A2O1A1O1Ixp25_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_234),
.B(n_34),
.C(n_31),
.D(n_237),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_271),
.A2(n_185),
.B1(n_239),
.B2(n_222),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_34),
.B(n_176),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_295),
.A2(n_120),
.B1(n_143),
.B2(n_199),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_266),
.B(n_70),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_263),
.A2(n_209),
.B1(n_199),
.B2(n_176),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_41),
.C(n_13),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_270),
.A2(n_41),
.B(n_2),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_327),
.A2(n_272),
.B(n_289),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_280),
.B(n_41),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_332),
.C(n_323),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_13),
.Y(n_332)
);

OA22x2_ASAP7_75t_L g366 ( 
.A1(n_338),
.A2(n_353),
.B1(n_316),
.B2(n_319),
.Y(n_366)
);

NOR3xp33_ASAP7_75t_SL g339 ( 
.A(n_305),
.B(n_279),
.C(n_267),
.Y(n_339)
);

NOR3xp33_ASAP7_75t_SL g386 ( 
.A(n_339),
.B(n_313),
.C(n_273),
.Y(n_386)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_333),
.Y(n_341)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_333),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_342),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_267),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_350),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_321),
.A2(n_270),
.B(n_294),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_310),
.A2(n_270),
.B1(n_298),
.B2(n_291),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_345),
.A2(n_324),
.B1(n_311),
.B2(n_304),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_308),
.B(n_270),
.Y(n_346)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_348),
.B(n_356),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_299),
.Y(n_349)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_349),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_303),
.B(n_284),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_351),
.B(n_365),
.Y(n_381)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_307),
.Y(n_352)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_352),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g353 ( 
.A(n_301),
.B(n_284),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_309),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_361),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_281),
.Y(n_355)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_315),
.A2(n_289),
.B(n_262),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_357),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_326),
.B(n_12),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_358),
.B(n_360),
.Y(n_383)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_307),
.Y(n_359)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_332),
.B(n_12),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_285),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_328),
.B(n_276),
.Y(n_362)
);

OAI21xp33_ASAP7_75t_L g377 ( 
.A1(n_362),
.A2(n_363),
.B(n_364),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_306),
.B(n_282),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_282),
.Y(n_364)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_378),
.B1(n_348),
.B2(n_356),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_330),
.Y(n_370)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_371),
.A2(n_374),
.B1(n_345),
.B2(n_349),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_363),
.B(n_300),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_335),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_340),
.A2(n_328),
.B1(n_329),
.B2(n_320),
.Y(n_374)
);

AOI322xp5_ASAP7_75t_SL g376 ( 
.A1(n_339),
.A2(n_318),
.A3(n_327),
.B1(n_276),
.B2(n_273),
.C1(n_264),
.C2(n_292),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_376),
.B(n_0),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_336),
.A2(n_325),
.B1(n_329),
.B2(n_313),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_312),
.Y(n_380)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_320),
.Y(n_384)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_336),
.B(n_364),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_385),
.B(n_386),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_331),
.C(n_334),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_337),
.C(n_365),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_350),
.Y(n_393)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_393),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_357),
.B1(n_362),
.B2(n_338),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_397),
.A2(n_398),
.B1(n_407),
.B2(n_411),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_399),
.A2(n_388),
.B1(n_366),
.B2(n_374),
.Y(n_426)
);

XNOR2x1_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_372),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_403),
.C(n_406),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_351),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_355),
.Y(n_404)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_346),
.C(n_335),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_367),
.A2(n_368),
.B1(n_378),
.B2(n_390),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_361),
.C(n_347),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_408),
.B(n_366),
.C(n_389),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_359),
.B1(n_352),
.B2(n_353),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_409),
.A2(n_415),
.B1(n_383),
.B2(n_391),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_368),
.A2(n_344),
.B(n_353),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_410),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_344),
.B1(n_334),
.B2(n_331),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_412),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_360),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_372),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_382),
.A2(n_12),
.B(n_2),
.Y(n_414)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_414),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_395),
.A2(n_375),
.B1(n_386),
.B2(n_382),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_417),
.A2(n_426),
.B1(n_395),
.B2(n_411),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_421),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_375),
.C(n_379),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_424),
.C(n_425),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_379),
.C(n_388),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_407),
.A2(n_366),
.B1(n_387),
.B2(n_391),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_414),
.B1(n_5),
.B2(n_6),
.Y(n_445)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_428),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_404),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_429),
.B(n_4),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_387),
.C(n_4),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_431),
.C(n_413),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_0),
.Y(n_431)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_432),
.Y(n_435)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_435),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_410),
.Y(n_437)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_437),
.Y(n_456)
);

AO22x1_ASAP7_75t_L g438 ( 
.A1(n_419),
.A2(n_412),
.B1(n_398),
.B2(n_399),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_438),
.A2(n_439),
.B1(n_422),
.B2(n_427),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_441),
.B(n_447),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_401),
.C(n_394),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_416),
.C(n_424),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_423),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_445),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_426),
.A2(n_400),
.B1(n_396),
.B2(n_405),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_444),
.A2(n_423),
.B1(n_433),
.B2(n_421),
.Y(n_455)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_434),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_448),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_422),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_445),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_455),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_436),
.A2(n_434),
.B1(n_418),
.B2(n_431),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_457),
.A2(n_459),
.B1(n_4),
.B2(n_6),
.Y(n_470)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_458),
.B(n_441),
.C(n_425),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_438),
.A2(n_444),
.B1(n_437),
.B2(n_443),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_437),
.A2(n_430),
.B(n_416),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_461),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_442),
.C(n_449),
.Y(n_461)
);

INVx11_ASAP7_75t_L g462 ( 
.A(n_453),
.Y(n_462)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_462),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_435),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_464),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_460),
.B(n_440),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_469),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_470),
.C(n_454),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_450),
.B(n_447),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_463),
.B(n_461),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_474),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_465),
.A2(n_459),
.B1(n_452),
.B2(n_455),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_475),
.A2(n_464),
.B1(n_456),
.B2(n_469),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_474),
.B(n_468),
.C(n_458),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_479),
.C(n_480),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_476),
.B(n_457),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_471),
.C(n_472),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_481),
.A2(n_478),
.B(n_9),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_483),
.A2(n_8),
.B(n_9),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_484),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_485),
.A2(n_8),
.B(n_10),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_486),
.B(n_482),
.Y(n_487)
);

OAI21xp33_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_10),
.B(n_11),
.Y(n_488)
);


endmodule