module fake_jpeg_6033_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_37),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_42),
.CON(n_54),
.SN(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_38),
.Y(n_73)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_44),
.Y(n_55)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_32),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_23),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_45),
.C(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_28),
.B1(n_21),
.B2(n_26),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_60),
.B1(n_62),
.B2(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_43),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_59),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_41),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_28),
.B1(n_21),
.B2(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_28),
.B1(n_21),
.B2(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_74),
.A2(n_64),
.B1(n_68),
.B2(n_19),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_36),
.B1(n_34),
.B2(n_39),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_73),
.B1(n_47),
.B2(n_19),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_36),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_96),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_30),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_21),
.B1(n_19),
.B2(n_39),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_43),
.B(n_38),
.C(n_31),
.Y(n_125)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_19),
.B1(n_39),
.B2(n_34),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_73),
.B1(n_34),
.B2(n_39),
.Y(n_115)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_101),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_110),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_49),
.C(n_62),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_126),
.C(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_116),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_114),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_122),
.B1(n_127),
.B2(n_64),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_124),
.B1(n_88),
.B2(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_72),
.C(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_86),
.B(n_18),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_136),
.B1(n_77),
.B2(n_88),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_143),
.C(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_140),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_150),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_76),
.C(n_85),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_85),
.B(n_76),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_105),
.B(n_114),
.Y(n_167)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_85),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

BUFx24_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_86),
.Y(n_154)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_79),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_170),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_120),
.B(n_101),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g198 ( 
.A(n_159),
.B(n_167),
.C(n_172),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_162),
.C(n_166),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_125),
.B(n_122),
.C(n_99),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_169),
.B1(n_178),
.B2(n_180),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_109),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_102),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_165),
.Y(n_188)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_125),
.C(n_121),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_124),
.C(n_123),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_99),
.B1(n_143),
.B2(n_131),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_99),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_113),
.B(n_116),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_130),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_139),
.C(n_138),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_119),
.B1(n_70),
.B2(n_68),
.Y(n_178)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_79),
.A3(n_64),
.B1(n_48),
.B2(n_95),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_35),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_83),
.B1(n_46),
.B2(n_38),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_155),
.B1(n_156),
.B2(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_94),
.B1(n_92),
.B2(n_77),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_185),
.B(n_192),
.Y(n_234)
);

AOI22x1_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_142),
.B1(n_135),
.B2(n_147),
.Y(n_187)
);

AOI22x1_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_94),
.B1(n_35),
.B2(n_63),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_196),
.C(n_197),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_202),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_153),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_148),
.C(n_84),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_18),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_18),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_153),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_132),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_205),
.B(n_175),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_23),
.B(n_30),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_132),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_178),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_211),
.B1(n_77),
.B2(n_30),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_161),
.B1(n_169),
.B2(n_159),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_212),
.A2(n_222),
.B1(n_225),
.B2(n_191),
.Y(n_251)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_161),
.B(n_164),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_217),
.B(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_181),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_218),
.B(n_201),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_173),
.B1(n_166),
.B2(n_161),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_226),
.B1(n_235),
.B2(n_204),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_232),
.Y(n_239)
);

OAI311xp33_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_22),
.A3(n_23),
.B1(n_153),
.C1(n_16),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_29),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_95),
.B(n_22),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_71),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_71),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_190),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_95),
.B1(n_17),
.B2(n_69),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_190),
.C(n_197),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_24),
.C(n_17),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_259),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_198),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_187),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_256),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_237),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_250),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_253),
.Y(n_264)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_205),
.B1(n_29),
.B2(n_16),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_227),
.B1(n_230),
.B2(n_214),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_260),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_71),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_59),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_258),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_24),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_220),
.B(n_24),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_265),
.Y(n_295)
);

XOR2x1_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_212),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_267),
.B(n_16),
.Y(n_292)
);

OAI322xp33_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_228),
.A3(n_213),
.B1(n_225),
.B2(n_235),
.C1(n_221),
.C2(n_24),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_279),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_238),
.A2(n_213),
.B1(n_17),
.B2(n_29),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_277),
.B1(n_11),
.B2(n_15),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_24),
.C(n_2),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_0),
.B(n_1),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_24),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_257),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_280),
.A2(n_292),
.B(n_270),
.C(n_265),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_274),
.A2(n_243),
.B1(n_239),
.B2(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_282),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_286),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_239),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_284),
.A2(n_290),
.B(n_261),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_242),
.C(n_10),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_291),
.C(n_293),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_271),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_273),
.B1(n_268),
.B2(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_272),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_17),
.B1(n_29),
.B2(n_16),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_281),
.B1(n_293),
.B2(n_292),
.Y(n_303)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_9),
.C(n_15),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_297),
.B(n_298),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_275),
.C(n_268),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_302),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_262),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_304),
.C(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_262),
.C(n_277),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_303),
.B(n_308),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_294),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_279),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_8),
.B1(n_12),
.B2(n_10),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_289),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_1),
.C(n_2),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_1),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_312),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_297),
.A2(n_304),
.B(n_306),
.Y(n_314)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_6),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_14),
.B1(n_10),
.B2(n_9),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_318),
.B1(n_3),
.B2(n_5),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_8),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_296),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_300),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_318)
);

AOI21xp33_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_3),
.B(n_5),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_299),
.C(n_305),
.Y(n_322)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_324),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_299),
.Y(n_324)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_3),
.B(n_5),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_327),
.A2(n_328),
.B(n_6),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_6),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_333),
.B(n_323),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_311),
.C(n_314),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

AO21x1_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_6),
.B(n_7),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_330),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_331),
.Y(n_339)
);


endmodule