module fake_netlist_5_1017_n_6007 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_649, n_552, n_547, n_43, n_721, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_725, n_139, n_38, n_105, n_280, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_302, n_265, n_526, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_692, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_724, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_138, n_264, n_109, n_669, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_727, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_691, n_717, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_700, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_722, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_726, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_720, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_713, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_256, n_305, n_533, n_52, n_278, n_110, n_6007);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_725;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_302;
input n_265;
input n_526;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_692;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_724;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_691;
input n_717;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_700;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_722;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_726;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_713;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_6007;

wire n_924;
wire n_977;
wire n_2253;
wire n_2756;
wire n_2417;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_5287;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_5978;
wire n_2395;
wire n_5161;
wire n_5776;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_877;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_1728;
wire n_2076;
wire n_1107;
wire n_5480;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_1242;
wire n_3283;
wire n_5469;
wire n_2323;
wire n_5744;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_5202;
wire n_5648;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_3214;
wire n_1517;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_5922;
wire n_1449;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_5848;
wire n_5406;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_882;
wire n_2384;
wire n_3156;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_5661;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_2276;
wire n_5852;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_845;
wire n_4255;
wire n_1796;
wire n_5577;
wire n_901;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_5689;
wire n_5894;
wire n_2079;
wire n_2238;
wire n_1151;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_5825;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_1000;
wire n_5686;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_748;
wire n_1667;
wire n_1058;
wire n_838;
wire n_3983;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_5909;
wire n_1385;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_5397;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_5709;
wire n_3208;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_5695;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_5860;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5862;
wire n_5189;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_1027;
wire n_4160;
wire n_2293;
wire n_5854;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_5936;
wire n_1199;
wire n_1038;
wire n_1841;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_1711;
wire n_870;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_965;
wire n_3790;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_5479;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_1194;
wire n_5888;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_5870;
wire n_1464;
wire n_4295;
wire n_5303;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_1121;
wire n_4391;
wire n_949;
wire n_5954;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_1195;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_757;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_1145;
wire n_5624;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_1153;
wire n_3856;
wire n_741;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_1207;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_940;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_978;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_5745;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4232;
wire n_4125;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_962;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_974;
wire n_5210;
wire n_4967;
wire n_5657;
wire n_957;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2729;
wire n_2261;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_4198;
wire n_2077;
wire n_2909;
wire n_5857;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_5756;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_5708;
wire n_3213;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_3474;
wire n_3984;
wire n_5927;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_4189;
wire n_5670;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_5965;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_948;
wire n_5751;
wire n_5664;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_5641;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_5963;
wire n_5980;
wire n_824;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_815;
wire n_4594;
wire n_3424;
wire n_5970;
wire n_1381;
wire n_1037;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_5690;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_5885;
wire n_2254;
wire n_1382;
wire n_925;
wire n_3546;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_950;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_968;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_5362;
wire n_4355;
wire n_3494;
wire n_5702;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_5527;
wire n_802;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_1305;
wire n_5266;
wire n_3178;
wire n_873;
wire n_5355;
wire n_2334;
wire n_4521;
wire n_4488;
wire n_5977;
wire n_2289;
wire n_3051;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_5551;
wire n_3715;
wire n_972;
wire n_5767;
wire n_3040;
wire n_1938;
wire n_5640;
wire n_1200;
wire n_2499;
wire n_3568;
wire n_5655;
wire n_5475;
wire n_3737;
wire n_1185;
wire n_991;
wire n_1967;
wire n_1329;
wire n_3255;
wire n_5692;
wire n_4856;
wire n_2997;
wire n_5921;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_883;
wire n_5322;
wire n_856;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_918;
wire n_4761;
wire n_942;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_5418;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_5933;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_763;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_4010;
wire n_1219;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_5644;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_789;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_4052;
wire n_5864;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_5460;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_5570;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_5983;
wire n_1661;
wire n_5804;
wire n_3565;
wire n_4701;
wire n_2575;
wire n_5910;
wire n_5040;
wire n_861;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_1899;
wire n_1003;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_1726;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_5717;
wire n_5464;
wire n_1657;
wire n_5886;
wire n_768;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3639;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_5610;
wire n_1109;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_2484;
wire n_808;
wire n_797;
wire n_5785;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_5994;
wire n_4538;
wire n_766;
wire n_1117;
wire n_2754;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3661;
wire n_3536;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_1137;
wire n_3934;
wire n_4985;
wire n_5788;
wire n_3922;
wire n_3846;
wire n_5897;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_5795;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_1890;
wire n_4220;
wire n_1944;
wire n_909;
wire n_5630;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_756;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_5775;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_760;
wire n_5731;
wire n_5581;
wire n_3691;
wire n_3628;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_5831;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_5884;
wire n_2447;
wire n_4764;
wire n_886;
wire n_5653;
wire n_1221;
wire n_5394;
wire n_2774;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_751;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_5889;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_5764;
wire n_5428;
wire n_3391;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_5543;
wire n_816;
wire n_5678;
wire n_5935;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_5950;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_5995;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_6006;
wire n_3245;
wire n_4417;
wire n_4899;
wire n_796;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1012;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_3509;
wire n_3352;
wire n_5671;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_1061;
wire n_3251;
wire n_2931;
wire n_5185;
wire n_1193;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_781;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_5945;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_5565;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_5780;
wire n_5643;
wire n_3238;
wire n_3210;
wire n_5846;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_805;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_3347;
wire n_1074;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_5401;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_1186;
wire n_5883;
wire n_5319;
wire n_1018;
wire n_2247;
wire n_1622;
wire n_1180;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5706;
wire n_5337;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_5364;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_5895;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_819;
wire n_5088;
wire n_2302;
wire n_5457;
wire n_951;
wire n_5532;
wire n_1494;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_933;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_5544;
wire n_3832;
wire n_3987;
wire n_902;
wire n_5987;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_5538;
wire n_5919;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_5410;
wire n_3332;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_3782;
wire n_2978;
wire n_4208;
wire n_2458;
wire n_2058;
wire n_3786;
wire n_2888;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_5503;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_5958;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_5654;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_5999;
wire n_4485;
wire n_4626;
wire n_1097;
wire n_1036;
wire n_798;
wire n_2659;
wire n_1414;
wire n_4975;
wire n_1852;
wire n_5602;
wire n_3089;
wire n_2470;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_1391;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_5903;
wire n_813;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_1064;
wire n_5842;
wire n_858;
wire n_2985;
wire n_5722;
wire n_5636;
wire n_5065;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_5667;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_5918;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_1211;
wire n_3367;
wire n_4464;
wire n_5877;
wire n_907;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_2356;
wire n_892;
wire n_4556;
wire n_5454;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_5913;
wire n_5621;
wire n_2919;
wire n_4327;
wire n_953;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_5573;
wire n_4353;
wire n_2042;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_5529;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_5800;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_847;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_822;
wire n_5645;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_5779;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_809;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_5697;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_747;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_851;
wire n_843;
wire n_3775;
wire n_4133;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_5882;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_5672;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_5693;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_5486;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_906;
wire n_919;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_5782;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_995;
wire n_1609;
wire n_5298;
wire n_5596;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_5728;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_5726;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_1043;
wire n_5095;
wire n_3002;
wire n_5324;
wire n_3897;
wire n_1159;
wire n_5928;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_5911;
wire n_2418;
wire n_5589;
wire n_5841;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_5712;
wire n_1420;
wire n_3330;
wire n_1132;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_5633;
wire n_2896;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_5583;
wire n_1349;
wire n_4460;
wire n_1031;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_834;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_874;
wire n_5652;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_993;
wire n_3154;
wire n_1551;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_970;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_3242;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_921;
wire n_5100;
wire n_1795;
wire n_5849;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_3524;
wire n_5616;
wire n_5034;
wire n_1708;
wire n_5988;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_5959;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_1252;
wire n_5754;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_5628;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_967;
wire n_2731;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_5981;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_5720;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_5325;
wire n_5696;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_5759;
wire n_4478;
wire n_5753;
wire n_2646;
wire n_5536;
wire n_1605;
wire n_5173;
wire n_1228;
wire n_3920;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_5027;
wire n_5647;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_5738;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_945;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_984;
wire n_1983;
wire n_5975;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1147;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_1201;
wire n_1114;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_1176;
wire n_5940;
wire n_1149;
wire n_1020;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_5555;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_5784;
wire n_5576;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_3898;
wire n_849;
wire n_1786;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_875;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_5578;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_1401;
wire n_969;
wire n_4113;
wire n_1019;
wire n_1998;
wire n_4686;
wire n_5530;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_5741;
wire n_5991;
wire n_3933;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_778;
wire n_4068;
wire n_1122;
wire n_4872;
wire n_6000;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_5792;
wire n_1187;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_1174;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_1737;
wire n_774;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_1059;
wire n_1133;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_5651;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_5819;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5998;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_5476;
wire n_2003;
wire n_5856;
wire n_1457;
wire n_5446;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_5944;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_872;
wire n_5684;
wire n_5861;
wire n_1297;
wire n_5976;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_5312;
wire n_985;
wire n_5850;
wire n_3425;
wire n_3217;
wire n_3404;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_1602;
wire n_1178;
wire n_5687;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1318;
wire n_780;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_5674;
wire n_3600;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_5682;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_898;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_5612;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_5898;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_941;
wire n_3862;
wire n_5214;
wire n_5487;
wire n_5563;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_5497;
wire n_4724;
wire n_5832;
wire n_1238;
wire n_1772;
wire n_752;
wire n_1476;
wire n_1108;
wire n_5526;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_862;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5593;
wire n_5021;
wire n_2772;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_5737;
wire n_786;
wire n_1142;
wire n_2579;
wire n_1770;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_5560;
wire n_1873;
wire n_3201;
wire n_1087;
wire n_5666;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_1247;
wire n_3050;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_5272;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_5361;
wire n_5683;
wire n_4171;
wire n_5847;
wire n_4045;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_5740;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_5729;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_844;
wire n_5905;
wire n_3497;
wire n_1601;
wire n_5409;
wire n_2940;
wire n_5688;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2505;
wire n_2427;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_5798;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_5415;
wire n_4676;
wire n_5770;
wire n_5892;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_5676;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_5769;
wire n_1130;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_5341;
wire n_5930;
wire n_5814;
wire n_4881;
wire n_5979;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_5622;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_5546;
wire n_927;
wire n_2689;
wire n_3259;
wire n_5482;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_904;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_5966;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_5431;
wire n_1508;
wire n_785;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_5908;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_5939;
wire n_3766;
wire n_1353;
wire n_800;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_5931;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_915;
wire n_864;
wire n_5420;
wire n_1264;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_5835;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1118;
wire n_1686;
wire n_5679;
wire n_947;
wire n_3710;
wire n_5938;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_5891;
wire n_1230;
wire n_4144;
wire n_5724;
wire n_5774;
wire n_2165;
wire n_929;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1257;
wire n_1182;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_5923;
wire n_5790;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_1483;
wire n_2983;
wire n_3810;
wire n_1289;
wire n_2715;
wire n_5598;
wire n_2085;
wire n_1669;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_1670;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_5677;
wire n_4168;
wire n_3446;
wire n_5997;
wire n_955;
wire n_5511;
wire n_5680;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_5533;
wire n_5838;
wire n_897;
wire n_5280;
wire n_1428;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_5206;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_1267;
wire n_1801;
wire n_5419;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_1473;
wire n_3755;
wire n_5803;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1556;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_736;
wire n_5097;
wire n_2750;
wire n_5730;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_5816;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_1248;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_5748;
wire n_2942;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_944;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_857;
wire n_5650;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_971;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_3481;
wire n_5481;
wire n_2808;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_5821;
wire n_4491;
wire n_2930;
wire n_5733;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_5871;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_5707;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_5836;
wire n_914;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_759;
wire n_5585;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_4082;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_1537;
wire n_5875;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_1647;
wire n_4685;
wire n_5968;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5812;
wire n_5515;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_1233;
wire n_5607;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_946;
wire n_1539;
wire n_5734;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_738;
wire n_1624;
wire n_4970;
wire n_3816;
wire n_1279;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_2960;
wire n_1090;
wire n_5438;
wire n_4627;
wire n_758;
wire n_2290;
wire n_2045;
wire n_3783;
wire n_3369;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_1049;
wire n_2145;
wire n_5725;
wire n_1639;
wire n_3030;
wire n_1068;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_5768;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_5685;
wire n_1923;
wire n_5773;
wire n_5138;
wire n_1017;
wire n_5374;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1828;
wire n_2320;
wire n_1045;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5485;
wire n_5766;
wire n_5216;
wire n_1009;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_5805;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_743;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_2595;
wire n_761;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_5554;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_5639;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_5417;
wire n_4614;
wire n_1265;
wire n_2681;
wire n_3103;
wire n_765;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1015;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_5488;
wire n_1101;
wire n_1106;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_5781;
wire n_1455;
wire n_767;
wire n_2490;
wire n_1407;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_5747;
wire n_5969;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_4802;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_5437;
wire n_5826;
wire n_3881;
wire n_2461;
wire n_4583;
wire n_2243;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_1630;
wire n_4891;
wire n_1023;
wire n_5603;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_5716;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_1056;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_5456;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_5727;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_1060;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_5833;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_1112;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_5967;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_5982;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2948;
wire n_2309;
wire n_5827;
wire n_1560;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_804;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_1504;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_3572;
wire n_992;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_842;
wire n_5434;
wire n_2082;
wire n_5941;
wire n_1643;
wire n_5879;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_5669;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_3078;
wire n_894;
wire n_3253;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4599;
wire n_5830;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_5760;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_5668;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_5765;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_5513;
wire n_4803;
wire n_5972;
wire n_4079;
wire n_4091;
wire n_1638;
wire n_5916;
wire n_5984;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_830;
wire n_5191;
wire n_3085;
wire n_5869;
wire n_5925;
wire n_1655;
wire n_749;
wire n_5359;
wire n_2574;
wire n_1134;
wire n_5293;
wire n_1358;
wire n_4316;
wire n_939;
wire n_3697;
wire n_1232;
wire n_734;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_5510;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_5200;
wire n_1653;
wire n_5659;
wire n_1506;
wire n_5618;
wire n_2867;
wire n_990;
wire n_1894;
wire n_975;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_5858;
wire n_5817;
wire n_3402;
wire n_5723;
wire n_5295;
wire n_4679;
wire n_4115;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_1970;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_3902;
wire n_4730;
wire n_937;
wire n_2779;
wire n_1584;
wire n_3654;
wire n_2164;
wire n_5996;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_5796;
wire n_895;
wire n_3358;
wire n_5791;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_732;
wire n_5906;
wire n_4743;
wire n_3805;
wire n_1067;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_5423;
wire n_799;
wire n_1213;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_869;
wire n_5736;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_5700;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_2363;
wire n_4072;
wire n_916;
wire n_5579;
wire n_1115;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_823;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_5642;
wire n_3553;
wire n_5880;
wire n_4746;
wire n_5713;
wire n_6005;
wire n_1683;
wire n_1530;
wire n_997;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_2996;
wire n_1268;
wire n_5793;
wire n_5591;
wire n_1320;
wire n_4050;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_5623;
wire n_1063;
wire n_5681;
wire n_4853;
wire n_981;
wire n_867;
wire n_2422;
wire n_2239;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_5732;
wire n_3852;
wire n_5178;
wire n_812;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_905;
wire n_5077;
wire n_782;
wire n_5872;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_5735;
wire n_1330;
wire n_3072;
wire n_3313;
wire n_3081;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_934;
wire n_5314;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_5953;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_5952;
wire n_4739;
wire n_5820;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_5718;
wire n_787;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_930;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_5777;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_5951;
wire n_2442;
wire n_928;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_5701;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_5797;
wire n_4839;
wire n_5222;
wire n_5743;
wire n_1028;
wire n_4016;
wire n_5772;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_5801;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_5971;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_5502;
wire n_2027;
wire n_5568;
wire n_2642;
wire n_2500;
wire n_1918;
wire n_5656;
wire n_863;
wire n_4831;
wire n_2513;
wire n_5974;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_5413;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_5752;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_1089;
wire n_5217;
wire n_1004;
wire n_5957;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5490;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_4580;
wire n_1263;
wire n_5912;
wire n_1126;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_5557;
wire n_5472;
wire n_2955;
wire n_4112;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_5396;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_956;
wire n_2134;
wire n_5960;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_1545;
wire n_2374;
wire n_5859;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_854;
wire n_1799;
wire n_2396;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_1705;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_1280;
wire n_3650;
wire n_5840;
wire n_2761;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_920;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_976;
wire n_1949;
wire n_1946;
wire n_2936;
wire n_5914;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_5542;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_5519;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_5586;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_5675;
wire n_926;
wire n_2180;
wire n_2249;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_5771;
wire n_1547;
wire n_777;
wire n_1755;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_2915;
wire n_1239;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_5844;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_4745;
wire n_2337;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_5344;
wire n_923;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_3986;
wire n_4376;
wire n_5705;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5574;
wire n_5126;
wire n_1039;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_1403;
wire n_5553;
wire n_4042;
wire n_4176;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_5368;
wire n_1202;
wire n_5626;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5876;
wire n_5114;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4472;
wire n_4462;
wire n_3433;
wire n_1072;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_5699;
wire n_2450;
wire n_3447;
wire n_5810;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_5366;
wire n_1162;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_931;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_5901;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_4553;
wire n_746;
wire n_784;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1244;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_5867;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_913;
wire n_3833;
wire n_5632;
wire n_865;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_5660;
wire n_4645;
wire n_1191;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_3128;
wire n_5426;
wire n_744;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_5778;
wire n_5625;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_3000;
wire n_5429;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_5818;
wire n_5646;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_3457;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_5719;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_1781;
wire n_2084;
wire n_3648;
wire n_5749;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_959;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_1079;
wire n_5489;
wire n_1593;
wire n_3767;
wire n_2873;
wire n_2540;
wire n_4589;
wire n_2299;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_742;
wire n_750;
wire n_5436;
wire n_5907;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_5569;
wire n_5439;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_5715;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_4818;
wire n_4514;
wire n_4800;
wire n_1366;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_3399;
wire n_2628;
wire n_1249;
wire n_5932;
wire n_1111;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_5828;
wire n_2831;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_5054;
wire n_5631;
wire n_2467;
wire n_1094;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_1209;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_5326;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_5809;
wire n_1897;
wire n_764;
wire n_1424;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_5915;
wire n_5452;
wire n_4754;
wire n_4554;
wire n_5595;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_5535;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_841;
wire n_1050;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_5761;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_5929;
wire n_3362;
wire n_1631;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_1179;
wire n_753;
wire n_1048;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_5868;
wire n_4034;
wire n_1688;
wire n_3327;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_5989;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_896;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_5520;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_5947;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_814;
wire n_2707;
wire n_5920;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_5808;
wire n_3342;
wire n_1062;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_1204;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_3780;
wire n_783;
wire n_1928;
wire n_5244;
wire n_5382;
wire n_1188;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_5384;
wire n_3608;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_2444;
wire n_5789;
wire n_1110;
wire n_3123;
wire n_5787;
wire n_5056;
wire n_1088;
wire n_5249;
wire n_3393;
wire n_866;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_5866;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_5899;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_5247;
wire n_5865;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_5924;
wire n_3182;
wire n_5822;
wire n_2564;
wire n_4947;
wire n_876;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_966;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_5658;
wire n_3408;
wire n_899;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_1514;
wire n_1771;
wire n_1005;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_1168;
wire n_5564;
wire n_2445;
wire n_1427;
wire n_1835;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_5539;
wire n_3308;
wire n_791;
wire n_1533;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_1480;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_810;
wire n_2965;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_2213;
wire n_1170;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_5703;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_5534;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_5904;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_5572;
wire n_5750;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_1762;
wire n_1013;
wire n_3023;
wire n_5881;
wire n_5815;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_5755;
wire n_825;
wire n_2819;
wire n_5949;
wire n_737;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_5955;
wire n_3959;
wire n_5763;
wire n_792;
wire n_3140;
wire n_5246;
wire n_5964;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_5665;
wire n_3069;
wire n_5498;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5783;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_6003;
wire n_5385;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_1129;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_961;
wire n_2250;
wire n_5845;
wire n_1225;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_5663;
wire n_994;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_5973;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_1223;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_5855;
wire n_2357;
wire n_1250;
wire n_5757;
wire n_3309;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_5704;
wire n_1086;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_5946;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_1113;
wire n_1277;
wire n_2591;
wire n_3384;
wire n_852;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5710;
wire n_5070;
wire n_1337;
wire n_4445;
wire n_5566;
wire n_5414;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_5834;
wire n_1076;
wire n_2823;
wire n_1408;
wire n_1761;
wire n_5874;
wire n_730;
wire n_5270;
wire n_5956;
wire n_795;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_5823;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_1583;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_5934;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_1032;
wire n_2614;
wire n_2991;
wire n_6001;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

INVx1_ASAP7_75t_L g729 ( 
.A(n_92),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_414),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_709),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_60),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_44),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_105),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_632),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_694),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_160),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_447),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_631),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_550),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_415),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_277),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_698),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_530),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_594),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_618),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_437),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_476),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_375),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_66),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_182),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_269),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_51),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_620),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_665),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_438),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_390),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_604),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_510),
.Y(n_759)
);

CKINVDCx16_ASAP7_75t_R g760 ( 
.A(n_120),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_430),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_687),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_128),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_299),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_658),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_13),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_123),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_160),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_439),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_579),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_170),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_408),
.Y(n_772)
);

BUFx5_ASAP7_75t_L g773 ( 
.A(n_333),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_710),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_130),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_163),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_29),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_661),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_609),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_208),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_38),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_477),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_177),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_307),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_706),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_711),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_104),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_727),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_277),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_465),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_62),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_592),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_288),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_52),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_130),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_664),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_565),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_439),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_116),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_339),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_708),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_716),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_122),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_385),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_51),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_189),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_65),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_389),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_140),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_492),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_616),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_721),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_451),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_728),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_113),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_695),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_691),
.Y(n_817)
);

BUFx10_ASAP7_75t_L g818 ( 
.A(n_265),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_241),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_689),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_204),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_10),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_553),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_336),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_724),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_247),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_669),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_571),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_314),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_177),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_200),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_81),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_650),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_183),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_126),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_21),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_638),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_315),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_700),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_20),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_393),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_335),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_122),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_567),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_349),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_684),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_363),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_85),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_333),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_95),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_726),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_639),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_581),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_618),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_43),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_164),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_517),
.Y(n_857)
);

BUFx10_ASAP7_75t_L g858 ( 
.A(n_693),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_450),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_113),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_560),
.Y(n_861)
);

BUFx10_ASAP7_75t_L g862 ( 
.A(n_157),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_167),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_454),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_166),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_622),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_702),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_74),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_199),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_202),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_677),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_718),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_252),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_510),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_565),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_555),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_435),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_266),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_211),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_221),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_322),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_346),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_237),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_262),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_600),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_260),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_697),
.Y(n_887)
);

BUFx10_ASAP7_75t_L g888 ( 
.A(n_722),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_191),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_85),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_410),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_430),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_100),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_553),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_598),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_523),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_380),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_221),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_3),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_582),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_56),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_252),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_269),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_194),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_585),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_480),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_251),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_63),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_511),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_292),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_144),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_427),
.Y(n_912)
);

BUFx10_ASAP7_75t_L g913 ( 
.A(n_467),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_242),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_123),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_83),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_635),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_666),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_76),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_345),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_336),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_529),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_38),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_380),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_571),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_44),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_169),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_560),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_110),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_176),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_117),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_655),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_292),
.Y(n_933)
);

CKINVDCx16_ASAP7_75t_R g934 ( 
.A(n_279),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_48),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_481),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_686),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_304),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_610),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_311),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_482),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_440),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_472),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_685),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_431),
.Y(n_945)
);

CKINVDCx14_ASAP7_75t_R g946 ( 
.A(n_186),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_138),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_282),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_134),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_60),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_184),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_634),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_714),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_549),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_356),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_57),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_272),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_337),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_279),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_212),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_265),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_1),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_37),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_328),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_585),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_192),
.Y(n_966)
);

BUFx10_ASAP7_75t_L g967 ( 
.A(n_362),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_331),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_159),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_257),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_348),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_157),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_314),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_297),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_56),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_391),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_654),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_688),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_488),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_354),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_341),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_548),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_327),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_90),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_472),
.Y(n_985)
);

INVxp67_ASAP7_75t_SL g986 ( 
.A(n_509),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_376),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_610),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_153),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_491),
.Y(n_990)
);

CKINVDCx14_ASAP7_75t_R g991 ( 
.A(n_646),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_337),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_449),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_386),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_165),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_219),
.Y(n_996)
);

BUFx10_ASAP7_75t_L g997 ( 
.A(n_66),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_247),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_701),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_696),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_550),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_154),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_37),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_163),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_578),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_450),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_465),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_116),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_705),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_533),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_21),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_91),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_63),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_30),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_612),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_725),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_660),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_647),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_699),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_609),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_147),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_115),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_395),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_300),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_605),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_601),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_161),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_231),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_97),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_538),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_690),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_9),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_246),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_554),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_505),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_227),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_383),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_681),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_428),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_601),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_395),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_334),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_651),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_88),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_347),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_76),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_625),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_386),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_469),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_501),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_451),
.Y(n_1051)
);

CKINVDCx16_ASAP7_75t_R g1052 ( 
.A(n_335),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_423),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_399),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_215),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_367),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_477),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_41),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_411),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_108),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_385),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_596),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_281),
.Y(n_1063)
);

CKINVDCx14_ASAP7_75t_R g1064 ( 
.A(n_40),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_167),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_283),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_1),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_354),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_355),
.Y(n_1069)
);

BUFx2_ASAP7_75t_SL g1070 ( 
.A(n_323),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_547),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_497),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_131),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_304),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_86),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_426),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_190),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_360),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_352),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_591),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_489),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_374),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_562),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_183),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_3),
.Y(n_1085)
);

BUFx10_ASAP7_75t_L g1086 ( 
.A(n_713),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_575),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_587),
.Y(n_1088)
);

BUFx2_ASAP7_75t_SL g1089 ( 
.A(n_633),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_442),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_411),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_303),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_494),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_662),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_18),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_70),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_415),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_274),
.Y(n_1098)
);

BUFx10_ASAP7_75t_L g1099 ( 
.A(n_641),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_595),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_549),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_351),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_667),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_577),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_364),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_617),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_227),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_45),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_452),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_438),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_84),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_90),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_458),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_234),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_501),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_707),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_201),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_583),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_715),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_717),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_374),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_282),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_239),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_148),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_219),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_615),
.Y(n_1126)
);

CKINVDCx14_ASAP7_75t_R g1127 ( 
.A(n_365),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_673),
.Y(n_1128)
);

BUFx5_ASAP7_75t_L g1129 ( 
.A(n_643),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_383),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_569),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_250),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_568),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_551),
.Y(n_1134)
);

BUFx10_ASAP7_75t_L g1135 ( 
.A(n_485),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_546),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_567),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_182),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_683),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_238),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_87),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_125),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_161),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_564),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_656),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_675),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_272),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_143),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_14),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_271),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_129),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_286),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_115),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_382),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_723),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_285),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_111),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_205),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_274),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_82),
.Y(n_1160)
);

INVx1_ASAP7_75t_SL g1161 ( 
.A(n_614),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_593),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_429),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_144),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_324),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_213),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_533),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_49),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_387),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_322),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_572),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_6),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_91),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_68),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_191),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_339),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_476),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_459),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_437),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_301),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_24),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_258),
.Y(n_1182)
);

CKINVDCx16_ASAP7_75t_R g1183 ( 
.A(n_166),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_370),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_49),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_202),
.Y(n_1186)
);

CKINVDCx16_ASAP7_75t_R g1187 ( 
.A(n_18),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_152),
.Y(n_1188)
);

BUFx5_ASAP7_75t_L g1189 ( 
.A(n_359),
.Y(n_1189)
);

CKINVDCx14_ASAP7_75t_R g1190 ( 
.A(n_271),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_425),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_513),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_626),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_107),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_16),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_165),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_266),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_82),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_543),
.Y(n_1199)
);

BUFx10_ASAP7_75t_L g1200 ( 
.A(n_350),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_602),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_78),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_537),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_179),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_569),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_463),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_692),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_526),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_146),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_614),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_131),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_200),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_599),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_413),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_270),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_253),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_111),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_293),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_416),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_720),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_147),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_71),
.Y(n_1222)
);

BUFx5_ASAP7_75t_L g1223 ( 
.A(n_620),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_59),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_27),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_173),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_379),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_181),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_140),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_676),
.Y(n_1230)
);

BUFx8_ASAP7_75t_SL g1231 ( 
.A(n_77),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_491),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_587),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_576),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_245),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_72),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_139),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_23),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_401),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_84),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_305),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_527),
.Y(n_1242)
);

CKINVDCx16_ASAP7_75t_R g1243 ( 
.A(n_74),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_514),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_86),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_535),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_246),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_103),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_268),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_475),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_158),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_305),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_204),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_703),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_590),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_712),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_427),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_313),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_559),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_150),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_207),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_589),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_308),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_611),
.Y(n_1264)
);

CKINVDCx16_ASAP7_75t_R g1265 ( 
.A(n_704),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_436),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_657),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_242),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_353),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_495),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_408),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_481),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_555),
.Y(n_1273)
);

INVxp67_ASAP7_75t_SL g1274 ( 
.A(n_401),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_293),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_98),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_529),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_14),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_356),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_180),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_719),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_129),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_53),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_473),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_43),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_311),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_578),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_485),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_773),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_773),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_773),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_814),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_773),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_773),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_829),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1231),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_773),
.Y(n_1297)
);

INVxp67_ASAP7_75t_SL g1298 ( 
.A(n_795),
.Y(n_1298)
);

INVxp33_ASAP7_75t_L g1299 ( 
.A(n_966),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_773),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_773),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_867),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1189),
.Y(n_1303)
);

INVxp67_ASAP7_75t_SL g1304 ( 
.A(n_795),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1189),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_871),
.Y(n_1306)
);

INVxp33_ASAP7_75t_L g1307 ( 
.A(n_1022),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1254),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_887),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1189),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_917),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_918),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1189),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_730),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_834),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1189),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1189),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1254),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1189),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_944),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1189),
.Y(n_1321)
);

INVxp33_ASAP7_75t_L g1322 ( 
.A(n_1126),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1223),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_946),
.B(n_0),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1223),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_952),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1223),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_863),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1223),
.Y(n_1329)
);

CKINVDCx20_ASAP7_75t_R g1330 ( 
.A(n_742),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1223),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1223),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_935),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1223),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1223),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_795),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1185),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1185),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_1185),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_767),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_767),
.Y(n_1341)
);

NOR2xp67_ASAP7_75t_L g1342 ( 
.A(n_1025),
.B(n_0),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_759),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_782),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_842),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_789),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_789),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_1114),
.B(n_2),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_953),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1064),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_916),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_916),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1075),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_842),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1075),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1116),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_760),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1079),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_828),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_842),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1079),
.Y(n_1361)
);

INVxp33_ASAP7_75t_L g1362 ( 
.A(n_1225),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1130),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_840),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_978),
.Y(n_1365)
);

INVxp33_ASAP7_75t_L g1366 ( 
.A(n_1105),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1130),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1136),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_842),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1136),
.Y(n_1370)
);

INVxp33_ASAP7_75t_SL g1371 ( 
.A(n_733),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1156),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1156),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_842),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1000),
.Y(n_1375)
);

BUFx8_ASAP7_75t_SL g1376 ( 
.A(n_1147),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_818),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1127),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1190),
.Y(n_1379)
);

INVxp33_ASAP7_75t_SL g1380 ( 
.A(n_733),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1160),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1160),
.Y(n_1382)
);

CKINVDCx16_ASAP7_75t_R g1383 ( 
.A(n_764),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_934),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_847),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_847),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_847),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1116),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_847),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_847),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_909),
.Y(n_1391)
);

INVxp33_ASAP7_75t_L g1392 ( 
.A(n_1272),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_909),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1230),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1017),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_909),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_909),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_909),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_818),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_920),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_920),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_920),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1018),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1254),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_920),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_818),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_920),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_857),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_968),
.Y(n_1409)
);

CKINVDCx14_ASAP7_75t_R g1410 ( 
.A(n_991),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_968),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_968),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_968),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_968),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_899),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_973),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_973),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_739),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_973),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_973),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_862),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_973),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_901),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_996),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1013),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1052),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_996),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1031),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_996),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_996),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_996),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1080),
.Y(n_1432)
);

INVxp67_ASAP7_75t_SL g1433 ( 
.A(n_1230),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1038),
.Y(n_1434)
);

CKINVDCx14_ASAP7_75t_R g1435 ( 
.A(n_858),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1080),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1080),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1043),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1080),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1080),
.Y(n_1440)
);

INVx4_ASAP7_75t_R g1441 ( 
.A(n_743),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1192),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1094),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1192),
.Y(n_1444)
);

INVxp33_ASAP7_75t_SL g1445 ( 
.A(n_739),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1192),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_740),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1192),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1192),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1229),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1229),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1229),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1229),
.Y(n_1453)
);

INVxp33_ASAP7_75t_SL g1454 ( 
.A(n_740),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1229),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_858),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1242),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1242),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_1183),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1242),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1242),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1242),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1103),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_731),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1129),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_963),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1187),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_729),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_732),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_734),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_737),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_738),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_746),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_747),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_985),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1119),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_748),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_753),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_758),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_772),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1243),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1129),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_741),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_866),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_775),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_776),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_780),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_741),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_783),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_790),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_791),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1003),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1015),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_794),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1072),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_868),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_798),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_803),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1083),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_805),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_807),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_821),
.Y(n_1502)
);

INVxp67_ASAP7_75t_SL g1503 ( 
.A(n_736),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_831),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_843),
.Y(n_1505)
);

INVxp33_ASAP7_75t_L g1506 ( 
.A(n_766),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_744),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_869),
.Y(n_1508)
);

CKINVDCx16_ASAP7_75t_R g1509 ( 
.A(n_1265),
.Y(n_1509)
);

INVxp67_ASAP7_75t_SL g1510 ( 
.A(n_762),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_853),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_854),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_858),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_855),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_856),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_859),
.Y(n_1516)
);

CKINVDCx16_ASAP7_75t_R g1517 ( 
.A(n_862),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_870),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1129),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_860),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_865),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1254),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_874),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_876),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_744),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_862),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_895),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_774),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_745),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_896),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_873),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_745),
.Y(n_1532)
);

INVxp33_ASAP7_75t_SL g1533 ( 
.A(n_749),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_788),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_908),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1087),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_911),
.Y(n_1537)
);

INVx1_ASAP7_75t_SL g1538 ( 
.A(n_1088),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_912),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_888),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_919),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_921),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_888),
.Y(n_1543)
);

INVxp33_ASAP7_75t_L g1544 ( 
.A(n_766),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_923),
.Y(n_1545)
);

INVxp67_ASAP7_75t_SL g1546 ( 
.A(n_802),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_926),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_929),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_875),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_936),
.Y(n_1550)
);

BUFx5_ASAP7_75t_L g1551 ( 
.A(n_812),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_942),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_943),
.Y(n_1553)
);

NOR2xp67_ASAP7_75t_L g1554 ( 
.A(n_1257),
.B(n_2),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_877),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1095),
.Y(n_1556)
);

CKINVDCx14_ASAP7_75t_R g1557 ( 
.A(n_888),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_804),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_948),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1129),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_957),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_959),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_878),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_960),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1129),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_965),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_913),
.Y(n_1567)
);

INVxp33_ASAP7_75t_SL g1568 ( 
.A(n_749),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1254),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_975),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_976),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_879),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_981),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_988),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_913),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_913),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_993),
.Y(n_1577)
);

INVxp67_ASAP7_75t_SL g1578 ( 
.A(n_816),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1096),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_995),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1001),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_750),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1006),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1007),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1014),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_817),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1020),
.Y(n_1587)
);

INVxp33_ASAP7_75t_SL g1588 ( 
.A(n_750),
.Y(n_1588)
);

INVxp33_ASAP7_75t_SL g1589 ( 
.A(n_751),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1129),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_947),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_880),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1021),
.Y(n_1593)
);

BUFx10_ASAP7_75t_L g1594 ( 
.A(n_743),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_882),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1033),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1047),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1048),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1060),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1115),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1138),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1073),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1085),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1093),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1097),
.Y(n_1605)
);

CKINVDCx16_ASAP7_75t_R g1606 ( 
.A(n_947),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1101),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_820),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1102),
.Y(n_1609)
);

INVxp33_ASAP7_75t_L g1610 ( 
.A(n_804),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1151),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1106),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_883),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_947),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_967),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1108),
.Y(n_1616)
);

INVxp67_ASAP7_75t_SL g1617 ( 
.A(n_837),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1110),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1112),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1129),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_884),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1134),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1165),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1154),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1166),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1171),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1180),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1196),
.Y(n_1628)
);

INVxp33_ASAP7_75t_L g1629 ( 
.A(n_810),
.Y(n_1629)
);

CKINVDCx16_ASAP7_75t_R g1630 ( 
.A(n_967),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1197),
.Y(n_1631)
);

INVxp33_ASAP7_75t_SL g1632 ( 
.A(n_751),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1198),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1129),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1199),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1206),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1209),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_810),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_885),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_886),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1210),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1212),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_890),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_822),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1213),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_891),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1215),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1216),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1232),
.Y(n_1649)
);

CKINVDCx16_ASAP7_75t_R g1650 ( 
.A(n_967),
.Y(n_1650)
);

CKINVDCx20_ASAP7_75t_R g1651 ( 
.A(n_1173),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_822),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1233),
.Y(n_1653)
);

CKINVDCx20_ASAP7_75t_R g1654 ( 
.A(n_1177),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1182),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1234),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_892),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_893),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1246),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_832),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1248),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1249),
.Y(n_1662)
);

BUFx5_ASAP7_75t_L g1663 ( 
.A(n_839),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_752),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1250),
.Y(n_1665)
);

INVx1_ASAP7_75t_SL g1666 ( 
.A(n_1191),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1253),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1258),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1262),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1259),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_997),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1260),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_752),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1275),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_754),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1277),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_846),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1278),
.Y(n_1678)
);

INVxp33_ASAP7_75t_L g1679 ( 
.A(n_832),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1283),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_852),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_872),
.Y(n_1682)
);

BUFx5_ASAP7_75t_L g1683 ( 
.A(n_932),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_937),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_894),
.Y(n_1685)
);

CKINVDCx20_ASAP7_75t_R g1686 ( 
.A(n_1271),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_977),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_999),
.Y(n_1688)
);

CKINVDCx14_ASAP7_75t_R g1689 ( 
.A(n_1086),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1009),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_897),
.Y(n_1691)
);

BUFx5_ASAP7_75t_L g1692 ( 
.A(n_1019),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1120),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1128),
.Y(n_1694)
);

NOR2xp67_ASAP7_75t_L g1695 ( 
.A(n_813),
.B(n_4),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_835),
.Y(n_1696)
);

CKINVDCx16_ASAP7_75t_R g1697 ( 
.A(n_997),
.Y(n_1697)
);

CKINVDCx16_ASAP7_75t_R g1698 ( 
.A(n_997),
.Y(n_1698)
);

INVxp33_ASAP7_75t_SL g1699 ( 
.A(n_754),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1146),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1220),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_835),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1281),
.Y(n_1703)
);

INVxp33_ASAP7_75t_L g1704 ( 
.A(n_864),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_827),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_827),
.Y(n_1706)
);

CKINVDCx16_ASAP7_75t_R g1707 ( 
.A(n_1032),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1139),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_864),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_889),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1139),
.Y(n_1711)
);

INVxp33_ASAP7_75t_SL g1712 ( 
.A(n_756),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1207),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1207),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_889),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_907),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_907),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_979),
.Y(n_1718)
);

INVxp33_ASAP7_75t_L g1719 ( 
.A(n_979),
.Y(n_1719)
);

INVxp33_ASAP7_75t_SL g1720 ( 
.A(n_756),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_980),
.Y(n_1721)
);

INVx4_ASAP7_75t_R g1722 ( 
.A(n_755),
.Y(n_1722)
);

INVxp33_ASAP7_75t_L g1723 ( 
.A(n_980),
.Y(n_1723)
);

NOR2xp67_ASAP7_75t_L g1724 ( 
.A(n_813),
.B(n_4),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1279),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1024),
.Y(n_1726)
);

INVxp33_ASAP7_75t_L g1727 ( 
.A(n_1024),
.Y(n_1727)
);

CKINVDCx16_ASAP7_75t_R g1728 ( 
.A(n_1032),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1030),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1030),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1076),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1032),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_755),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1076),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1078),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1078),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1090),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1090),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1098),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1086),
.Y(n_1740)
);

CKINVDCx5p33_ASAP7_75t_R g1741 ( 
.A(n_898),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1098),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_757),
.Y(n_1743)
);

INVxp33_ASAP7_75t_L g1744 ( 
.A(n_1113),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1113),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1181),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1181),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1186),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1357),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1385),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1324),
.B(n_1292),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1308),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1345),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1388),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1388),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1308),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1456),
.B(n_786),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1410),
.B(n_1086),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1298),
.B(n_786),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1481),
.Y(n_1760)
);

BUFx6f_ASAP7_75t_L g1761 ( 
.A(n_1308),
.Y(n_1761)
);

INVx4_ASAP7_75t_SL g1762 ( 
.A(n_1308),
.Y(n_1762)
);

OAI22x1_ASAP7_75t_SL g1763 ( 
.A1(n_1314),
.A2(n_757),
.B1(n_763),
.B2(n_761),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1318),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1410),
.B(n_1099),
.Y(n_1765)
);

BUFx8_ASAP7_75t_L g1766 ( 
.A(n_1315),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1318),
.Y(n_1767)
);

BUFx12f_ASAP7_75t_L g1768 ( 
.A(n_1296),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1325),
.A2(n_1331),
.B(n_1290),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1304),
.B(n_735),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1318),
.Y(n_1771)
);

BUFx12f_ASAP7_75t_L g1772 ( 
.A(n_1384),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1345),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1386),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1425),
.Y(n_1775)
);

BUFx12f_ASAP7_75t_L g1776 ( 
.A(n_1384),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1354),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1354),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1318),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1404),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_L g1781 ( 
.A(n_1404),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1387),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1302),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1389),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1390),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1484),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1404),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1391),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1306),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1393),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1522),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1366),
.A2(n_881),
.B1(n_933),
.B2(n_793),
.Y(n_1792)
);

INVx5_ASAP7_75t_L g1793 ( 
.A(n_1522),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1522),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1456),
.B(n_833),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1339),
.B(n_1464),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1503),
.B(n_735),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1371),
.A2(n_1082),
.B1(n_1274),
.B2(n_986),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1435),
.B(n_1557),
.Y(n_1799)
);

OAI22x1_ASAP7_75t_SL g1800 ( 
.A1(n_1314),
.A2(n_763),
.B1(n_768),
.B2(n_761),
.Y(n_1800)
);

BUFx12f_ASAP7_75t_L g1801 ( 
.A(n_1350),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1360),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1360),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1569),
.Y(n_1804)
);

OAI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1325),
.A2(n_1224),
.B(n_1186),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1396),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1369),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1510),
.B(n_1528),
.Y(n_1808)
);

CKINVDCx6p67_ASAP7_75t_R g1809 ( 
.A(n_1383),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1496),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1369),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1534),
.B(n_765),
.Y(n_1812)
);

INVxp67_ASAP7_75t_L g1813 ( 
.A(n_1488),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1546),
.B(n_1578),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1513),
.B(n_941),
.Y(n_1815)
);

CKINVDCx20_ASAP7_75t_R g1816 ( 
.A(n_1330),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1586),
.B(n_765),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1397),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1569),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1398),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1569),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1400),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1569),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1435),
.B(n_1099),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1374),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1374),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1449),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1449),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1426),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1733),
.Y(n_1830)
);

BUFx8_ASAP7_75t_SL g1831 ( 
.A(n_1376),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1558),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1309),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1401),
.Y(n_1834)
);

BUFx8_ASAP7_75t_SL g1835 ( 
.A(n_1376),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1733),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1608),
.B(n_778),
.Y(n_1837)
);

OA21x2_ASAP7_75t_L g1838 ( 
.A1(n_1289),
.A2(n_1252),
.B(n_1224),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1402),
.Y(n_1839)
);

BUFx12f_ASAP7_75t_L g1840 ( 
.A(n_1350),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1508),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1733),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1733),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1557),
.B(n_1099),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1405),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_L g1846 ( 
.A(n_1407),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1409),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1411),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1412),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1689),
.B(n_1135),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1558),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1413),
.Y(n_1852)
);

INVx5_ASAP7_75t_L g1853 ( 
.A(n_1594),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1414),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1416),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1467),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1417),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1617),
.B(n_778),
.Y(n_1858)
);

CKINVDCx6p67_ASAP7_75t_R g1859 ( 
.A(n_1459),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1371),
.A2(n_902),
.B1(n_903),
.B2(n_900),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1419),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1513),
.B(n_1540),
.Y(n_1862)
);

OA21x2_ASAP7_75t_L g1863 ( 
.A1(n_1291),
.A2(n_1252),
.B(n_1045),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1525),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1677),
.B(n_1688),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1420),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1529),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1681),
.B(n_1267),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1422),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1424),
.Y(n_1870)
);

BUFx12f_ASAP7_75t_L g1871 ( 
.A(n_1378),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1427),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1429),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1430),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1594),
.B(n_941),
.Y(n_1875)
);

OAI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1331),
.A2(n_1089),
.B(n_796),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1431),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1432),
.Y(n_1878)
);

INVx5_ASAP7_75t_L g1879 ( 
.A(n_1594),
.Y(n_1879)
);

OAI22x1_ASAP7_75t_SL g1880 ( 
.A1(n_1330),
.A2(n_769),
.B1(n_770),
.B2(n_768),
.Y(n_1880)
);

BUFx8_ASAP7_75t_L g1881 ( 
.A(n_1418),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1380),
.B(n_1045),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1311),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1682),
.B(n_785),
.Y(n_1884)
);

BUFx12f_ASAP7_75t_L g1885 ( 
.A(n_1378),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1436),
.Y(n_1886)
);

INVx4_ASAP7_75t_L g1887 ( 
.A(n_1312),
.Y(n_1887)
);

BUFx3_ASAP7_75t_L g1888 ( 
.A(n_1340),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1320),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1437),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1326),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1684),
.B(n_785),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1532),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1638),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1439),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1440),
.Y(n_1896)
);

BUFx12f_ASAP7_75t_L g1897 ( 
.A(n_1379),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1582),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1442),
.Y(n_1899)
);

INVx5_ASAP7_75t_L g1900 ( 
.A(n_1638),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1444),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1664),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1446),
.Y(n_1903)
);

OAI22x1_ASAP7_75t_L g1904 ( 
.A1(n_1406),
.A2(n_770),
.B1(n_771),
.B2(n_769),
.Y(n_1904)
);

BUFx6f_ASAP7_75t_L g1905 ( 
.A(n_1448),
.Y(n_1905)
);

BUFx12f_ASAP7_75t_L g1906 ( 
.A(n_1379),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1644),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1450),
.Y(n_1908)
);

INVx4_ASAP7_75t_L g1909 ( 
.A(n_1349),
.Y(n_1909)
);

CKINVDCx5p33_ASAP7_75t_R g1910 ( 
.A(n_1365),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1689),
.B(n_1135),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1451),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1452),
.Y(n_1913)
);

BUFx6f_ASAP7_75t_L g1914 ( 
.A(n_1453),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1455),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1457),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1380),
.B(n_1055),
.Y(n_1917)
);

BUFx8_ASAP7_75t_SL g1918 ( 
.A(n_1343),
.Y(n_1918)
);

AND2x2_ASAP7_75t_SL g1919 ( 
.A(n_1509),
.B(n_1070),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1445),
.A2(n_905),
.B1(n_906),
.B2(n_904),
.Y(n_1920)
);

INVx5_ASAP7_75t_L g1921 ( 
.A(n_1644),
.Y(n_1921)
);

AOI22x1_ASAP7_75t_SL g1922 ( 
.A1(n_1343),
.A2(n_777),
.B1(n_779),
.B2(n_771),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1458),
.Y(n_1923)
);

INVx5_ASAP7_75t_L g1924 ( 
.A(n_1652),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1460),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1461),
.Y(n_1926)
);

INVx2_ASAP7_75t_SL g1927 ( 
.A(n_1518),
.Y(n_1927)
);

AOI22x1_ASAP7_75t_SL g1928 ( 
.A1(n_1344),
.A2(n_779),
.B1(n_781),
.B2(n_777),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1462),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1687),
.B(n_1690),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1652),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1540),
.B(n_1055),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1336),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_L g1934 ( 
.A(n_1660),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1543),
.B(n_938),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1660),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1293),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1294),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1297),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1337),
.Y(n_1940)
);

BUFx8_ASAP7_75t_SL g1941 ( 
.A(n_1344),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1693),
.B(n_1267),
.Y(n_1942)
);

INVx4_ASAP7_75t_L g1943 ( 
.A(n_1375),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1300),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_1696),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1395),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1543),
.B(n_1141),
.Y(n_1947)
);

INVx4_ASAP7_75t_L g1948 ( 
.A(n_1403),
.Y(n_1948)
);

OA21x2_ASAP7_75t_L g1949 ( 
.A1(n_1301),
.A2(n_1305),
.B(n_1303),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1696),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1673),
.Y(n_1951)
);

INVx2_ASAP7_75t_SL g1952 ( 
.A(n_1531),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1356),
.B(n_1135),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1702),
.Y(n_1954)
);

INVx6_ASAP7_75t_L g1955 ( 
.A(n_1740),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1310),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1338),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_SL g1958 ( 
.A(n_1517),
.B(n_1200),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1341),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1740),
.B(n_1141),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1694),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1702),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1709),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1709),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1710),
.Y(n_1965)
);

BUFx12f_ASAP7_75t_L g1966 ( 
.A(n_1549),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1313),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1710),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1316),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1555),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1317),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1700),
.Y(n_1972)
);

BUFx8_ASAP7_75t_SL g1973 ( 
.A(n_1359),
.Y(n_1973)
);

OA21x2_ASAP7_75t_L g1974 ( 
.A1(n_1319),
.A2(n_914),
.B(n_910),
.Y(n_1974)
);

INVx3_ASAP7_75t_L g1975 ( 
.A(n_1468),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1394),
.B(n_1200),
.Y(n_1976)
);

CKINVDCx20_ASAP7_75t_R g1977 ( 
.A(n_1359),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1321),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1323),
.Y(n_1979)
);

INVx6_ASAP7_75t_L g1980 ( 
.A(n_1551),
.Y(n_1980)
);

INVx5_ASAP7_75t_L g1981 ( 
.A(n_1465),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1327),
.Y(n_1982)
);

INVx5_ASAP7_75t_L g1983 ( 
.A(n_1465),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1329),
.Y(n_1984)
);

INVx4_ASAP7_75t_L g1985 ( 
.A(n_1428),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1332),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1701),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1334),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1703),
.Y(n_1989)
);

OAI22x1_ASAP7_75t_L g1990 ( 
.A1(n_1421),
.A2(n_784),
.B1(n_787),
.B2(n_781),
.Y(n_1990)
);

HB1xp67_ASAP7_75t_L g1991 ( 
.A(n_1675),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1335),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1743),
.Y(n_1993)
);

INVx4_ASAP7_75t_L g1994 ( 
.A(n_1434),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1469),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1715),
.Y(n_1996)
);

INVx4_ASAP7_75t_L g1997 ( 
.A(n_1438),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1433),
.B(n_796),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1716),
.Y(n_1999)
);

BUFx12f_ASAP7_75t_L g2000 ( 
.A(n_1563),
.Y(n_2000)
);

OA21x2_ASAP7_75t_L g2001 ( 
.A1(n_1705),
.A2(n_922),
.B(n_915),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1717),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1447),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1470),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1471),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1551),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_1377),
.B(n_801),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1592),
.Y(n_2008)
);

BUFx12f_ASAP7_75t_L g2009 ( 
.A(n_1595),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1399),
.B(n_1295),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1483),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1507),
.Y(n_2012)
);

BUFx3_ASAP7_75t_L g2013 ( 
.A(n_1346),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1328),
.B(n_801),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1706),
.B(n_825),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1445),
.A2(n_925),
.B1(n_927),
.B2(n_924),
.Y(n_2016)
);

BUFx6f_ASAP7_75t_L g2017 ( 
.A(n_1718),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1443),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1551),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1708),
.B(n_825),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1721),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1613),
.B(n_1200),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1726),
.Y(n_2023)
);

AND2x6_ASAP7_75t_L g2024 ( 
.A(n_1482),
.B(n_940),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1472),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1621),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1711),
.B(n_1713),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1551),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1473),
.Y(n_2029)
);

INVx5_ASAP7_75t_L g2030 ( 
.A(n_1482),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1474),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1551),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1366),
.A2(n_1142),
.B1(n_1161),
.B2(n_1061),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_1463),
.Y(n_2034)
);

BUFx8_ASAP7_75t_SL g2035 ( 
.A(n_1364),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_1695),
.Y(n_2036)
);

INVx5_ASAP7_75t_L g2037 ( 
.A(n_1519),
.Y(n_2037)
);

CKINVDCx20_ASAP7_75t_R g2038 ( 
.A(n_1364),
.Y(n_2038)
);

INVx4_ASAP7_75t_L g2039 ( 
.A(n_1476),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1551),
.Y(n_2040)
);

AOI22xp5_ASAP7_75t_SL g2041 ( 
.A1(n_1392),
.A2(n_787),
.B1(n_792),
.B2(n_784),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1663),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1663),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1729),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1663),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1333),
.B(n_851),
.Y(n_2046)
);

BUFx3_ASAP7_75t_L g2047 ( 
.A(n_1347),
.Y(n_2047)
);

CKINVDCx16_ASAP7_75t_R g2048 ( 
.A(n_1575),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1730),
.Y(n_2049)
);

BUFx3_ASAP7_75t_L g2050 ( 
.A(n_1351),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1352),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1714),
.B(n_851),
.Y(n_2052)
);

BUFx8_ASAP7_75t_L g2053 ( 
.A(n_1353),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1663),
.Y(n_2054)
);

BUFx3_ASAP7_75t_L g2055 ( 
.A(n_1355),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_1639),
.Y(n_2056)
);

NOR2xp33_ASAP7_75t_L g2057 ( 
.A(n_1454),
.B(n_1016),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_1731),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1392),
.A2(n_1164),
.B1(n_1288),
.B2(n_1069),
.Y(n_2059)
);

AND2x4_ASAP7_75t_L g2060 ( 
.A(n_1358),
.B(n_1016),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1454),
.B(n_1145),
.Y(n_2061)
);

BUFx8_ASAP7_75t_SL g2062 ( 
.A(n_1408),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1361),
.B(n_1145),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1477),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1478),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1363),
.B(n_1155),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1663),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1663),
.B(n_1155),
.Y(n_2068)
);

BUFx6f_ASAP7_75t_L g2069 ( 
.A(n_1734),
.Y(n_2069)
);

BUFx12f_ASAP7_75t_L g2070 ( 
.A(n_1640),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1683),
.B(n_1256),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1683),
.B(n_1256),
.Y(n_2072)
);

BUFx12f_ASAP7_75t_L g2073 ( 
.A(n_1643),
.Y(n_2073)
);

OA21x2_ASAP7_75t_L g2074 ( 
.A1(n_1519),
.A2(n_930),
.B(n_928),
.Y(n_2074)
);

BUFx12f_ASAP7_75t_L g2075 ( 
.A(n_1646),
.Y(n_2075)
);

BUFx12f_ASAP7_75t_L g2076 ( 
.A(n_1657),
.Y(n_2076)
);

BUFx6f_ASAP7_75t_L g2077 ( 
.A(n_1735),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1479),
.Y(n_2078)
);

BUFx12f_ASAP7_75t_L g2079 ( 
.A(n_1658),
.Y(n_2079)
);

BUFx12f_ASAP7_75t_L g2080 ( 
.A(n_1685),
.Y(n_2080)
);

BUFx8_ASAP7_75t_SL g2081 ( 
.A(n_1408),
.Y(n_2081)
);

INVx4_ASAP7_75t_L g2082 ( 
.A(n_1691),
.Y(n_2082)
);

BUFx8_ASAP7_75t_SL g2083 ( 
.A(n_1415),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1683),
.Y(n_2084)
);

BUFx6f_ASAP7_75t_L g2085 ( 
.A(n_1736),
.Y(n_2085)
);

BUFx2_ASAP7_75t_L g2086 ( 
.A(n_1741),
.Y(n_2086)
);

OAI22x1_ASAP7_75t_R g2087 ( 
.A1(n_1415),
.A2(n_797),
.B1(n_799),
.B2(n_792),
.Y(n_2087)
);

BUFx3_ASAP7_75t_L g2088 ( 
.A(n_1367),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1737),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_1572),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1480),
.Y(n_2091)
);

OAI22x1_ASAP7_75t_L g2092 ( 
.A1(n_1526),
.A2(n_799),
.B1(n_800),
.B2(n_797),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1738),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1724),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1368),
.Y(n_2095)
);

AND2x4_ASAP7_75t_L g2096 ( 
.A(n_1370),
.B(n_931),
.Y(n_2096)
);

BUFx3_ASAP7_75t_L g2097 ( 
.A(n_1372),
.Y(n_2097)
);

BUFx8_ASAP7_75t_SL g2098 ( 
.A(n_1423),
.Y(n_2098)
);

BUFx8_ASAP7_75t_L g2099 ( 
.A(n_1373),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1683),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1683),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1485),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1683),
.B(n_939),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1692),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1692),
.Y(n_2105)
);

INVx3_ASAP7_75t_L g2106 ( 
.A(n_1486),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1487),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1692),
.B(n_945),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1489),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1560),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1490),
.Y(n_2111)
);

INVx4_ASAP7_75t_L g2112 ( 
.A(n_1572),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1491),
.Y(n_2113)
);

BUFx6f_ASAP7_75t_L g2114 ( 
.A(n_1739),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1560),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_1494),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1565),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1811),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1811),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1751),
.B(n_1692),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1995),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1828),
.Y(n_2122)
);

INVx4_ASAP7_75t_L g2123 ( 
.A(n_1981),
.Y(n_2123)
);

BUFx8_ASAP7_75t_L g2124 ( 
.A(n_1801),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1751),
.B(n_1692),
.Y(n_2125)
);

OAI21x1_ASAP7_75t_L g2126 ( 
.A1(n_1876),
.A2(n_1590),
.B(n_1565),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2004),
.Y(n_2127)
);

INVx3_ASAP7_75t_L g2128 ( 
.A(n_1752),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2103),
.B(n_1630),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1828),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1754),
.B(n_1497),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2005),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2025),
.Y(n_2133)
);

NOR2x1_ASAP7_75t_L g2134 ( 
.A(n_2082),
.B(n_1381),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2068),
.B(n_1692),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2029),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1753),
.Y(n_2137)
);

BUFx6f_ASAP7_75t_L g2138 ( 
.A(n_1752),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2064),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2065),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1773),
.Y(n_2141)
);

INVx4_ASAP7_75t_L g2142 ( 
.A(n_1981),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1777),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1752),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2078),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_1796),
.B(n_1533),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2091),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2102),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2107),
.Y(n_2149)
);

BUFx8_ASAP7_75t_L g2150 ( 
.A(n_1840),
.Y(n_2150)
);

BUFx3_ASAP7_75t_L g2151 ( 
.A(n_1754),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1752),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_1756),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2109),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1799),
.B(n_1506),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2036),
.B(n_1506),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2068),
.B(n_1590),
.Y(n_2157)
);

BUFx2_ASAP7_75t_L g2158 ( 
.A(n_1766),
.Y(n_2158)
);

AND2x2_ASAP7_75t_SL g2159 ( 
.A(n_1919),
.B(n_1606),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2111),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2113),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1961),
.Y(n_2162)
);

INVx6_ASAP7_75t_L g2163 ( 
.A(n_1955),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1972),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2036),
.B(n_1544),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2094),
.B(n_1544),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1987),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1989),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1967),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1967),
.Y(n_2170)
);

BUFx2_ASAP7_75t_L g2171 ( 
.A(n_1766),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2071),
.B(n_1620),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2071),
.B(n_1620),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1778),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1978),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2072),
.B(n_1634),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1756),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1756),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1802),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1803),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_1749),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2094),
.B(n_1610),
.Y(n_2182)
);

NOR2x1_ASAP7_75t_L g2183 ( 
.A(n_2082),
.B(n_1382),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1756),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_2103),
.B(n_1650),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2072),
.B(n_1634),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2108),
.B(n_1610),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_1796),
.B(n_1533),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_1761),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_SL g2190 ( 
.A(n_1958),
.B(n_1568),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1807),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2108),
.B(n_1629),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1825),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_1850),
.B(n_1629),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1978),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1978),
.Y(n_2196)
);

CKINVDCx11_ASAP7_75t_R g2197 ( 
.A(n_1816),
.Y(n_2197)
);

INVx3_ASAP7_75t_L g2198 ( 
.A(n_1761),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1761),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1978),
.Y(n_2200)
);

AND2x6_ASAP7_75t_L g2201 ( 
.A(n_1824),
.B(n_1498),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_1761),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1826),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1984),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1755),
.B(n_1500),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_1764),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1984),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_1755),
.B(n_1501),
.Y(n_2208)
);

AND2x2_ASAP7_75t_SL g2209 ( 
.A(n_1919),
.B(n_1697),
.Y(n_2209)
);

HB1xp67_ASAP7_75t_L g2210 ( 
.A(n_1749),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1984),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1847),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1814),
.B(n_1679),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1847),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_1764),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1886),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1814),
.B(n_1679),
.Y(n_2217)
);

BUFx3_ASAP7_75t_L g2218 ( 
.A(n_1955),
.Y(n_2218)
);

AOI22xp5_ASAP7_75t_L g2219 ( 
.A1(n_2057),
.A2(n_1568),
.B1(n_1589),
.B2(n_1588),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_1911),
.B(n_1844),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1984),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2024),
.B(n_1704),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_1888),
.B(n_1502),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1888),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1886),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1764),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1890),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1959),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2024),
.B(n_1808),
.Y(n_2229)
);

BUFx6f_ASAP7_75t_L g2230 ( 
.A(n_1764),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1890),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1795),
.B(n_1698),
.Y(n_2232)
);

INVxp67_ASAP7_75t_L g2233 ( 
.A(n_2057),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2024),
.B(n_1808),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1959),
.Y(n_2235)
);

INVx3_ASAP7_75t_L g2236 ( 
.A(n_1767),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2013),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_1853),
.B(n_1704),
.Y(n_2238)
);

BUFx6f_ASAP7_75t_L g2239 ( 
.A(n_1767),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2013),
.Y(n_2240)
);

OA21x2_ASAP7_75t_L g2241 ( 
.A1(n_1805),
.A2(n_1745),
.B(n_1742),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_1918),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1767),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1769),
.Y(n_2244)
);

INVx2_ASAP7_75t_SL g2245 ( 
.A(n_1998),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2047),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1767),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1931),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1931),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1931),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_1795),
.B(n_1707),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_1931),
.Y(n_2252)
);

BUFx6f_ASAP7_75t_L g2253 ( 
.A(n_1771),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2047),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2050),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2024),
.B(n_1719),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2050),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1853),
.B(n_1719),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2051),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2024),
.B(n_1723),
.Y(n_2260)
);

INVx3_ASAP7_75t_L g2261 ( 
.A(n_1771),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2051),
.Y(n_2262)
);

INVx4_ASAP7_75t_L g2263 ( 
.A(n_1981),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2055),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2055),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2088),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_1775),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2088),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1853),
.B(n_1879),
.Y(n_2269)
);

NAND2xp33_ASAP7_75t_L g2270 ( 
.A(n_1759),
.B(n_949),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_1955),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2095),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2095),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1853),
.B(n_1723),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2097),
.Y(n_2275)
);

BUFx6f_ASAP7_75t_L g2276 ( 
.A(n_1771),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2097),
.Y(n_2277)
);

BUFx2_ASAP7_75t_L g2278 ( 
.A(n_1775),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1937),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_1879),
.B(n_1727),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_1879),
.B(n_2010),
.Y(n_2281)
);

BUFx8_ASAP7_75t_L g2282 ( 
.A(n_1871),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_1798),
.A2(n_1589),
.B1(n_1632),
.B2(n_1588),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1938),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1939),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1944),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1956),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_1933),
.B(n_1504),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_1771),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1934),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1934),
.Y(n_2291)
);

BUFx6f_ASAP7_75t_L g2292 ( 
.A(n_1780),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1969),
.Y(n_2293)
);

BUFx2_ASAP7_75t_L g2294 ( 
.A(n_1829),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1934),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1934),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1971),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_1998),
.B(n_1728),
.Y(n_2298)
);

BUFx6f_ASAP7_75t_L g2299 ( 
.A(n_1780),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_1865),
.B(n_1632),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1979),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1936),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1982),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_1918),
.Y(n_2304)
);

NAND2xp33_ASAP7_75t_R g2305 ( 
.A(n_1974),
.B(n_2001),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1936),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_1780),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1986),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_L g2309 ( 
.A(n_1780),
.Y(n_2309)
);

BUFx8_ASAP7_75t_L g2310 ( 
.A(n_1885),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1988),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1992),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_1879),
.B(n_1727),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1936),
.Y(n_2314)
);

INVx3_ASAP7_75t_L g2315 ( 
.A(n_1781),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_1865),
.B(n_1770),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_1829),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1940),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1936),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1757),
.B(n_1759),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1957),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1945),
.Y(n_2322)
);

INVx3_ASAP7_75t_L g2323 ( 
.A(n_1781),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1830),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2010),
.B(n_1953),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1830),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_1945),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_1856),
.Y(n_2328)
);

AND2x4_ASAP7_75t_L g2329 ( 
.A(n_1975),
.B(n_1505),
.Y(n_2329)
);

AND2x6_ASAP7_75t_L g2330 ( 
.A(n_1758),
.B(n_1511),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1830),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1830),
.Y(n_2332)
);

INVx5_ASAP7_75t_L g2333 ( 
.A(n_1980),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1836),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1757),
.B(n_1744),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1836),
.Y(n_2336)
);

HB1xp67_ASAP7_75t_L g2337 ( 
.A(n_1856),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1836),
.Y(n_2338)
);

AND2x4_ASAP7_75t_L g2339 ( 
.A(n_1975),
.B(n_1512),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_1945),
.Y(n_2340)
);

INVx3_ASAP7_75t_L g2341 ( 
.A(n_1781),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1836),
.Y(n_2342)
);

XOR2xp5_ASAP7_75t_L g2343 ( 
.A(n_1816),
.B(n_1977),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_1976),
.B(n_1744),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2031),
.B(n_1514),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_2031),
.B(n_1515),
.Y(n_2346)
);

NOR2x1_ASAP7_75t_L g2347 ( 
.A(n_2112),
.B(n_1516),
.Y(n_2347)
);

OA21x2_ASAP7_75t_L g2348 ( 
.A1(n_1750),
.A2(n_1747),
.B(n_1746),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2106),
.B(n_1520),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1842),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_1781),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_1791),
.Y(n_2352)
);

HB1xp67_ASAP7_75t_L g2353 ( 
.A(n_2003),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2106),
.B(n_1521),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1945),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1842),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_1950),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_1950),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1842),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1770),
.B(n_1748),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1842),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1843),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1843),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1843),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_1813),
.B(n_1299),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1843),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1950),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1774),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_1791),
.Y(n_2369)
);

INVx5_ASAP7_75t_L g2370 ( 
.A(n_1980),
.Y(n_2370)
);

OAI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_1882),
.A2(n_1917),
.B1(n_1920),
.B2(n_1860),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_1797),
.B(n_1699),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_1782),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1784),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_1797),
.B(n_1699),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1785),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1950),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1788),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_1954),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_1790),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1806),
.Y(n_2381)
);

HB1xp67_ASAP7_75t_L g2382 ( 
.A(n_2003),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_1954),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1818),
.Y(n_2384)
);

BUFx6f_ASAP7_75t_L g2385 ( 
.A(n_1791),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1954),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1954),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1820),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_1813),
.B(n_1299),
.Y(n_2389)
);

INVx3_ASAP7_75t_L g2390 ( 
.A(n_1791),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_1794),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1822),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1834),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_1963),
.Y(n_2394)
);

BUFx6f_ASAP7_75t_L g2395 ( 
.A(n_1794),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1839),
.Y(n_2396)
);

BUFx8_ASAP7_75t_L g2397 ( 
.A(n_1897),
.Y(n_2397)
);

BUFx6f_ASAP7_75t_L g2398 ( 
.A(n_1794),
.Y(n_2398)
);

AND2x4_ASAP7_75t_L g2399 ( 
.A(n_2116),
.B(n_1523),
.Y(n_2399)
);

INVx5_ASAP7_75t_L g2400 ( 
.A(n_1980),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_1849),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_1812),
.B(n_1712),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_1864),
.B(n_1307),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_1864),
.B(n_1307),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_1963),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_1852),
.Y(n_2406)
);

AND2x6_ASAP7_75t_L g2407 ( 
.A(n_1765),
.B(n_1524),
.Y(n_2407)
);

BUFx3_ASAP7_75t_L g2408 ( 
.A(n_1838),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_1812),
.B(n_1712),
.Y(n_2409)
);

HB1xp67_ASAP7_75t_L g2410 ( 
.A(n_2011),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1855),
.Y(n_2411)
);

BUFx6f_ASAP7_75t_L g2412 ( 
.A(n_1794),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_1867),
.B(n_1322),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1861),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_1867),
.B(n_1322),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1866),
.Y(n_2416)
);

BUFx6f_ASAP7_75t_L g2417 ( 
.A(n_1804),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1963),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_1817),
.B(n_1720),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1869),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_1963),
.Y(n_2421)
);

OA21x2_ASAP7_75t_L g2422 ( 
.A1(n_1870),
.A2(n_1530),
.B(n_1527),
.Y(n_2422)
);

INVx3_ASAP7_75t_L g2423 ( 
.A(n_1804),
.Y(n_2423)
);

BUFx6f_ASAP7_75t_L g2424 ( 
.A(n_1804),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_1964),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_1817),
.B(n_1720),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_1804),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_1872),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1873),
.Y(n_2429)
);

HB1xp67_ASAP7_75t_L g2430 ( 
.A(n_2011),
.Y(n_2430)
);

INVxp33_ASAP7_75t_SL g2431 ( 
.A(n_2041),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1874),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1878),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1964),
.Y(n_2434)
);

AND2x4_ASAP7_75t_L g2435 ( 
.A(n_2116),
.B(n_1535),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_1964),
.Y(n_2436)
);

OAI22xp5_ASAP7_75t_SL g2437 ( 
.A1(n_1977),
.A2(n_1466),
.B1(n_1475),
.B2(n_1423),
.Y(n_2437)
);

BUFx2_ASAP7_75t_L g2438 ( 
.A(n_2038),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_1819),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1896),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_1981),
.Y(n_2441)
);

BUFx6f_ASAP7_75t_L g2442 ( 
.A(n_1819),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_1898),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_1964),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_1837),
.B(n_1537),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_1965),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_1837),
.B(n_1539),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_1965),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_1819),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1899),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_1965),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_1901),
.Y(n_2452)
);

AND2x6_ASAP7_75t_L g2453 ( 
.A(n_1815),
.B(n_1541),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_1908),
.Y(n_2454)
);

BUFx3_ASAP7_75t_L g2455 ( 
.A(n_1838),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_1858),
.B(n_1362),
.Y(n_2456)
);

BUFx3_ASAP7_75t_L g2457 ( 
.A(n_1838),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_1893),
.B(n_1362),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1913),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_1858),
.B(n_1542),
.Y(n_2460)
);

NAND2xp33_ASAP7_75t_L g2461 ( 
.A(n_1868),
.B(n_950),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_1926),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_1819),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_1823),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_1965),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1845),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_1893),
.B(n_1567),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2110),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_1902),
.B(n_1576),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2110),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_1823),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_1779),
.B(n_1545),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_1823),
.Y(n_2473)
);

HB1xp67_ASAP7_75t_L g2474 ( 
.A(n_1898),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_1845),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2115),
.Y(n_2476)
);

INVx1_ASAP7_75t_SL g2477 ( 
.A(n_1941),
.Y(n_2477)
);

INVx2_ASAP7_75t_SL g2478 ( 
.A(n_1815),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_1779),
.B(n_1547),
.Y(n_2479)
);

OA21x2_ASAP7_75t_L g2480 ( 
.A1(n_2015),
.A2(n_1550),
.B(n_1548),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_1845),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_1845),
.Y(n_2482)
);

INVx3_ASAP7_75t_L g2483 ( 
.A(n_1823),
.Y(n_2483)
);

CKINVDCx6p67_ASAP7_75t_R g2484 ( 
.A(n_1809),
.Y(n_2484)
);

CKINVDCx20_ASAP7_75t_R g2485 ( 
.A(n_2038),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_1787),
.B(n_1552),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2115),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_1846),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_1846),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_1902),
.B(n_1591),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_1862),
.B(n_1614),
.Y(n_2491)
);

BUFx6f_ASAP7_75t_L g2492 ( 
.A(n_1827),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2117),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_1827),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_1787),
.B(n_1553),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2117),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_1846),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_1827),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_SL g2499 ( 
.A(n_2056),
.B(n_1538),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_1821),
.B(n_1949),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_1846),
.Y(n_2501)
);

BUFx2_ASAP7_75t_L g2502 ( 
.A(n_1862),
.Y(n_2502)
);

INVx3_ASAP7_75t_L g2503 ( 
.A(n_1827),
.Y(n_2503)
);

INVxp67_ASAP7_75t_L g2504 ( 
.A(n_2061),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_1854),
.Y(n_2505)
);

BUFx6f_ASAP7_75t_L g2506 ( 
.A(n_1854),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_1848),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_1854),
.Y(n_2508)
);

INVx4_ASAP7_75t_L g2509 ( 
.A(n_1983),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_1857),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_1854),
.Y(n_2511)
);

HB1xp67_ASAP7_75t_L g2512 ( 
.A(n_1951),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_2007),
.B(n_1342),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_1877),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2007),
.B(n_1348),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_1905),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_1905),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_1905),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_1932),
.B(n_1615),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_1932),
.B(n_1671),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_1905),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_1821),
.B(n_1559),
.Y(n_2522)
);

HB1xp67_ASAP7_75t_L g2523 ( 
.A(n_1951),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_1947),
.B(n_1732),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_L g2525 ( 
.A(n_1914),
.Y(n_2525)
);

AOI22xp5_ASAP7_75t_L g2526 ( 
.A1(n_2061),
.A2(n_1554),
.B1(n_1669),
.B2(n_1666),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_1947),
.B(n_951),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_1914),
.Y(n_2528)
);

BUFx3_ASAP7_75t_L g2529 ( 
.A(n_1863),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_1949),
.B(n_1561),
.Y(n_2530)
);

HB1xp67_ASAP7_75t_L g2531 ( 
.A(n_1991),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_1895),
.Y(n_2532)
);

INVx3_ASAP7_75t_L g2533 ( 
.A(n_1983),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_1914),
.Y(n_2534)
);

BUFx6f_ASAP7_75t_L g2535 ( 
.A(n_1914),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_1915),
.Y(n_2536)
);

AND2x4_ASAP7_75t_L g2537 ( 
.A(n_1960),
.B(n_1562),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_1915),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_1960),
.B(n_1678),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_1915),
.Y(n_2540)
);

OAI21x1_ASAP7_75t_L g2541 ( 
.A1(n_1949),
.A2(n_1680),
.B(n_1566),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_1941),
.Y(n_2542)
);

INVx3_ASAP7_75t_L g2543 ( 
.A(n_1915),
.Y(n_2543)
);

AND2x6_ASAP7_75t_L g2544 ( 
.A(n_2006),
.B(n_1564),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1923),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_1903),
.Y(n_2546)
);

INVxp33_ASAP7_75t_L g2547 ( 
.A(n_2365),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2156),
.B(n_2022),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2244),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2244),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2241),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2241),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2121),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2241),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2348),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_2197),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2127),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2132),
.Y(n_2558)
);

INVx3_ASAP7_75t_L g2559 ( 
.A(n_2348),
.Y(n_2559)
);

NAND3xp33_ASAP7_75t_L g2560 ( 
.A(n_2300),
.B(n_1917),
.C(n_1882),
.Y(n_2560)
);

AOI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2375),
.A2(n_1974),
.B1(n_2001),
.B2(n_2074),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2468),
.Y(n_2562)
);

BUFx6f_ASAP7_75t_L g2563 ( 
.A(n_2408),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2133),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2468),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2136),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_2197),
.Y(n_2567)
);

BUFx3_ASAP7_75t_L g2568 ( 
.A(n_2151),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2470),
.Y(n_2569)
);

CKINVDCx11_ASAP7_75t_R g2570 ( 
.A(n_2484),
.Y(n_2570)
);

AO22x2_ASAP7_75t_L g2571 ( 
.A1(n_2371),
.A2(n_2233),
.B1(n_2504),
.B2(n_2234),
.Y(n_2571)
);

BUFx2_ASAP7_75t_L g2572 ( 
.A(n_2278),
.Y(n_2572)
);

BUFx2_ASAP7_75t_L g2573 ( 
.A(n_2294),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2165),
.B(n_1786),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2470),
.Y(n_2575)
);

AOI22xp33_ASAP7_75t_L g2576 ( 
.A1(n_2316),
.A2(n_1974),
.B1(n_1863),
.B2(n_2001),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2316),
.B(n_2074),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2139),
.Y(n_2578)
);

BUFx10_ASAP7_75t_L g2579 ( 
.A(n_2242),
.Y(n_2579)
);

NAND3xp33_ASAP7_75t_L g2580 ( 
.A(n_2300),
.B(n_2016),
.C(n_2012),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2140),
.Y(n_2581)
);

OAI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2229),
.A2(n_2012),
.B1(n_1952),
.B2(n_1927),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2145),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2372),
.B(n_2402),
.Y(n_2584)
);

AOI22xp33_ASAP7_75t_L g2585 ( 
.A1(n_2530),
.A2(n_1863),
.B1(n_2074),
.B2(n_2033),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2147),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2187),
.B(n_1887),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2148),
.Y(n_2588)
);

BUFx6f_ASAP7_75t_L g2589 ( 
.A(n_2408),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_SL g2590 ( 
.A(n_2409),
.B(n_2112),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2166),
.B(n_1810),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2348),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_2491),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2419),
.B(n_1783),
.Y(n_2594)
);

OR2x2_ASAP7_75t_L g2595 ( 
.A(n_2443),
.B(n_1991),
.Y(n_2595)
);

INVx4_ASAP7_75t_L g2596 ( 
.A(n_2163),
.Y(n_2596)
);

AOI21x1_ASAP7_75t_L g2597 ( 
.A1(n_2500),
.A2(n_2028),
.B(n_2019),
.Y(n_2597)
);

INVx1_ASAP7_75t_SL g2598 ( 
.A(n_2328),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2192),
.B(n_1887),
.Y(n_2599)
);

INVx4_ASAP7_75t_L g2600 ( 
.A(n_2163),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_SL g2601 ( 
.A(n_2426),
.B(n_1789),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2146),
.B(n_1909),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2146),
.B(n_1909),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_SL g2604 ( 
.A(n_2120),
.B(n_2125),
.Y(n_2604)
);

BUFx4f_ASAP7_75t_L g2605 ( 
.A(n_2484),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2149),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_SL g2607 ( 
.A(n_2245),
.B(n_1833),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2154),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2476),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2455),
.A2(n_2033),
.B1(n_2059),
.B2(n_1792),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2160),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2161),
.Y(n_2612)
);

AND2x2_ASAP7_75t_SL g2613 ( 
.A(n_2159),
.B(n_2090),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2476),
.Y(n_2614)
);

INVx1_ASAP7_75t_SL g2615 ( 
.A(n_2389),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2188),
.B(n_1943),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2487),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2162),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2164),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2167),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2188),
.B(n_1943),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2168),
.Y(n_2622)
);

INVx4_ASAP7_75t_L g2623 ( 
.A(n_2163),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2182),
.B(n_1841),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2318),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2455),
.Y(n_2626)
);

BUFx3_ASAP7_75t_L g2627 ( 
.A(n_2151),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2487),
.Y(n_2628)
);

INVx1_ASAP7_75t_SL g2629 ( 
.A(n_2403),
.Y(n_2629)
);

BUFx2_ASAP7_75t_L g2630 ( 
.A(n_2181),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2493),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2493),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2321),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2245),
.B(n_1883),
.Y(n_2634)
);

INVx4_ASAP7_75t_L g2635 ( 
.A(n_2218),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2375),
.B(n_1948),
.Y(n_2636)
);

OR2x6_ASAP7_75t_L g2637 ( 
.A(n_2158),
.B(n_2171),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2288),
.Y(n_2638)
);

AND2x6_ASAP7_75t_L g2639 ( 
.A(n_2457),
.B(n_1935),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2457),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2496),
.Y(n_2641)
);

BUFx6f_ASAP7_75t_L g2642 ( 
.A(n_2529),
.Y(n_2642)
);

INVx2_ASAP7_75t_SL g2643 ( 
.A(n_2325),
.Y(n_2643)
);

INVx2_ASAP7_75t_L g2644 ( 
.A(n_2496),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2288),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_2242),
.Y(n_2646)
);

OR2x6_ASAP7_75t_L g2647 ( 
.A(n_2438),
.B(n_1966),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2118),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2118),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_SL g2650 ( 
.A(n_2478),
.B(n_1889),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2288),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2344),
.B(n_1970),
.Y(n_2652)
);

INVx3_ASAP7_75t_L g2653 ( 
.A(n_2529),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_L g2654 ( 
.A(n_2456),
.B(n_1948),
.Y(n_2654)
);

INVxp33_ASAP7_75t_L g2655 ( 
.A(n_2404),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2131),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2119),
.Y(n_2657)
);

AOI22xp33_ASAP7_75t_L g2658 ( 
.A1(n_2480),
.A2(n_2059),
.B1(n_1792),
.B2(n_1990),
.Y(n_2658)
);

INVx1_ASAP7_75t_SL g2659 ( 
.A(n_2413),
.Y(n_2659)
);

INVx2_ASAP7_75t_SL g2660 ( 
.A(n_2131),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2119),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2131),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2122),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2205),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2205),
.Y(n_2665)
);

INVx2_ASAP7_75t_SL g2666 ( 
.A(n_2205),
.Y(n_2666)
);

INVx3_ASAP7_75t_L g2667 ( 
.A(n_2128),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2208),
.Y(n_2668)
);

INVx6_ASAP7_75t_L g2669 ( 
.A(n_2124),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2122),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_L g2671 ( 
.A(n_2456),
.B(n_1985),
.Y(n_2671)
);

INVx4_ASAP7_75t_L g2672 ( 
.A(n_2218),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2320),
.B(n_2194),
.Y(n_2673)
);

BUFx4f_ASAP7_75t_L g2674 ( 
.A(n_2201),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2213),
.B(n_1985),
.Y(n_2675)
);

INVx2_ASAP7_75t_SL g2676 ( 
.A(n_2208),
.Y(n_2676)
);

OAI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2217),
.A2(n_1993),
.B1(n_806),
.B2(n_808),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2208),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2368),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2130),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2130),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2478),
.B(n_2222),
.Y(n_2682)
);

BUFx10_ASAP7_75t_L g2683 ( 
.A(n_2304),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2445),
.B(n_1994),
.Y(n_2684)
);

INVx2_ASAP7_75t_SL g2685 ( 
.A(n_2519),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2373),
.Y(n_2686)
);

NAND2xp33_ASAP7_75t_L g2687 ( 
.A(n_2201),
.B(n_1891),
.Y(n_2687)
);

INVx3_ASAP7_75t_L g2688 ( 
.A(n_2128),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2155),
.B(n_2008),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2212),
.Y(n_2690)
);

AND3x2_ASAP7_75t_L g2691 ( 
.A(n_2190),
.B(n_1760),
.C(n_1993),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2374),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_SL g2693 ( 
.A(n_2256),
.B(n_1910),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2260),
.B(n_1946),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2376),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2212),
.Y(n_2696)
);

INVxp33_ASAP7_75t_SL g2697 ( 
.A(n_2343),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2214),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2214),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_2335),
.B(n_1994),
.Y(n_2700)
);

AND3x2_ASAP7_75t_L g2701 ( 
.A(n_2443),
.B(n_2086),
.C(n_2026),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2378),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2447),
.B(n_1997),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2460),
.B(n_1997),
.Y(n_2704)
);

AND2x4_ASAP7_75t_L g2705 ( 
.A(n_2271),
.B(n_2060),
.Y(n_2705)
);

NOR2xp33_ASAP7_75t_L g2706 ( 
.A(n_2520),
.B(n_2524),
.Y(n_2706)
);

XOR2xp5_ASAP7_75t_L g2707 ( 
.A(n_2437),
.B(n_1466),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2157),
.B(n_2018),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2172),
.B(n_2039),
.Y(n_2709)
);

NOR2x1_ASAP7_75t_L g2710 ( 
.A(n_2271),
.B(n_2039),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2216),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2173),
.B(n_2014),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2380),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2415),
.B(n_2014),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2129),
.B(n_2034),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2216),
.Y(n_2716)
);

NAND2xp33_ASAP7_75t_L g2717 ( 
.A(n_2201),
.B(n_1868),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2225),
.Y(n_2718)
);

AND2x4_ASAP7_75t_L g2719 ( 
.A(n_2223),
.B(n_2224),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2225),
.Y(n_2720)
);

INVx3_ASAP7_75t_L g2721 ( 
.A(n_2128),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2304),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2458),
.B(n_2046),
.Y(n_2723)
);

NOR2xp33_ASAP7_75t_L g2724 ( 
.A(n_2129),
.B(n_2046),
.Y(n_2724)
);

OAI22xp33_ASAP7_75t_L g2725 ( 
.A1(n_2360),
.A2(n_806),
.B1(n_808),
.B2(n_800),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2176),
.B(n_2186),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2227),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2227),
.Y(n_2728)
);

OAI22xp33_ASAP7_75t_SL g2729 ( 
.A1(n_2513),
.A2(n_1892),
.B1(n_1942),
.B2(n_1884),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_2153),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_2542),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2238),
.B(n_2060),
.Y(n_2732)
);

AOI22xp33_ASAP7_75t_L g2733 ( 
.A1(n_2480),
.A2(n_1904),
.B1(n_2092),
.B2(n_2096),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2231),
.Y(n_2734)
);

BUFx6f_ASAP7_75t_SL g2735 ( 
.A(n_2159),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2381),
.Y(n_2736)
);

INVx6_ASAP7_75t_L g2737 ( 
.A(n_2124),
.Y(n_2737)
);

BUFx3_ASAP7_75t_L g2738 ( 
.A(n_2502),
.Y(n_2738)
);

INVx4_ASAP7_75t_L g2739 ( 
.A(n_2506),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2231),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2258),
.B(n_2063),
.Y(n_2741)
);

INVx3_ASAP7_75t_L g2742 ( 
.A(n_2153),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2274),
.B(n_2063),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2137),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2137),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_2220),
.B(n_2066),
.Y(n_2746)
);

INVx2_ASAP7_75t_SL g2747 ( 
.A(n_2539),
.Y(n_2747)
);

NAND2xp33_ASAP7_75t_L g2748 ( 
.A(n_2201),
.B(n_1884),
.Y(n_2748)
);

AND3x2_ASAP7_75t_L g2749 ( 
.A(n_2474),
.B(n_1875),
.C(n_2066),
.Y(n_2749)
);

OR2x6_ASAP7_75t_L g2750 ( 
.A(n_2353),
.B(n_2000),
.Y(n_2750)
);

INVx2_ASAP7_75t_SL g2751 ( 
.A(n_2537),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_SL g2752 ( 
.A(n_2280),
.B(n_1892),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2141),
.Y(n_2753)
);

INVx2_ASAP7_75t_SL g2754 ( 
.A(n_2537),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2141),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2313),
.B(n_2201),
.Y(n_2756)
);

NOR2x1p5_ASAP7_75t_L g2757 ( 
.A(n_2542),
.B(n_1859),
.Y(n_2757)
);

INVx3_ASAP7_75t_L g2758 ( 
.A(n_2153),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2185),
.B(n_1942),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2279),
.B(n_1875),
.Y(n_2760)
);

AOI22xp5_ASAP7_75t_L g2761 ( 
.A1(n_2461),
.A2(n_2009),
.B1(n_2073),
.B2(n_2070),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2284),
.B(n_2015),
.Y(n_2762)
);

INVx1_ASAP7_75t_SL g2763 ( 
.A(n_2485),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2198),
.Y(n_2764)
);

AOI22xp33_ASAP7_75t_L g2765 ( 
.A1(n_2480),
.A2(n_2541),
.B1(n_2270),
.B2(n_2461),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2537),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2143),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2384),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2388),
.Y(n_2769)
);

BUFx8_ASAP7_75t_SL g2770 ( 
.A(n_2485),
.Y(n_2770)
);

INVx2_ASAP7_75t_SL g2771 ( 
.A(n_2223),
.Y(n_2771)
);

CKINVDCx6p67_ASAP7_75t_R g2772 ( 
.A(n_2209),
.Y(n_2772)
);

INVx2_ASAP7_75t_SL g2773 ( 
.A(n_2223),
.Y(n_2773)
);

BUFx2_ASAP7_75t_L g2774 ( 
.A(n_2181),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2143),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_SL g2776 ( 
.A(n_2135),
.B(n_2219),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2467),
.B(n_2469),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2392),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2185),
.B(n_2096),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2490),
.B(n_2048),
.Y(n_2780)
);

INVx2_ASAP7_75t_SL g2781 ( 
.A(n_2353),
.Y(n_2781)
);

AO22x2_ASAP7_75t_L g2782 ( 
.A1(n_2513),
.A2(n_1928),
.B1(n_1922),
.B2(n_2087),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2174),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2174),
.Y(n_2784)
);

INVx3_ASAP7_75t_L g2785 ( 
.A(n_2198),
.Y(n_2785)
);

CKINVDCx6p67_ASAP7_75t_R g2786 ( 
.A(n_2209),
.Y(n_2786)
);

INVx2_ASAP7_75t_SL g2787 ( 
.A(n_2382),
.Y(n_2787)
);

INVx3_ASAP7_75t_L g2788 ( 
.A(n_2198),
.Y(n_2788)
);

AOI22xp5_ASAP7_75t_L g2789 ( 
.A1(n_2330),
.A2(n_2076),
.B1(n_2079),
.B2(n_2075),
.Y(n_2789)
);

AND3x2_ASAP7_75t_L g2790 ( 
.A(n_2474),
.B(n_1571),
.C(n_1570),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2393),
.Y(n_2791)
);

INVxp33_ASAP7_75t_L g2792 ( 
.A(n_2210),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2285),
.B(n_2020),
.Y(n_2793)
);

OAI22xp33_ASAP7_75t_L g2794 ( 
.A1(n_2526),
.A2(n_811),
.B1(n_815),
.B2(n_809),
.Y(n_2794)
);

AND2x6_ASAP7_75t_L g2795 ( 
.A(n_2281),
.B(n_2032),
.Y(n_2795)
);

CKINVDCx5p33_ASAP7_75t_R g2796 ( 
.A(n_2124),
.Y(n_2796)
);

INVx5_ASAP7_75t_L g2797 ( 
.A(n_2533),
.Y(n_2797)
);

BUFx6f_ASAP7_75t_L g2798 ( 
.A(n_2138),
.Y(n_2798)
);

BUFx6f_ASAP7_75t_L g2799 ( 
.A(n_2138),
.Y(n_2799)
);

OAI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2515),
.A2(n_2020),
.B1(n_2052),
.B2(n_1930),
.Y(n_2800)
);

NAND3xp33_ASAP7_75t_L g2801 ( 
.A(n_2270),
.B(n_2527),
.C(n_2515),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2179),
.Y(n_2802)
);

NAND2xp33_ASAP7_75t_L g2803 ( 
.A(n_2330),
.B(n_2052),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_2527),
.B(n_2080),
.Y(n_2804)
);

INVx2_ASAP7_75t_SL g2805 ( 
.A(n_2382),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_2169),
.B(n_1762),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2396),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2179),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2401),
.Y(n_2809)
);

BUFx6f_ASAP7_75t_L g2810 ( 
.A(n_2138),
.Y(n_2810)
);

INVxp67_ASAP7_75t_L g2811 ( 
.A(n_2512),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2180),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2180),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2191),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2191),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2193),
.Y(n_2816)
);

INVx2_ASAP7_75t_SL g2817 ( 
.A(n_2410),
.Y(n_2817)
);

BUFx8_ASAP7_75t_SL g2818 ( 
.A(n_2150),
.Y(n_2818)
);

INVx6_ASAP7_75t_L g2819 ( 
.A(n_2150),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2193),
.Y(n_2820)
);

INVxp67_ASAP7_75t_SL g2821 ( 
.A(n_2541),
.Y(n_2821)
);

AND3x1_ASAP7_75t_L g2822 ( 
.A(n_2499),
.B(n_2531),
.C(n_2523),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2170),
.B(n_1762),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2203),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2453),
.A2(n_811),
.B1(n_815),
.B2(n_809),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2203),
.Y(n_2826)
);

BUFx2_ASAP7_75t_L g2827 ( 
.A(n_2210),
.Y(n_2827)
);

INVx2_ASAP7_75t_SL g2828 ( 
.A(n_2410),
.Y(n_2828)
);

INVx3_ASAP7_75t_L g2829 ( 
.A(n_2199),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2406),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_SL g2831 ( 
.A(n_2228),
.B(n_1762),
.Y(n_2831)
);

INVx3_ASAP7_75t_L g2832 ( 
.A(n_2199),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2507),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2507),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2411),
.Y(n_2835)
);

AOI22xp5_ASAP7_75t_L g2836 ( 
.A1(n_2330),
.A2(n_1906),
.B1(n_1772),
.B2(n_1776),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2510),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2414),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2510),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_2150),
.Y(n_2840)
);

BUFx6f_ASAP7_75t_L g2841 ( 
.A(n_2138),
.Y(n_2841)
);

INVx1_ASAP7_75t_SL g2842 ( 
.A(n_2430),
.Y(n_2842)
);

CKINVDCx5p33_ASAP7_75t_R g2843 ( 
.A(n_2282),
.Y(n_2843)
);

BUFx6f_ASAP7_75t_L g2844 ( 
.A(n_2152),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2298),
.B(n_1930),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2514),
.Y(n_2846)
);

INVxp33_ASAP7_75t_L g2847 ( 
.A(n_2267),
.Y(n_2847)
);

AND2x6_ASAP7_75t_L g2848 ( 
.A(n_2134),
.B(n_2040),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2416),
.Y(n_2849)
);

BUFx6f_ASAP7_75t_L g2850 ( 
.A(n_2152),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2199),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2420),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2514),
.Y(n_2853)
);

NAND2xp33_ASAP7_75t_R g2854 ( 
.A(n_2431),
.B(n_819),
.Y(n_2854)
);

OAI21xp33_ASAP7_75t_SL g2855 ( 
.A1(n_2298),
.A2(n_2027),
.B(n_1574),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2532),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2428),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2330),
.A2(n_2043),
.B1(n_2045),
.B2(n_2042),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2430),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2429),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_L g2861 ( 
.A(n_2235),
.B(n_954),
.Y(n_2861)
);

INVx2_ASAP7_75t_SL g2862 ( 
.A(n_2267),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_SL g2863 ( 
.A(n_2237),
.B(n_2240),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2286),
.B(n_2054),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2287),
.B(n_2067),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2532),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2546),
.Y(n_2867)
);

INVx1_ASAP7_75t_SL g2868 ( 
.A(n_2317),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2432),
.Y(n_2869)
);

CKINVDCx20_ASAP7_75t_R g2870 ( 
.A(n_2282),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2546),
.Y(n_2871)
);

NOR2xp33_ASAP7_75t_L g2872 ( 
.A(n_2246),
.B(n_955),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2422),
.Y(n_2873)
);

CKINVDCx5p33_ASAP7_75t_R g2874 ( 
.A(n_2282),
.Y(n_2874)
);

AND2x4_ASAP7_75t_L g2875 ( 
.A(n_2254),
.B(n_1573),
.Y(n_2875)
);

INVx4_ASAP7_75t_L g2876 ( 
.A(n_2506),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2433),
.Y(n_2877)
);

NOR2xp33_ASAP7_75t_L g2878 ( 
.A(n_2255),
.B(n_956),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2422),
.Y(n_2879)
);

INVx3_ASAP7_75t_L g2880 ( 
.A(n_2226),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2422),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2440),
.Y(n_2882)
);

BUFx4f_ASAP7_75t_L g2883 ( 
.A(n_2330),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2248),
.Y(n_2884)
);

NAND3xp33_ASAP7_75t_L g2885 ( 
.A(n_2283),
.B(n_961),
.C(n_958),
.Y(n_2885)
);

BUFx6f_ASAP7_75t_L g2886 ( 
.A(n_2152),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2293),
.B(n_2084),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2257),
.B(n_962),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2453),
.A2(n_823),
.B1(n_824),
.B2(n_819),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2297),
.Y(n_2890)
);

INVx8_ASAP7_75t_L g2891 ( 
.A(n_2407),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2301),
.Y(n_2892)
);

INVx4_ASAP7_75t_L g2893 ( 
.A(n_2506),
.Y(n_2893)
);

BUFx4f_ASAP7_75t_L g2894 ( 
.A(n_2407),
.Y(n_2894)
);

INVx5_ASAP7_75t_L g2895 ( 
.A(n_2533),
.Y(n_2895)
);

INVx4_ASAP7_75t_L g2896 ( 
.A(n_2506),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2303),
.Y(n_2897)
);

OAI22xp33_ASAP7_75t_L g2898 ( 
.A1(n_2512),
.A2(n_2531),
.B1(n_2523),
.B2(n_2317),
.Y(n_2898)
);

AOI22xp33_ASAP7_75t_L g2899 ( 
.A1(n_2453),
.A2(n_824),
.B1(n_826),
.B2(n_823),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_SL g2900 ( 
.A(n_2259),
.B(n_2100),
.Y(n_2900)
);

BUFx2_ASAP7_75t_L g2901 ( 
.A(n_2337),
.Y(n_2901)
);

AOI22xp33_ASAP7_75t_L g2902 ( 
.A1(n_2453),
.A2(n_830),
.B1(n_836),
.B2(n_826),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2308),
.Y(n_2903)
);

INVx4_ASAP7_75t_L g2904 ( 
.A(n_2525),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2453),
.A2(n_836),
.B1(n_838),
.B2(n_830),
.Y(n_2905)
);

AND3x2_ASAP7_75t_L g2906 ( 
.A(n_2337),
.B(n_1580),
.C(n_1577),
.Y(n_2906)
);

INVx2_ASAP7_75t_SL g2907 ( 
.A(n_2262),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2311),
.Y(n_2908)
);

BUFx4f_ASAP7_75t_L g2909 ( 
.A(n_2407),
.Y(n_2909)
);

INVx3_ASAP7_75t_L g2910 ( 
.A(n_2226),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2312),
.B(n_2101),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2407),
.B(n_2104),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2450),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2407),
.B(n_2105),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2525),
.Y(n_2915)
);

BUFx3_ASAP7_75t_L g2916 ( 
.A(n_2264),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2452),
.B(n_1912),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2454),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2459),
.B(n_1916),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_SL g2920 ( 
.A(n_2265),
.B(n_1983),
.Y(n_2920)
);

INVx2_ASAP7_75t_L g2921 ( 
.A(n_2462),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2492),
.Y(n_2922)
);

AOI21x1_ASAP7_75t_L g2923 ( 
.A1(n_2175),
.A2(n_1929),
.B(n_2027),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2266),
.Y(n_2924)
);

CKINVDCx5p33_ASAP7_75t_R g2925 ( 
.A(n_2310),
.Y(n_2925)
);

INVx3_ASAP7_75t_L g2926 ( 
.A(n_2226),
.Y(n_2926)
);

NOR2xp33_ASAP7_75t_L g2927 ( 
.A(n_2268),
.B(n_964),
.Y(n_2927)
);

AND2x4_ASAP7_75t_L g2928 ( 
.A(n_2272),
.B(n_1581),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_SL g2929 ( 
.A(n_2273),
.B(n_1983),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2275),
.B(n_969),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2277),
.B(n_970),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2248),
.Y(n_2932)
);

BUFx6f_ASAP7_75t_SL g2933 ( 
.A(n_2329),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2249),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2195),
.B(n_1923),
.Y(n_2935)
);

AND3x2_ASAP7_75t_L g2936 ( 
.A(n_2329),
.B(n_1584),
.C(n_1583),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2196),
.B(n_1923),
.Y(n_2937)
);

BUFx6f_ASAP7_75t_SL g2938 ( 
.A(n_2329),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2249),
.Y(n_2939)
);

HB1xp67_ASAP7_75t_L g2940 ( 
.A(n_2339),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2339),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2339),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2345),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2250),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2250),
.Y(n_2945)
);

NAND2xp33_ASAP7_75t_SL g2946 ( 
.A(n_2232),
.B(n_2251),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2345),
.Y(n_2947)
);

BUFx6f_ASAP7_75t_L g2948 ( 
.A(n_2152),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_2252),
.B(n_2030),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2345),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2252),
.Y(n_2951)
);

AND2x2_ASAP7_75t_SL g2952 ( 
.A(n_2346),
.B(n_1585),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2290),
.B(n_2030),
.Y(n_2953)
);

NAND3xp33_ASAP7_75t_L g2954 ( 
.A(n_2347),
.B(n_972),
.C(n_971),
.Y(n_2954)
);

BUFx2_ASAP7_75t_L g2955 ( 
.A(n_2183),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_2290),
.B(n_2030),
.Y(n_2956)
);

INVx2_ASAP7_75t_SL g2957 ( 
.A(n_2346),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_SL g2958 ( 
.A(n_2291),
.B(n_2030),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2346),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2291),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2349),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2349),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2295),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2232),
.B(n_974),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2295),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2349),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2296),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2251),
.B(n_982),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2200),
.B(n_1923),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2296),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2302),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2204),
.B(n_1925),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2207),
.B(n_1925),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_SL g2974 ( 
.A(n_2302),
.B(n_2037),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2306),
.Y(n_2975)
);

INVx1_ASAP7_75t_SL g2976 ( 
.A(n_2477),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2354),
.Y(n_2977)
);

INVx5_ASAP7_75t_L g2978 ( 
.A(n_2533),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2211),
.B(n_1925),
.Y(n_2979)
);

NAND2xp33_ASAP7_75t_SL g2980 ( 
.A(n_2305),
.B(n_838),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2354),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2221),
.B(n_1925),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2833),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2777),
.B(n_2354),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2574),
.B(n_2399),
.Y(n_2985)
);

AND2x6_ASAP7_75t_L g2986 ( 
.A(n_2563),
.B(n_2305),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2726),
.B(n_2306),
.Y(n_2987)
);

AND2x6_ASAP7_75t_L g2988 ( 
.A(n_2563),
.B(n_2314),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2575),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2833),
.Y(n_2990)
);

BUFx3_ASAP7_75t_L g2991 ( 
.A(n_2572),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2626),
.B(n_2314),
.Y(n_2992)
);

AND2x4_ASAP7_75t_L g2993 ( 
.A(n_2568),
.B(n_2399),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2626),
.B(n_2319),
.Y(n_2994)
);

AND2x4_ASAP7_75t_L g2995 ( 
.A(n_2568),
.B(n_2627),
.Y(n_2995)
);

INVx8_ASAP7_75t_L g2996 ( 
.A(n_2933),
.Y(n_2996)
);

INVx4_ASAP7_75t_L g2997 ( 
.A(n_2563),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2834),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2673),
.B(n_2319),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2653),
.B(n_2322),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2834),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2837),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2837),
.Y(n_3003)
);

AND2x4_ASAP7_75t_L g3004 ( 
.A(n_2627),
.B(n_2751),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2563),
.Y(n_3005)
);

AND2x4_ASAP7_75t_L g3006 ( 
.A(n_2754),
.B(n_2399),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2853),
.Y(n_3007)
);

INVx4_ASAP7_75t_L g3008 ( 
.A(n_2589),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2853),
.Y(n_3009)
);

NOR2xp33_ASAP7_75t_L g3010 ( 
.A(n_2654),
.B(n_1475),
.Y(n_3010)
);

INVxp67_ASAP7_75t_L g3011 ( 
.A(n_2591),
.Y(n_3011)
);

AND2x4_ASAP7_75t_L g3012 ( 
.A(n_2766),
.B(n_2435),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2571),
.A2(n_2431),
.B1(n_2544),
.B2(n_2435),
.Y(n_3013)
);

INVx3_ASAP7_75t_L g3014 ( 
.A(n_2589),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2624),
.B(n_2615),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2629),
.B(n_2435),
.Y(n_3016)
);

INVxp67_ASAP7_75t_SL g3017 ( 
.A(n_2589),
.Y(n_3017)
);

INVx2_ASAP7_75t_SL g3018 ( 
.A(n_2573),
.Y(n_3018)
);

AO22x2_ASAP7_75t_L g3019 ( 
.A1(n_2560),
.A2(n_1800),
.B1(n_1880),
.B2(n_1763),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2659),
.B(n_1492),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2575),
.Y(n_3021)
);

AO21x2_ASAP7_75t_L g3022 ( 
.A1(n_2561),
.A2(n_2126),
.B(n_2498),
.Y(n_3022)
);

INVx1_ASAP7_75t_SL g3023 ( 
.A(n_2868),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2856),
.Y(n_3024)
);

NAND3xp33_ASAP7_75t_L g3025 ( 
.A(n_2759),
.B(n_2479),
.C(n_2472),
.Y(n_3025)
);

NOR2xp33_ASAP7_75t_L g3026 ( 
.A(n_2654),
.B(n_1492),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2653),
.B(n_2322),
.Y(n_3027)
);

BUFx3_ASAP7_75t_L g3028 ( 
.A(n_2738),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2856),
.Y(n_3029)
);

AND2x4_ASAP7_75t_L g3030 ( 
.A(n_2660),
.B(n_2327),
.Y(n_3030)
);

AO22x2_ASAP7_75t_L g3031 ( 
.A1(n_2707),
.A2(n_1493),
.B1(n_1499),
.B2(n_1495),
.Y(n_3031)
);

AND2x4_ASAP7_75t_L g3032 ( 
.A(n_2666),
.B(n_2327),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2577),
.B(n_2340),
.Y(n_3033)
);

INVx4_ASAP7_75t_L g3034 ( 
.A(n_2589),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2617),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2866),
.Y(n_3036)
);

AND2x4_ASAP7_75t_L g3037 ( 
.A(n_2676),
.B(n_2340),
.Y(n_3037)
);

INVx4_ASAP7_75t_L g3038 ( 
.A(n_2640),
.Y(n_3038)
);

INVx4_ASAP7_75t_L g3039 ( 
.A(n_2640),
.Y(n_3039)
);

AND2x6_ASAP7_75t_L g3040 ( 
.A(n_2640),
.B(n_2355),
.Y(n_3040)
);

NOR2xp33_ASAP7_75t_L g3041 ( 
.A(n_2671),
.B(n_1493),
.Y(n_3041)
);

OR2x6_ASAP7_75t_L g3042 ( 
.A(n_2669),
.B(n_1768),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2617),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2866),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2867),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2675),
.B(n_2355),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2867),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2871),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2640),
.Y(n_3049)
);

AND2x4_ASAP7_75t_L g3050 ( 
.A(n_2771),
.B(n_2357),
.Y(n_3050)
);

BUFx6f_ASAP7_75t_L g3051 ( 
.A(n_2642),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2642),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2952),
.B(n_2269),
.Y(n_3053)
);

HB1xp67_ASAP7_75t_L g3054 ( 
.A(n_2630),
.Y(n_3054)
);

OAI22xp5_ASAP7_75t_L g3055 ( 
.A1(n_2610),
.A2(n_2658),
.B1(n_2571),
.B2(n_2580),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2652),
.B(n_1495),
.Y(n_3056)
);

NOR2xp33_ASAP7_75t_L g3057 ( 
.A(n_2671),
.B(n_1499),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2548),
.B(n_1536),
.Y(n_3058)
);

INVx4_ASAP7_75t_L g3059 ( 
.A(n_2642),
.Y(n_3059)
);

INVx4_ASAP7_75t_L g3060 ( 
.A(n_2642),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2675),
.B(n_2357),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2712),
.B(n_2358),
.Y(n_3062)
);

INVx2_ASAP7_75t_SL g3063 ( 
.A(n_2774),
.Y(n_3063)
);

AND2x6_ASAP7_75t_L g3064 ( 
.A(n_2873),
.B(n_2358),
.Y(n_3064)
);

BUFx6f_ASAP7_75t_L g3065 ( 
.A(n_2798),
.Y(n_3065)
);

INVx4_ASAP7_75t_L g3066 ( 
.A(n_2596),
.Y(n_3066)
);

BUFx6f_ASAP7_75t_L g3067 ( 
.A(n_2798),
.Y(n_3067)
);

INVx5_ASAP7_75t_L g3068 ( 
.A(n_2639),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2631),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2584),
.B(n_2367),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2689),
.B(n_1536),
.Y(n_3071)
);

INVx5_ASAP7_75t_L g3072 ( 
.A(n_2639),
.Y(n_3072)
);

BUFx2_ASAP7_75t_L g3073 ( 
.A(n_2827),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2602),
.B(n_1556),
.Y(n_3074)
);

OR2x2_ASAP7_75t_SL g3075 ( 
.A(n_2636),
.B(n_1556),
.Y(n_3075)
);

CKINVDCx20_ASAP7_75t_R g3076 ( 
.A(n_2770),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2871),
.Y(n_3077)
);

BUFx10_ASAP7_75t_L g3078 ( 
.A(n_2804),
.Y(n_3078)
);

NOR2x1p5_ASAP7_75t_L g3079 ( 
.A(n_2616),
.B(n_2310),
.Y(n_3079)
);

INVx4_ASAP7_75t_L g3080 ( 
.A(n_2596),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_2547),
.B(n_1579),
.Y(n_3081)
);

AND2x4_ASAP7_75t_L g3082 ( 
.A(n_2773),
.B(n_2367),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2783),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2783),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_SL g3085 ( 
.A(n_2952),
.B(n_2333),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2784),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2784),
.Y(n_3087)
);

AND2x4_ASAP7_75t_L g3088 ( 
.A(n_2643),
.B(n_2377),
.Y(n_3088)
);

AO21x2_ASAP7_75t_L g3089 ( 
.A1(n_2682),
.A2(n_2604),
.B(n_2803),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2802),
.Y(n_3090)
);

NAND2x1p5_ASAP7_75t_L g3091 ( 
.A(n_2600),
.B(n_2543),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2802),
.Y(n_3092)
);

BUFx6f_ASAP7_75t_L g3093 ( 
.A(n_2798),
.Y(n_3093)
);

BUFx3_ASAP7_75t_L g3094 ( 
.A(n_2738),
.Y(n_3094)
);

AND2x4_ASAP7_75t_L g3095 ( 
.A(n_2719),
.B(n_2377),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_2547),
.B(n_1579),
.Y(n_3096)
);

NAND2x1p5_ASAP7_75t_L g3097 ( 
.A(n_2600),
.B(n_2543),
.Y(n_3097)
);

BUFx6f_ASAP7_75t_SL g3098 ( 
.A(n_2579),
.Y(n_3098)
);

BUFx6f_ASAP7_75t_L g3099 ( 
.A(n_2798),
.Y(n_3099)
);

OR2x2_ASAP7_75t_SL g3100 ( 
.A(n_2621),
.B(n_1600),
.Y(n_3100)
);

NOR2xp33_ASAP7_75t_L g3101 ( 
.A(n_2602),
.B(n_1600),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2603),
.B(n_1601),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_SL g3103 ( 
.A(n_2603),
.B(n_2333),
.Y(n_3103)
);

HB1xp67_ASAP7_75t_L g3104 ( 
.A(n_2901),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2655),
.B(n_2714),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2808),
.Y(n_3106)
);

NOR2xp33_ASAP7_75t_L g3107 ( 
.A(n_2584),
.B(n_1601),
.Y(n_3107)
);

OAI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_2610),
.A2(n_2658),
.B1(n_2571),
.B2(n_2585),
.Y(n_3108)
);

BUFx2_ASAP7_75t_L g3109 ( 
.A(n_2598),
.Y(n_3109)
);

INVx2_ASAP7_75t_SL g3110 ( 
.A(n_2862),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_2719),
.B(n_2379),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2808),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2759),
.B(n_2379),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2704),
.B(n_2383),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_2655),
.B(n_1611),
.Y(n_3115)
);

OR2x2_ASAP7_75t_L g3116 ( 
.A(n_2595),
.B(n_2842),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2587),
.B(n_2333),
.Y(n_3117)
);

INVx1_ASAP7_75t_SL g3118 ( 
.A(n_2723),
.Y(n_3118)
);

NOR2xp33_ASAP7_75t_L g3119 ( 
.A(n_2599),
.B(n_1611),
.Y(n_3119)
);

INVx3_ASAP7_75t_L g3120 ( 
.A(n_2667),
.Y(n_3120)
);

AND2x2_ASAP7_75t_SL g3121 ( 
.A(n_2613),
.B(n_1973),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2812),
.Y(n_3122)
);

BUFx10_ASAP7_75t_L g3123 ( 
.A(n_2804),
.Y(n_3123)
);

AND2x4_ASAP7_75t_L g3124 ( 
.A(n_2635),
.B(n_2383),
.Y(n_3124)
);

NAND2xp33_ASAP7_75t_L g3125 ( 
.A(n_2891),
.B(n_2544),
.Y(n_3125)
);

AND2x4_ASAP7_75t_L g3126 ( 
.A(n_2635),
.B(n_2386),
.Y(n_3126)
);

BUFx6f_ASAP7_75t_L g3127 ( 
.A(n_2799),
.Y(n_3127)
);

AND2x4_ASAP7_75t_SL g3128 ( 
.A(n_2579),
.B(n_1623),
.Y(n_3128)
);

INVx3_ASAP7_75t_L g3129 ( 
.A(n_2667),
.Y(n_3129)
);

BUFx6f_ASAP7_75t_L g3130 ( 
.A(n_2799),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2812),
.Y(n_3131)
);

BUFx3_ASAP7_75t_L g3132 ( 
.A(n_2770),
.Y(n_3132)
);

BUFx3_ASAP7_75t_L g3133 ( 
.A(n_2781),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2813),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2813),
.Y(n_3135)
);

OAI22xp5_ASAP7_75t_SL g3136 ( 
.A1(n_2613),
.A2(n_1651),
.B1(n_1654),
.B2(n_1623),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2814),
.Y(n_3137)
);

CKINVDCx11_ASAP7_75t_R g3138 ( 
.A(n_2570),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2814),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2815),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2815),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_L g3142 ( 
.A(n_2704),
.B(n_1651),
.Y(n_3142)
);

AOI22xp5_ASAP7_75t_L g3143 ( 
.A1(n_2980),
.A2(n_2544),
.B1(n_2387),
.B2(n_2394),
.Y(n_3143)
);

INVx3_ASAP7_75t_L g3144 ( 
.A(n_2688),
.Y(n_3144)
);

AND2x2_ASAP7_75t_L g3145 ( 
.A(n_2706),
.B(n_1654),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2631),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2816),
.Y(n_3147)
);

NOR2xp33_ASAP7_75t_L g3148 ( 
.A(n_2684),
.B(n_1655),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2787),
.Y(n_3149)
);

INVx3_ASAP7_75t_L g3150 ( 
.A(n_2688),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2632),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_SL g3152 ( 
.A(n_2703),
.B(n_2333),
.Y(n_3152)
);

AND2x4_ASAP7_75t_L g3153 ( 
.A(n_2672),
.B(n_2705),
.Y(n_3153)
);

NAND3xp33_ASAP7_75t_L g3154 ( 
.A(n_2776),
.B(n_2495),
.C(n_2486),
.Y(n_3154)
);

INVx1_ASAP7_75t_SL g3155 ( 
.A(n_2805),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_2706),
.B(n_2792),
.Y(n_3156)
);

HB1xp67_ASAP7_75t_L g3157 ( 
.A(n_2817),
.Y(n_3157)
);

INVxp33_ASAP7_75t_SL g3158 ( 
.A(n_2646),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2816),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2709),
.B(n_2386),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_2776),
.A2(n_2639),
.B1(n_2752),
.B2(n_2801),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2820),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2632),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2820),
.Y(n_3164)
);

OR2x2_ASAP7_75t_L g3165 ( 
.A(n_2811),
.B(n_2522),
.Y(n_3165)
);

AND2x4_ASAP7_75t_L g3166 ( 
.A(n_2672),
.B(n_2387),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2824),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2641),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2824),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2826),
.Y(n_3170)
);

NOR2x1p5_ASAP7_75t_L g3171 ( 
.A(n_2772),
.B(n_2310),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2800),
.B(n_2405),
.Y(n_3172)
);

INVx5_ASAP7_75t_L g3173 ( 
.A(n_2639),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2826),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2940),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2700),
.B(n_2405),
.Y(n_3176)
);

BUFx2_ASAP7_75t_L g3177 ( 
.A(n_2811),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2729),
.B(n_2394),
.Y(n_3178)
);

AND2x6_ASAP7_75t_L g3179 ( 
.A(n_2873),
.B(n_2418),
.Y(n_3179)
);

HB1xp67_ASAP7_75t_L g3180 ( 
.A(n_2828),
.Y(n_3180)
);

BUFx6f_ASAP7_75t_L g3181 ( 
.A(n_2799),
.Y(n_3181)
);

INVx5_ASAP7_75t_L g3182 ( 
.A(n_2639),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2641),
.Y(n_3183)
);

BUFx6f_ASAP7_75t_L g3184 ( 
.A(n_2799),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2940),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2690),
.Y(n_3186)
);

AO21x2_ASAP7_75t_L g3187 ( 
.A1(n_2682),
.A2(n_2604),
.B(n_2717),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_2845),
.B(n_2418),
.Y(n_3188)
);

INVx3_ASAP7_75t_L g3189 ( 
.A(n_2721),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_2792),
.B(n_1655),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2690),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2644),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2845),
.B(n_2421),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_2847),
.B(n_2780),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2644),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_SL g3196 ( 
.A(n_2674),
.B(n_2397),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_2700),
.B(n_2370),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2744),
.Y(n_3198)
);

AOI22xp33_ASAP7_75t_L g3199 ( 
.A1(n_2752),
.A2(n_2544),
.B1(n_2425),
.B2(n_2434),
.Y(n_3199)
);

OR2x2_ASAP7_75t_SL g3200 ( 
.A(n_2885),
.B(n_1686),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2745),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_2582),
.B(n_2370),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_L g3203 ( 
.A(n_2847),
.B(n_2708),
.Y(n_3203)
);

NOR2xp33_ASAP7_75t_L g3204 ( 
.A(n_2708),
.B(n_1686),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2753),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2755),
.Y(n_3206)
);

AOI22xp33_ASAP7_75t_L g3207 ( 
.A1(n_2825),
.A2(n_2544),
.B1(n_2425),
.B2(n_2434),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2767),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2775),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2551),
.B(n_2421),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2696),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_2859),
.B(n_1725),
.Y(n_3212)
);

INVx5_ASAP7_75t_L g3213 ( 
.A(n_2810),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_L g3214 ( 
.A(n_2594),
.B(n_1725),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2648),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_L g3216 ( 
.A(n_2594),
.B(n_1973),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2698),
.Y(n_3217)
);

BUFx2_ASAP7_75t_L g3218 ( 
.A(n_2763),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2699),
.Y(n_3219)
);

AND2x4_ASAP7_75t_L g3220 ( 
.A(n_2705),
.B(n_2436),
.Y(n_3220)
);

BUFx6f_ASAP7_75t_L g3221 ( 
.A(n_2810),
.Y(n_3221)
);

BUFx10_ASAP7_75t_L g3222 ( 
.A(n_2715),
.Y(n_3222)
);

HB1xp67_ASAP7_75t_L g3223 ( 
.A(n_2685),
.Y(n_3223)
);

AOI22xp33_ASAP7_75t_L g3224 ( 
.A1(n_2825),
.A2(n_2444),
.B1(n_2446),
.B2(n_2436),
.Y(n_3224)
);

AND2x4_ASAP7_75t_L g3225 ( 
.A(n_2957),
.B(n_2444),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2648),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_SL g3227 ( 
.A(n_2715),
.B(n_2370),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_2889),
.A2(n_2448),
.B1(n_2451),
.B2(n_2446),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2711),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2716),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2649),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2649),
.Y(n_3232)
);

AND2x6_ASAP7_75t_L g3233 ( 
.A(n_2879),
.B(n_2881),
.Y(n_3233)
);

AO22x2_ASAP7_75t_L g3234 ( 
.A1(n_2590),
.A2(n_2062),
.B1(n_2081),
.B2(n_2035),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_2593),
.B(n_1832),
.Y(n_3235)
);

CKINVDCx20_ASAP7_75t_R g3236 ( 
.A(n_2818),
.Y(n_3236)
);

BUFx4f_ASAP7_75t_L g3237 ( 
.A(n_2669),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_SL g3238 ( 
.A(n_2724),
.B(n_2370),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2657),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2657),
.Y(n_3240)
);

BUFx6f_ASAP7_75t_L g3241 ( 
.A(n_2810),
.Y(n_3241)
);

BUFx3_ASAP7_75t_L g3242 ( 
.A(n_2605),
.Y(n_3242)
);

OR2x6_ASAP7_75t_L g3243 ( 
.A(n_2669),
.B(n_2397),
.Y(n_3243)
);

BUFx6f_ASAP7_75t_L g3244 ( 
.A(n_2810),
.Y(n_3244)
);

AND2x4_ASAP7_75t_L g3245 ( 
.A(n_2916),
.B(n_2448),
.Y(n_3245)
);

INVx4_ASAP7_75t_SL g3246 ( 
.A(n_2737),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2718),
.Y(n_3247)
);

AND2x2_ASAP7_75t_SL g3248 ( 
.A(n_2889),
.B(n_2899),
.Y(n_3248)
);

INVx1_ASAP7_75t_SL g3249 ( 
.A(n_2946),
.Y(n_3249)
);

BUFx3_ASAP7_75t_L g3250 ( 
.A(n_2605),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2720),
.Y(n_3251)
);

BUFx6f_ASAP7_75t_L g3252 ( 
.A(n_2841),
.Y(n_3252)
);

AND2x4_ASAP7_75t_L g3253 ( 
.A(n_2916),
.B(n_2451),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2551),
.B(n_2465),
.Y(n_3254)
);

HB1xp67_ASAP7_75t_L g3255 ( 
.A(n_2747),
.Y(n_3255)
);

NAND3x1_ASAP7_75t_L g3256 ( 
.A(n_2761),
.B(n_1835),
.C(n_1831),
.Y(n_3256)
);

AND2x2_ASAP7_75t_L g3257 ( 
.A(n_2964),
.B(n_1832),
.Y(n_3257)
);

BUFx6f_ASAP7_75t_L g3258 ( 
.A(n_2841),
.Y(n_3258)
);

OR2x2_ASAP7_75t_L g3259 ( 
.A(n_2898),
.B(n_1851),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2661),
.Y(n_3260)
);

BUFx6f_ASAP7_75t_L g3261 ( 
.A(n_2841),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2552),
.B(n_2465),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2727),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2661),
.Y(n_3264)
);

BUFx6f_ASAP7_75t_L g3265 ( 
.A(n_2841),
.Y(n_3265)
);

INVx2_ASAP7_75t_SL g3266 ( 
.A(n_2790),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_SL g3267 ( 
.A(n_2724),
.B(n_2400),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_2721),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2728),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_2964),
.B(n_1851),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2734),
.Y(n_3271)
);

AND2x4_ASAP7_75t_L g3272 ( 
.A(n_2638),
.B(n_2498),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2740),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2663),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2663),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_2968),
.B(n_1587),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_2590),
.B(n_2400),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2552),
.B(n_2494),
.Y(n_3278)
);

AND3x1_ASAP7_75t_L g3279 ( 
.A(n_2733),
.B(n_1596),
.C(n_1593),
.Y(n_3279)
);

BUFx6f_ASAP7_75t_L g3280 ( 
.A(n_2844),
.Y(n_3280)
);

NOR2xp33_ASAP7_75t_L g3281 ( 
.A(n_2601),
.B(n_2035),
.Y(n_3281)
);

NOR2xp33_ASAP7_75t_L g3282 ( 
.A(n_2601),
.B(n_2062),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2670),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2670),
.Y(n_3284)
);

INVx4_ASAP7_75t_L g3285 ( 
.A(n_2623),
.Y(n_3285)
);

INVx5_ASAP7_75t_L g3286 ( 
.A(n_2844),
.Y(n_3286)
);

AND2x4_ASAP7_75t_L g3287 ( 
.A(n_2645),
.B(n_2651),
.Y(n_3287)
);

BUFx6f_ASAP7_75t_L g3288 ( 
.A(n_2844),
.Y(n_3288)
);

AOI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2748),
.A2(n_2475),
.B1(n_2481),
.B2(n_2466),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2554),
.B(n_2494),
.Y(n_3290)
);

AND2x4_ASAP7_75t_L g3291 ( 
.A(n_2656),
.B(n_1597),
.Y(n_3291)
);

OR2x2_ASAP7_75t_L g3292 ( 
.A(n_2898),
.B(n_1598),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_2968),
.B(n_1599),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2680),
.Y(n_3294)
);

CKINVDCx20_ASAP7_75t_R g3295 ( 
.A(n_2818),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_2693),
.B(n_2081),
.Y(n_3296)
);

BUFx3_ASAP7_75t_L g3297 ( 
.A(n_2875),
.Y(n_3297)
);

AND2x4_ASAP7_75t_L g3298 ( 
.A(n_2662),
.B(n_1602),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_2680),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2681),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2681),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_2839),
.Y(n_3302)
);

AND2x2_ASAP7_75t_L g3303 ( 
.A(n_2779),
.B(n_1603),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_2884),
.Y(n_3304)
);

INVx1_ASAP7_75t_SL g3305 ( 
.A(n_2976),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_2884),
.Y(n_3306)
);

BUFx3_ASAP7_75t_L g3307 ( 
.A(n_2875),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_2932),
.Y(n_3308)
);

NAND3xp33_ASAP7_75t_L g3309 ( 
.A(n_2585),
.B(n_2576),
.C(n_2733),
.Y(n_3309)
);

INVx3_ASAP7_75t_L g3310 ( 
.A(n_2730),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_2932),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_2846),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2553),
.Y(n_3313)
);

AND2x4_ASAP7_75t_L g3314 ( 
.A(n_2664),
.B(n_1604),
.Y(n_3314)
);

NOR2xp33_ASAP7_75t_L g3315 ( 
.A(n_2693),
.B(n_2083),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2557),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2558),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2554),
.B(n_2494),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2762),
.B(n_2503),
.Y(n_3319)
);

INVx3_ASAP7_75t_L g3320 ( 
.A(n_2730),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2564),
.Y(n_3321)
);

OAI22xp33_ASAP7_75t_SL g3322 ( 
.A1(n_2694),
.A2(n_844),
.B1(n_845),
.B2(n_841),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_SL g3323 ( 
.A(n_2822),
.B(n_2400),
.Y(n_3323)
);

AND2x4_ASAP7_75t_L g3324 ( 
.A(n_2665),
.B(n_1605),
.Y(n_3324)
);

BUFx6f_ASAP7_75t_SL g3325 ( 
.A(n_2683),
.Y(n_3325)
);

CKINVDCx5p33_ASAP7_75t_R g3326 ( 
.A(n_2722),
.Y(n_3326)
);

INVx2_ASAP7_75t_SL g3327 ( 
.A(n_2790),
.Y(n_3327)
);

NAND2xp33_ASAP7_75t_L g3328 ( 
.A(n_2891),
.B(n_2400),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2793),
.B(n_2503),
.Y(n_3329)
);

CKINVDCx5p33_ASAP7_75t_R g3330 ( 
.A(n_2731),
.Y(n_3330)
);

AND2x4_ASAP7_75t_L g3331 ( 
.A(n_2668),
.B(n_2678),
.Y(n_3331)
);

AO22x2_ASAP7_75t_L g3332 ( 
.A1(n_2694),
.A2(n_2098),
.B1(n_2083),
.B2(n_1607),
.Y(n_3332)
);

INVx2_ASAP7_75t_SL g3333 ( 
.A(n_2906),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2732),
.B(n_2503),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_L g3335 ( 
.A(n_2779),
.B(n_2098),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2576),
.B(n_2482),
.Y(n_3336)
);

NAND2x1p5_ASAP7_75t_L g3337 ( 
.A(n_2623),
.B(n_2528),
.Y(n_3337)
);

BUFx2_ASAP7_75t_L g3338 ( 
.A(n_2855),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_2934),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_2955),
.B(n_1609),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_2566),
.Y(n_3341)
);

INVxp67_ASAP7_75t_L g3342 ( 
.A(n_2861),
.Y(n_3342)
);

NOR2xp33_ASAP7_75t_L g3343 ( 
.A(n_2650),
.B(n_1881),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2578),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2581),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2583),
.Y(n_3346)
);

BUFx3_ASAP7_75t_L g3347 ( 
.A(n_2928),
.Y(n_3347)
);

AND2x4_ASAP7_75t_L g3348 ( 
.A(n_2941),
.B(n_1612),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_2934),
.Y(n_3349)
);

BUFx2_ASAP7_75t_L g3350 ( 
.A(n_2906),
.Y(n_3350)
);

BUFx6f_ASAP7_75t_L g3351 ( 
.A(n_2844),
.Y(n_3351)
);

OR2x2_ASAP7_75t_L g3352 ( 
.A(n_2760),
.B(n_1616),
.Y(n_3352)
);

AND2x2_ASAP7_75t_L g3353 ( 
.A(n_2741),
.B(n_1618),
.Y(n_3353)
);

INVx1_ASAP7_75t_SL g3354 ( 
.A(n_2691),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_2549),
.B(n_2488),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_2586),
.Y(n_3356)
);

INVx4_ASAP7_75t_L g3357 ( 
.A(n_2850),
.Y(n_3357)
);

BUFx4_ASAP7_75t_L g3358 ( 
.A(n_2570),
.Y(n_3358)
);

INVx5_ASAP7_75t_L g3359 ( 
.A(n_2850),
.Y(n_3359)
);

BUFx6f_ASAP7_75t_L g3360 ( 
.A(n_2850),
.Y(n_3360)
);

INVx3_ASAP7_75t_L g3361 ( 
.A(n_2742),
.Y(n_3361)
);

BUFx6f_ASAP7_75t_L g3362 ( 
.A(n_2850),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2588),
.Y(n_3363)
);

INVx2_ASAP7_75t_SL g3364 ( 
.A(n_2928),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2606),
.Y(n_3365)
);

BUFx4_ASAP7_75t_L g3366 ( 
.A(n_2737),
.Y(n_3366)
);

AND2x6_ASAP7_75t_L g3367 ( 
.A(n_2879),
.B(n_2324),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_2549),
.B(n_2489),
.Y(n_3368)
);

AND2x6_ASAP7_75t_L g3369 ( 
.A(n_2881),
.B(n_2326),
.Y(n_3369)
);

OAI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_2899),
.A2(n_2905),
.B1(n_2902),
.B2(n_2765),
.Y(n_3370)
);

INVx3_ASAP7_75t_L g3371 ( 
.A(n_2742),
.Y(n_3371)
);

BUFx2_ASAP7_75t_L g3372 ( 
.A(n_2750),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2939),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_2939),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_2550),
.B(n_2497),
.Y(n_3375)
);

INVx4_ASAP7_75t_L g3376 ( 
.A(n_2886),
.Y(n_3376)
);

BUFx2_ASAP7_75t_L g3377 ( 
.A(n_2750),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_2650),
.B(n_1881),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_2743),
.B(n_1619),
.Y(n_3379)
);

BUFx6f_ASAP7_75t_L g3380 ( 
.A(n_2886),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_2550),
.B(n_2501),
.Y(n_3381)
);

BUFx3_ASAP7_75t_L g3382 ( 
.A(n_2737),
.Y(n_3382)
);

AND2x4_ASAP7_75t_L g3383 ( 
.A(n_2942),
.B(n_1622),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_2944),
.Y(n_3384)
);

AO22x2_ASAP7_75t_L g3385 ( 
.A1(n_2794),
.A2(n_1624),
.B1(n_1626),
.B2(n_1625),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_L g3386 ( 
.A(n_2607),
.B(n_1831),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2555),
.B(n_2505),
.Y(n_3387)
);

INVx3_ASAP7_75t_L g3388 ( 
.A(n_2758),
.Y(n_3388)
);

INVx1_ASAP7_75t_SL g3389 ( 
.A(n_2691),
.Y(n_3389)
);

CKINVDCx5p33_ASAP7_75t_R g3390 ( 
.A(n_2697),
.Y(n_3390)
);

NAND2x1p5_ASAP7_75t_L g3391 ( 
.A(n_2674),
.B(n_2535),
.Y(n_3391)
);

OR2x2_ASAP7_75t_L g3392 ( 
.A(n_2786),
.B(n_1627),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2608),
.Y(n_3393)
);

OAI21xp33_ASAP7_75t_SL g3394 ( 
.A1(n_2821),
.A2(n_2126),
.B(n_1631),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_2611),
.Y(n_3395)
);

INVx8_ASAP7_75t_L g3396 ( 
.A(n_2933),
.Y(n_3396)
);

CKINVDCx5p33_ASAP7_75t_R g3397 ( 
.A(n_2556),
.Y(n_3397)
);

BUFx2_ASAP7_75t_L g3398 ( 
.A(n_2750),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_2944),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2555),
.B(n_2508),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_2945),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2945),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_SL g3403 ( 
.A(n_2902),
.B(n_2525),
.Y(n_3403)
);

BUFx6f_ASAP7_75t_L g3404 ( 
.A(n_2886),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_2612),
.Y(n_3405)
);

INVx2_ASAP7_75t_SL g3406 ( 
.A(n_2936),
.Y(n_3406)
);

INVx2_ASAP7_75t_SL g3407 ( 
.A(n_2936),
.Y(n_3407)
);

HB1xp67_ASAP7_75t_L g3408 ( 
.A(n_2938),
.Y(n_3408)
);

INVx1_ASAP7_75t_SL g3409 ( 
.A(n_2746),
.Y(n_3409)
);

BUFx2_ASAP7_75t_L g3410 ( 
.A(n_2647),
.Y(n_3410)
);

INVx4_ASAP7_75t_L g3411 ( 
.A(n_2886),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_2607),
.B(n_1835),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2618),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_2619),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_2951),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2620),
.Y(n_3416)
);

BUFx3_ASAP7_75t_L g3417 ( 
.A(n_2819),
.Y(n_3417)
);

BUFx8_ASAP7_75t_SL g3418 ( 
.A(n_2870),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_2951),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_SL g3420 ( 
.A(n_2905),
.B(n_2525),
.Y(n_3420)
);

BUFx10_ASAP7_75t_L g3421 ( 
.A(n_2701),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_2960),
.Y(n_3422)
);

INVx5_ASAP7_75t_L g3423 ( 
.A(n_2948),
.Y(n_3423)
);

BUFx2_ASAP7_75t_L g3424 ( 
.A(n_2647),
.Y(n_3424)
);

NOR2xp33_ASAP7_75t_L g3425 ( 
.A(n_2634),
.B(n_2331),
.Y(n_3425)
);

INVx2_ASAP7_75t_SL g3426 ( 
.A(n_3109),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3303),
.B(n_2622),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3276),
.B(n_2625),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3015),
.B(n_2746),
.Y(n_3429)
);

AOI22xp5_ASAP7_75t_L g3430 ( 
.A1(n_3010),
.A2(n_2735),
.B1(n_2687),
.B2(n_2634),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3304),
.Y(n_3431)
);

AND2x2_ASAP7_75t_SL g3432 ( 
.A(n_3248),
.B(n_2789),
.Y(n_3432)
);

NAND2xp33_ASAP7_75t_L g3433 ( 
.A(n_2986),
.B(n_2891),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_3342),
.B(n_2794),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3306),
.Y(n_3435)
);

NOR3xp33_ASAP7_75t_L g3436 ( 
.A(n_3142),
.B(n_2677),
.C(n_2725),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3293),
.B(n_2633),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_SL g3438 ( 
.A(n_3222),
.B(n_2907),
.Y(n_3438)
);

AND2x4_ASAP7_75t_SL g3439 ( 
.A(n_3153),
.B(n_2683),
.Y(n_3439)
);

NOR2xp33_ASAP7_75t_L g3440 ( 
.A(n_3026),
.B(n_2735),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3308),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3188),
.B(n_2559),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3156),
.B(n_2977),
.Y(n_3443)
);

INVx2_ASAP7_75t_L g3444 ( 
.A(n_3311),
.Y(n_3444)
);

O2A1O1Ixp33_ASAP7_75t_L g3445 ( 
.A1(n_3055),
.A2(n_2677),
.B(n_2725),
.C(n_2863),
.Y(n_3445)
);

OAI21xp33_ASAP7_75t_L g3446 ( 
.A1(n_3074),
.A2(n_2872),
.B(n_2861),
.Y(n_3446)
);

AO22x1_ASAP7_75t_L g3447 ( 
.A1(n_3101),
.A2(n_3102),
.B1(n_3041),
.B2(n_3057),
.Y(n_3447)
);

AND2x4_ASAP7_75t_L g3448 ( 
.A(n_2995),
.B(n_2943),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_3148),
.B(n_2924),
.Y(n_3449)
);

AOI22xp33_ASAP7_75t_L g3450 ( 
.A1(n_3055),
.A2(n_2981),
.B1(n_2950),
.B2(n_2959),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_SL g3451 ( 
.A(n_3222),
.B(n_2710),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3313),
.Y(n_3452)
);

INVx2_ASAP7_75t_SL g3453 ( 
.A(n_2991),
.Y(n_3453)
);

INVx2_ASAP7_75t_SL g3454 ( 
.A(n_3018),
.Y(n_3454)
);

INVx2_ASAP7_75t_SL g3455 ( 
.A(n_3073),
.Y(n_3455)
);

OAI221xp5_ASAP7_75t_L g3456 ( 
.A1(n_3011),
.A2(n_2854),
.B1(n_2836),
.B2(n_2686),
.C(n_2695),
.Y(n_3456)
);

NOR2xp33_ASAP7_75t_L g3457 ( 
.A(n_3119),
.B(n_2872),
.Y(n_3457)
);

INVx3_ASAP7_75t_L g3458 ( 
.A(n_3005),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3353),
.B(n_2679),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3370),
.A2(n_2966),
.B1(n_2961),
.B2(n_2962),
.Y(n_3460)
);

OAI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3370),
.A2(n_2765),
.B1(n_2894),
.B2(n_2883),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_3249),
.B(n_2692),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3118),
.B(n_2878),
.Y(n_3463)
);

AND2x4_ASAP7_75t_L g3464 ( 
.A(n_2995),
.B(n_2947),
.Y(n_3464)
);

AOI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3328),
.A2(n_2821),
.B(n_2883),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3379),
.B(n_2984),
.Y(n_3466)
);

AND2x2_ASAP7_75t_L g3467 ( 
.A(n_3194),
.B(n_2985),
.Y(n_3467)
);

AND2x6_ASAP7_75t_SL g3468 ( 
.A(n_3386),
.B(n_2647),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_3339),
.Y(n_3469)
);

INVx2_ASAP7_75t_SL g3470 ( 
.A(n_3133),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3257),
.B(n_2702),
.Y(n_3471)
);

AOI22xp5_ASAP7_75t_L g3472 ( 
.A1(n_3107),
.A2(n_2954),
.B1(n_2878),
.B2(n_2927),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3105),
.B(n_2888),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3349),
.Y(n_3474)
);

AO22x1_ASAP7_75t_L g3475 ( 
.A1(n_3305),
.A2(n_3023),
.B1(n_3214),
.B2(n_3204),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_SL g3476 ( 
.A(n_3249),
.B(n_2713),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3118),
.B(n_2888),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3270),
.B(n_2736),
.Y(n_3478)
);

AOI22xp33_ASAP7_75t_L g3479 ( 
.A1(n_3108),
.A2(n_2768),
.B1(n_2778),
.B2(n_2769),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_SL g3480 ( 
.A(n_3203),
.B(n_2791),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_2987),
.B(n_2807),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3373),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_SL g3483 ( 
.A(n_3155),
.B(n_3023),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_2987),
.B(n_2809),
.Y(n_3484)
);

INVx2_ASAP7_75t_SL g3485 ( 
.A(n_3149),
.Y(n_3485)
);

AOI22xp5_ASAP7_75t_L g3486 ( 
.A1(n_3409),
.A2(n_2930),
.B1(n_2931),
.B2(n_2927),
.Y(n_3486)
);

A2O1A1Ixp33_ASAP7_75t_L g3487 ( 
.A1(n_3161),
.A2(n_2894),
.B(n_2909),
.C(n_2931),
.Y(n_3487)
);

OAI221xp5_ASAP7_75t_L g3488 ( 
.A1(n_3136),
.A2(n_2854),
.B1(n_2838),
.B2(n_2849),
.C(n_2835),
.Y(n_3488)
);

AOI21xp5_ASAP7_75t_L g3489 ( 
.A1(n_3033),
.A2(n_2909),
.B(n_2912),
.Y(n_3489)
);

AOI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3409),
.A2(n_2930),
.B1(n_2938),
.B2(n_2756),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_3374),
.Y(n_3491)
);

CKINVDCx5p33_ASAP7_75t_R g3492 ( 
.A(n_3326),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3188),
.B(n_2830),
.Y(n_3493)
);

AOI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3145),
.A2(n_2857),
.B1(n_2860),
.B2(n_2852),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_SL g3495 ( 
.A(n_3155),
.B(n_2869),
.Y(n_3495)
);

O2A1O1Ixp33_ASAP7_75t_L g3496 ( 
.A1(n_3322),
.A2(n_2863),
.B(n_2882),
.C(n_2877),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3193),
.B(n_2913),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3193),
.B(n_3319),
.Y(n_3498)
);

AOI22xp33_ASAP7_75t_L g3499 ( 
.A1(n_3108),
.A2(n_2921),
.B1(n_2918),
.B2(n_2892),
.Y(n_3499)
);

AOI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3016),
.A2(n_2897),
.B1(n_2903),
.B2(n_2890),
.Y(n_3500)
);

AOI22xp33_ASAP7_75t_L g3501 ( 
.A1(n_3338),
.A2(n_2908),
.B1(n_2900),
.B2(n_2795),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3316),
.Y(n_3502)
);

BUFx12f_ASAP7_75t_L g3503 ( 
.A(n_3138),
.Y(n_3503)
);

BUFx3_ASAP7_75t_L g3504 ( 
.A(n_3028),
.Y(n_3504)
);

BUFx6f_ASAP7_75t_L g3505 ( 
.A(n_3065),
.Y(n_3505)
);

OR2x6_ASAP7_75t_L g3506 ( 
.A(n_2996),
.B(n_2819),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3340),
.B(n_2782),
.Y(n_3507)
);

INVx5_ASAP7_75t_L g3508 ( 
.A(n_3005),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3319),
.B(n_2749),
.Y(n_3509)
);

NOR2xp67_ASAP7_75t_L g3510 ( 
.A(n_3330),
.B(n_2796),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3113),
.B(n_2749),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3056),
.B(n_2782),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3384),
.Y(n_3513)
);

BUFx6f_ASAP7_75t_L g3514 ( 
.A(n_3065),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_SL g3515 ( 
.A(n_2993),
.B(n_2917),
.Y(n_3515)
);

AOI22xp33_ASAP7_75t_L g3516 ( 
.A1(n_3287),
.A2(n_2900),
.B1(n_2795),
.B2(n_2848),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_SL g3517 ( 
.A1(n_3136),
.A2(n_2567),
.B1(n_2843),
.B2(n_2840),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3399),
.Y(n_3518)
);

OAI22xp5_ASAP7_75t_L g3519 ( 
.A1(n_3309),
.A2(n_2592),
.B1(n_2559),
.B2(n_2782),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3071),
.B(n_3020),
.Y(n_3520)
);

O2A1O1Ixp5_ASAP7_75t_L g3521 ( 
.A1(n_3197),
.A2(n_2923),
.B(n_2597),
.C(n_2914),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3401),
.Y(n_3522)
);

INVx2_ASAP7_75t_SL g3523 ( 
.A(n_3063),
.Y(n_3523)
);

OR2x2_ASAP7_75t_L g3524 ( 
.A(n_3116),
.B(n_2637),
.Y(n_3524)
);

NAND2xp33_ASAP7_75t_L g3525 ( 
.A(n_2986),
.B(n_2795),
.Y(n_3525)
);

OAI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_3309),
.A2(n_2858),
.B(n_2592),
.Y(n_3526)
);

NOR2xp67_ASAP7_75t_L g3527 ( 
.A(n_3397),
.B(n_2874),
.Y(n_3527)
);

A2O1A1Ixp33_ASAP7_75t_L g3528 ( 
.A1(n_3425),
.A2(n_2919),
.B(n_2865),
.C(n_2887),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_3402),
.Y(n_3529)
);

HB1xp67_ASAP7_75t_L g3530 ( 
.A(n_3054),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3113),
.B(n_2795),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3062),
.B(n_2795),
.Y(n_3532)
);

NOR3xp33_ASAP7_75t_L g3533 ( 
.A(n_3335),
.B(n_2925),
.C(n_2920),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_SL g3534 ( 
.A(n_2993),
.B(n_2948),
.Y(n_3534)
);

INVx3_ASAP7_75t_L g3535 ( 
.A(n_3005),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_2999),
.B(n_2562),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_2999),
.B(n_3062),
.Y(n_3537)
);

OR2x2_ASAP7_75t_L g3538 ( 
.A(n_3058),
.B(n_2637),
.Y(n_3538)
);

NOR2xp33_ASAP7_75t_L g3539 ( 
.A(n_3104),
.B(n_2701),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3081),
.B(n_2757),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3329),
.B(n_2565),
.Y(n_3541)
);

AND2x2_ASAP7_75t_L g3542 ( 
.A(n_3096),
.B(n_2637),
.Y(n_3542)
);

OAI22xp5_ASAP7_75t_L g3543 ( 
.A1(n_3013),
.A2(n_2963),
.B1(n_2965),
.B2(n_2960),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3177),
.B(n_2819),
.Y(n_3544)
);

AOI22xp5_ASAP7_75t_L g3545 ( 
.A1(n_3013),
.A2(n_2848),
.B1(n_2929),
.B2(n_2920),
.Y(n_3545)
);

AOI22xp33_ASAP7_75t_L g3546 ( 
.A1(n_3287),
.A2(n_2848),
.B1(n_2911),
.B2(n_2864),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3352),
.B(n_3317),
.Y(n_3547)
);

AOI22xp5_ASAP7_75t_L g3548 ( 
.A1(n_3006),
.A2(n_2848),
.B1(n_2929),
.B2(n_2831),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3321),
.B(n_2848),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3415),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3341),
.B(n_2569),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3344),
.B(n_2609),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3345),
.B(n_2614),
.Y(n_3553)
);

A2O1A1Ixp33_ASAP7_75t_L g3554 ( 
.A1(n_3154),
.A2(n_2628),
.B(n_2965),
.C(n_2963),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_3346),
.Y(n_3555)
);

AOI22xp5_ASAP7_75t_L g3556 ( 
.A1(n_3006),
.A2(n_3012),
.B1(n_3053),
.B2(n_3364),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_3419),
.Y(n_3557)
);

INVx2_ASAP7_75t_SL g3558 ( 
.A(n_3110),
.Y(n_3558)
);

CKINVDCx5p33_ASAP7_75t_R g3559 ( 
.A(n_3158),
.Y(n_3559)
);

OAI22xp5_ASAP7_75t_SL g3560 ( 
.A1(n_3121),
.A2(n_1148),
.B1(n_1162),
.B2(n_861),
.Y(n_3560)
);

CKINVDCx5p33_ASAP7_75t_R g3561 ( 
.A(n_3390),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3356),
.B(n_2967),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_SL g3563 ( 
.A(n_3153),
.B(n_2948),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_SL g3564 ( 
.A(n_3004),
.B(n_2948),
.Y(n_3564)
);

BUFx8_ASAP7_75t_L g3565 ( 
.A(n_3098),
.Y(n_3565)
);

CKINVDCx20_ASAP7_75t_R g3566 ( 
.A(n_3076),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3363),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3365),
.B(n_3393),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3395),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3405),
.Y(n_3570)
);

INVx4_ASAP7_75t_L g3571 ( 
.A(n_3049),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3413),
.Y(n_3572)
);

AND2x4_ASAP7_75t_SL g3573 ( 
.A(n_3157),
.B(n_2739),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3331),
.A2(n_2967),
.B1(n_2971),
.B2(n_2970),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3414),
.Y(n_3575)
);

OAI22xp5_ASAP7_75t_L g3576 ( 
.A1(n_3279),
.A2(n_2971),
.B1(n_2975),
.B2(n_2970),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3416),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_2983),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3115),
.B(n_1628),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3114),
.B(n_2975),
.Y(n_3580)
);

AND2x2_ASAP7_75t_SL g3581 ( 
.A(n_3196),
.B(n_2397),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3114),
.B(n_2758),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3061),
.B(n_2764),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_2990),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_SL g3585 ( 
.A(n_3004),
.B(n_2739),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3061),
.B(n_2764),
.Y(n_3586)
);

BUFx3_ASAP7_75t_L g3587 ( 
.A(n_3094),
.Y(n_3587)
);

A2O1A1Ixp33_ASAP7_75t_L g3588 ( 
.A1(n_3154),
.A2(n_2788),
.B(n_2829),
.C(n_2785),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3046),
.B(n_2785),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_SL g3590 ( 
.A(n_3012),
.B(n_2876),
.Y(n_3590)
);

AOI22xp5_ASAP7_75t_L g3591 ( 
.A1(n_3296),
.A2(n_2831),
.B1(n_2953),
.B2(n_2949),
.Y(n_3591)
);

INVx2_ASAP7_75t_SL g3592 ( 
.A(n_3180),
.Y(n_3592)
);

BUFx3_ASAP7_75t_L g3593 ( 
.A(n_2996),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3331),
.B(n_3088),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3354),
.B(n_2788),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_2998),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3001),
.Y(n_3597)
);

INVx2_ASAP7_75t_SL g3598 ( 
.A(n_3305),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3422),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_2989),
.Y(n_3600)
);

AOI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_3272),
.A2(n_2953),
.B1(n_2956),
.B2(n_2949),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_3322),
.B(n_2876),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3070),
.B(n_2986),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3088),
.B(n_2829),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_SL g3605 ( 
.A(n_3354),
.B(n_2893),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3165),
.B(n_2832),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3070),
.B(n_2832),
.Y(n_3607)
);

AND2x6_ASAP7_75t_L g3608 ( 
.A(n_3049),
.B(n_2922),
.Y(n_3608)
);

AOI22xp33_ASAP7_75t_L g3609 ( 
.A1(n_3272),
.A2(n_2958),
.B1(n_2974),
.B2(n_2956),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_SL g3610 ( 
.A(n_3389),
.B(n_2893),
.Y(n_3610)
);

BUFx3_ASAP7_75t_L g3611 ( 
.A(n_2996),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3212),
.B(n_3190),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3002),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3003),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3007),
.Y(n_3615)
);

NOR2xp33_ASAP7_75t_L g3616 ( 
.A(n_3389),
.B(n_2851),
.Y(n_3616)
);

AO22x1_ASAP7_75t_L g3617 ( 
.A1(n_3343),
.A2(n_2099),
.B1(n_2053),
.B2(n_844),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_SL g3618 ( 
.A(n_3049),
.B(n_2896),
.Y(n_3618)
);

AOI22xp5_ASAP7_75t_L g3619 ( 
.A1(n_3315),
.A2(n_2974),
.B1(n_2958),
.B2(n_2880),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_3218),
.B(n_3392),
.Y(n_3620)
);

AOI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_2986),
.A2(n_2926),
.B1(n_2910),
.B2(n_2880),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3009),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_L g3623 ( 
.A(n_3078),
.B(n_2851),
.Y(n_3623)
);

INVx3_ASAP7_75t_L g3624 ( 
.A(n_3051),
.Y(n_3624)
);

OR2x2_ASAP7_75t_L g3625 ( 
.A(n_3075),
.B(n_2935),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_3033),
.A2(n_2896),
.B(n_2904),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3024),
.Y(n_3627)
);

OR2x2_ASAP7_75t_L g3628 ( 
.A(n_3100),
.B(n_2937),
.Y(n_3628)
);

OR2x6_ASAP7_75t_L g3629 ( 
.A(n_3396),
.B(n_3243),
.Y(n_3629)
);

AOI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3348),
.A2(n_2926),
.B1(n_2910),
.B2(n_2823),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3160),
.B(n_2904),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3029),
.Y(n_3632)
);

AOI22xp33_ASAP7_75t_L g3633 ( 
.A1(n_3348),
.A2(n_2823),
.B1(n_2806),
.B2(n_2969),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3175),
.B(n_2915),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3185),
.B(n_2915),
.Y(n_3635)
);

AOI22xp5_ASAP7_75t_L g3636 ( 
.A1(n_3220),
.A2(n_3111),
.B1(n_3095),
.B2(n_3279),
.Y(n_3636)
);

BUFx2_ASAP7_75t_L g3637 ( 
.A(n_3223),
.Y(n_3637)
);

O2A1O1Ixp33_ASAP7_75t_L g3638 ( 
.A1(n_3259),
.A2(n_2806),
.B(n_2973),
.C(n_2972),
.Y(n_3638)
);

INVx2_ASAP7_75t_SL g3639 ( 
.A(n_3255),
.Y(n_3639)
);

BUFx3_ASAP7_75t_L g3640 ( 
.A(n_3396),
.Y(n_3640)
);

INVx3_ASAP7_75t_L g3641 ( 
.A(n_3051),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3233),
.B(n_3210),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3233),
.B(n_2979),
.Y(n_3643)
);

OAI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_3068),
.A2(n_845),
.B1(n_848),
.B2(n_841),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3233),
.B(n_2982),
.Y(n_3645)
);

INVx3_ASAP7_75t_L g3646 ( 
.A(n_3051),
.Y(n_3646)
);

NAND3xp33_ASAP7_75t_SL g3647 ( 
.A(n_3378),
.B(n_849),
.C(n_848),
.Y(n_3647)
);

BUFx3_ASAP7_75t_L g3648 ( 
.A(n_3396),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_3065),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3233),
.B(n_2511),
.Y(n_3650)
);

AOI22xp33_ASAP7_75t_L g3651 ( 
.A1(n_3383),
.A2(n_2517),
.B1(n_2518),
.B2(n_2516),
.Y(n_3651)
);

AOI22xp5_ASAP7_75t_L g3652 ( 
.A1(n_3220),
.A2(n_2534),
.B1(n_2536),
.B2(n_2521),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3210),
.B(n_2538),
.Y(n_3653)
);

INVx3_ASAP7_75t_L g3654 ( 
.A(n_2997),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_3235),
.B(n_1633),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3291),
.B(n_1635),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3254),
.B(n_2545),
.Y(n_3657)
);

INVx1_ASAP7_75t_L g3658 ( 
.A(n_3036),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_SL g3659 ( 
.A(n_3078),
.B(n_2797),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_SL g3660 ( 
.A(n_3123),
.B(n_2797),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3123),
.B(n_983),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3254),
.B(n_2332),
.Y(n_3662)
);

NOR2xp33_ASAP7_75t_L g3663 ( 
.A(n_3292),
.B(n_984),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3262),
.B(n_2334),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_SL g3665 ( 
.A(n_3213),
.B(n_2797),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3044),
.Y(n_3666)
);

INVx2_ASAP7_75t_SL g3667 ( 
.A(n_3266),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3176),
.B(n_2336),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3017),
.B(n_2338),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3021),
.Y(n_3670)
);

BUFx2_ASAP7_75t_L g3671 ( 
.A(n_3297),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3245),
.B(n_2342),
.Y(n_3672)
);

BUFx3_ASAP7_75t_L g3673 ( 
.A(n_3382),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_SL g3674 ( 
.A(n_3213),
.B(n_2797),
.Y(n_3674)
);

NOR2xp33_ASAP7_75t_L g3675 ( 
.A(n_3216),
.B(n_987),
.Y(n_3675)
);

BUFx6f_ASAP7_75t_L g3676 ( 
.A(n_3067),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_SL g3677 ( 
.A(n_3213),
.B(n_2895),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3245),
.B(n_3253),
.Y(n_3678)
);

OAI21xp5_ASAP7_75t_L g3679 ( 
.A1(n_3394),
.A2(n_2356),
.B(n_2350),
.Y(n_3679)
);

INVx3_ASAP7_75t_L g3680 ( 
.A(n_2997),
.Y(n_3680)
);

AOI22xp5_ASAP7_75t_SL g3681 ( 
.A1(n_3281),
.A2(n_850),
.B1(n_861),
.B2(n_849),
.Y(n_3681)
);

NOR3xp33_ASAP7_75t_SL g3682 ( 
.A(n_3282),
.B(n_1008),
.C(n_850),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3253),
.B(n_2359),
.Y(n_3683)
);

HB1xp67_ASAP7_75t_L g3684 ( 
.A(n_3307),
.Y(n_3684)
);

BUFx6f_ASAP7_75t_L g3685 ( 
.A(n_3067),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3262),
.B(n_2361),
.Y(n_3686)
);

INVx2_ASAP7_75t_SL g3687 ( 
.A(n_3327),
.Y(n_3687)
);

NAND3xp33_ASAP7_75t_SL g3688 ( 
.A(n_3196),
.B(n_1010),
.C(n_1008),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3200),
.B(n_989),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3035),
.Y(n_3690)
);

AND2x6_ASAP7_75t_L g3691 ( 
.A(n_3014),
.B(n_2362),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3030),
.B(n_2363),
.Y(n_3692)
);

INVx8_ASAP7_75t_L g3693 ( 
.A(n_2988),
.Y(n_3693)
);

AOI22xp33_ASAP7_75t_L g3694 ( 
.A1(n_3383),
.A2(n_2366),
.B1(n_2364),
.B2(n_1999),
.Y(n_3694)
);

NAND2x1p5_ASAP7_75t_L g3695 ( 
.A(n_3008),
.B(n_2895),
.Y(n_3695)
);

AND3x1_ASAP7_75t_L g3696 ( 
.A(n_3333),
.B(n_1637),
.C(n_1636),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3030),
.B(n_2236),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3043),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3032),
.B(n_2236),
.Y(n_3699)
);

INVxp67_ASAP7_75t_SL g3700 ( 
.A(n_3067),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3069),
.Y(n_3701)
);

NOR2xp33_ASAP7_75t_L g3702 ( 
.A(n_3350),
.B(n_990),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3334),
.B(n_3178),
.Y(n_3703)
);

OR2x6_ASAP7_75t_L g3704 ( 
.A(n_3243),
.B(n_1641),
.Y(n_3704)
);

INVxp67_ASAP7_75t_SL g3705 ( 
.A(n_3093),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3045),
.Y(n_3706)
);

INVxp33_ASAP7_75t_L g3707 ( 
.A(n_3408),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3146),
.Y(n_3708)
);

INVxp67_ASAP7_75t_L g3709 ( 
.A(n_3385),
.Y(n_3709)
);

NAND2x1_ASAP7_75t_L g3710 ( 
.A(n_2988),
.B(n_2236),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3047),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3048),
.Y(n_3712)
);

INVx3_ASAP7_75t_L g3713 ( 
.A(n_3008),
.Y(n_3713)
);

OR2x6_ASAP7_75t_L g3714 ( 
.A(n_3243),
.B(n_1642),
.Y(n_3714)
);

INVx2_ASAP7_75t_L g3715 ( 
.A(n_3151),
.Y(n_3715)
);

NOR2xp33_ASAP7_75t_SL g3716 ( 
.A(n_3237),
.B(n_2053),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3178),
.B(n_2261),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3077),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3083),
.Y(n_3719)
);

NOR3xp33_ASAP7_75t_SL g3720 ( 
.A(n_3412),
.B(n_1011),
.C(n_1010),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3084),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_3286),
.B(n_2895),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_3347),
.B(n_992),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3086),
.Y(n_3724)
);

HB1xp67_ASAP7_75t_L g3725 ( 
.A(n_3246),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3163),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3087),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3032),
.B(n_2261),
.Y(n_3728)
);

INVx8_ASAP7_75t_L g3729 ( 
.A(n_2988),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3037),
.B(n_2261),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3168),
.Y(n_3731)
);

NOR2x2_ASAP7_75t_L g3732 ( 
.A(n_3042),
.B(n_1441),
.Y(n_3732)
);

AND2x6_ASAP7_75t_SL g3733 ( 
.A(n_3042),
.B(n_1645),
.Y(n_3733)
);

O2A1O1Ixp5_ASAP7_75t_L g3734 ( 
.A1(n_3103),
.A2(n_2323),
.B(n_2341),
.C(n_2315),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3037),
.B(n_2315),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_SL g3736 ( 
.A(n_3286),
.B(n_2895),
.Y(n_3736)
);

NOR2xp33_ASAP7_75t_L g3737 ( 
.A(n_3242),
.B(n_994),
.Y(n_3737)
);

NOR2xp67_ASAP7_75t_SL g3738 ( 
.A(n_3068),
.B(n_2978),
.Y(n_3738)
);

NOR2xp33_ASAP7_75t_L g3739 ( 
.A(n_3250),
.B(n_998),
.Y(n_3739)
);

NAND3xp33_ASAP7_75t_L g3740 ( 
.A(n_3025),
.B(n_3172),
.C(n_3198),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3050),
.B(n_2315),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3090),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3050),
.B(n_2323),
.Y(n_3743)
);

AOI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3095),
.A2(n_2177),
.B1(n_2178),
.B2(n_2144),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_SL g3745 ( 
.A(n_3286),
.B(n_2978),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3082),
.B(n_2323),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3082),
.B(n_2341),
.Y(n_3747)
);

NOR2xp33_ASAP7_75t_L g3748 ( 
.A(n_3128),
.B(n_1002),
.Y(n_3748)
);

AOI22xp33_ASAP7_75t_L g3749 ( 
.A1(n_3291),
.A2(n_1999),
.B1(n_2002),
.B2(n_1996),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3225),
.B(n_2341),
.Y(n_3750)
);

CKINVDCx5p33_ASAP7_75t_R g3751 ( 
.A(n_3418),
.Y(n_3751)
);

HB1xp67_ASAP7_75t_L g3752 ( 
.A(n_3246),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3092),
.Y(n_3753)
);

A2O1A1Ixp33_ASAP7_75t_L g3754 ( 
.A1(n_3025),
.A2(n_1648),
.B(n_1649),
.C(n_1647),
.Y(n_3754)
);

AND2x2_ASAP7_75t_L g3755 ( 
.A(n_3298),
.B(n_1653),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_3225),
.B(n_2351),
.Y(n_3756)
);

NOR2xp33_ASAP7_75t_L g3757 ( 
.A(n_3298),
.B(n_1004),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3314),
.B(n_3324),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3106),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_SL g3760 ( 
.A(n_3359),
.B(n_2978),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3314),
.B(n_2351),
.Y(n_3761)
);

OAI221xp5_ASAP7_75t_L g3762 ( 
.A1(n_3406),
.A2(n_1012),
.B1(n_1148),
.B2(n_1144),
.C(n_1011),
.Y(n_3762)
);

INVx3_ASAP7_75t_L g3763 ( 
.A(n_3034),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3324),
.B(n_2351),
.Y(n_3764)
);

NOR2xp33_ASAP7_75t_L g3765 ( 
.A(n_3407),
.B(n_1005),
.Y(n_3765)
);

NOR2xp33_ASAP7_75t_SL g3766 ( 
.A(n_3237),
.B(n_2099),
.Y(n_3766)
);

BUFx6f_ASAP7_75t_L g3767 ( 
.A(n_3093),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3183),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3192),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3111),
.B(n_2352),
.Y(n_3770)
);

AOI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3323),
.A2(n_2177),
.B1(n_2178),
.B2(n_2144),
.Y(n_3771)
);

NOR2x1p5_ASAP7_75t_L g3772 ( 
.A(n_3417),
.B(n_1012),
.Y(n_3772)
);

INVx8_ASAP7_75t_L g3773 ( 
.A(n_2988),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3112),
.B(n_2352),
.Y(n_3774)
);

AOI22xp33_ASAP7_75t_L g3775 ( 
.A1(n_3403),
.A2(n_3420),
.B1(n_3201),
.B2(n_3206),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3195),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_L g3777 ( 
.A(n_3034),
.B(n_1023),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_SL g3778 ( 
.A(n_3359),
.B(n_2978),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3122),
.B(n_2352),
.Y(n_3779)
);

NOR3xp33_ASAP7_75t_SL g3780 ( 
.A(n_3019),
.B(n_1149),
.C(n_1144),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3215),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3226),
.Y(n_3782)
);

BUFx6f_ASAP7_75t_SL g3783 ( 
.A(n_3042),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3131),
.B(n_2390),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3134),
.B(n_2390),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3135),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3137),
.B(n_2390),
.Y(n_3787)
);

INVx1_ASAP7_75t_SL g3788 ( 
.A(n_3366),
.Y(n_3788)
);

CKINVDCx5p33_ASAP7_75t_R g3789 ( 
.A(n_3098),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3139),
.Y(n_3790)
);

NAND2xp33_ASAP7_75t_L g3791 ( 
.A(n_3040),
.B(n_3068),
.Y(n_3791)
);

AOI22xp33_ASAP7_75t_L g3792 ( 
.A1(n_3205),
.A2(n_1999),
.B1(n_2002),
.B2(n_1996),
.Y(n_3792)
);

INVxp67_ASAP7_75t_L g3793 ( 
.A(n_3385),
.Y(n_3793)
);

OR2x2_ASAP7_75t_L g3794 ( 
.A(n_3208),
.B(n_1656),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3140),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3231),
.Y(n_3796)
);

AOI22xp33_ASAP7_75t_L g3797 ( 
.A1(n_3209),
.A2(n_1999),
.B1(n_2002),
.B2(n_1996),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3232),
.Y(n_3798)
);

BUFx6f_ASAP7_75t_L g3799 ( 
.A(n_3093),
.Y(n_3799)
);

INVx2_ASAP7_75t_SL g3800 ( 
.A(n_3421),
.Y(n_3800)
);

INVx5_ASAP7_75t_L g3801 ( 
.A(n_3040),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_SL g3802 ( 
.A(n_3359),
.B(n_2535),
.Y(n_3802)
);

AOI22xp33_ASAP7_75t_L g3803 ( 
.A1(n_3302),
.A2(n_2002),
.B1(n_2017),
.B2(n_1996),
.Y(n_3803)
);

AOI221xp5_ASAP7_75t_L g3804 ( 
.A1(n_3031),
.A2(n_1152),
.B1(n_1153),
.B2(n_1150),
.C(n_1149),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3239),
.Y(n_3805)
);

BUFx2_ASAP7_75t_L g3806 ( 
.A(n_3372),
.Y(n_3806)
);

CKINVDCx5p33_ASAP7_75t_R g3807 ( 
.A(n_3325),
.Y(n_3807)
);

AND2x2_ASAP7_75t_L g3808 ( 
.A(n_3019),
.B(n_1659),
.Y(n_3808)
);

INVx2_ASAP7_75t_SL g3809 ( 
.A(n_3504),
.Y(n_3809)
);

CKINVDCx20_ASAP7_75t_R g3810 ( 
.A(n_3566),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3457),
.B(n_3132),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3473),
.B(n_3312),
.Y(n_3812)
);

NOR2xp33_ASAP7_75t_R g3813 ( 
.A(n_3492),
.B(n_3236),
.Y(n_3813)
);

BUFx6f_ASAP7_75t_L g3814 ( 
.A(n_3505),
.Y(n_3814)
);

HB1xp67_ASAP7_75t_L g3815 ( 
.A(n_3598),
.Y(n_3815)
);

NOR2xp33_ASAP7_75t_L g3816 ( 
.A(n_3447),
.B(n_3421),
.Y(n_3816)
);

INVx4_ASAP7_75t_L g3817 ( 
.A(n_3508),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3452),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3502),
.Y(n_3819)
);

BUFx6f_ASAP7_75t_L g3820 ( 
.A(n_3505),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3555),
.Y(n_3821)
);

AOI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_3446),
.A2(n_3031),
.B1(n_3332),
.B2(n_3234),
.Y(n_3822)
);

AOI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3675),
.A2(n_3436),
.B1(n_3520),
.B2(n_3472),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_SL g3824 ( 
.A(n_3486),
.B(n_3038),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3466),
.B(n_3014),
.Y(n_3825)
);

O2A1O1Ixp33_ASAP7_75t_L g3826 ( 
.A1(n_3647),
.A2(n_3202),
.B(n_3227),
.C(n_3079),
.Y(n_3826)
);

INVx2_ASAP7_75t_SL g3827 ( 
.A(n_3587),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3463),
.B(n_3052),
.Y(n_3828)
);

NOR2xp33_ASAP7_75t_L g3829 ( 
.A(n_3449),
.B(n_3377),
.Y(n_3829)
);

INVx2_ASAP7_75t_SL g3830 ( 
.A(n_3673),
.Y(n_3830)
);

NOR2xp33_ASAP7_75t_L g3831 ( 
.A(n_3434),
.B(n_3398),
.Y(n_3831)
);

BUFx6f_ASAP7_75t_L g3832 ( 
.A(n_3505),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3567),
.Y(n_3833)
);

INVx2_ASAP7_75t_SL g3834 ( 
.A(n_3426),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3569),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3477),
.B(n_3052),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3570),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3467),
.B(n_3211),
.Y(n_3838)
);

INVx2_ASAP7_75t_L g3839 ( 
.A(n_3572),
.Y(n_3839)
);

NOR2xp33_ASAP7_75t_L g3840 ( 
.A(n_3620),
.B(n_3410),
.Y(n_3840)
);

OR2x2_ASAP7_75t_L g3841 ( 
.A(n_3547),
.B(n_3424),
.Y(n_3841)
);

BUFx6f_ASAP7_75t_L g3842 ( 
.A(n_3514),
.Y(n_3842)
);

INVx3_ASAP7_75t_L g3843 ( 
.A(n_3693),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3448),
.B(n_3079),
.Y(n_3844)
);

CKINVDCx5p33_ASAP7_75t_R g3845 ( 
.A(n_3561),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3575),
.Y(n_3846)
);

CKINVDCx5p33_ASAP7_75t_R g3847 ( 
.A(n_3559),
.Y(n_3847)
);

AOI22xp33_ASAP7_75t_L g3848 ( 
.A1(n_3432),
.A2(n_3332),
.B1(n_3234),
.B2(n_3217),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3428),
.B(n_3219),
.Y(n_3849)
);

AND2x2_ASAP7_75t_SL g3850 ( 
.A(n_3581),
.B(n_3038),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3437),
.B(n_3229),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3577),
.Y(n_3852)
);

CKINVDCx5p33_ASAP7_75t_R g3853 ( 
.A(n_3751),
.Y(n_3853)
);

OR2x2_ASAP7_75t_L g3854 ( 
.A(n_3612),
.B(n_3230),
.Y(n_3854)
);

AND2x4_ASAP7_75t_L g3855 ( 
.A(n_3448),
.B(n_3066),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3568),
.Y(n_3856)
);

OR2x2_ASAP7_75t_SL g3857 ( 
.A(n_3538),
.B(n_3358),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3578),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3431),
.Y(n_3859)
);

BUFx3_ASAP7_75t_L g3860 ( 
.A(n_3593),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3427),
.B(n_3247),
.Y(n_3861)
);

BUFx2_ASAP7_75t_L g3862 ( 
.A(n_3455),
.Y(n_3862)
);

AND3x2_ASAP7_75t_SL g3863 ( 
.A(n_3681),
.B(n_3260),
.C(n_3240),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3435),
.Y(n_3864)
);

BUFx3_ASAP7_75t_L g3865 ( 
.A(n_3611),
.Y(n_3865)
);

AOI22xp33_ASAP7_75t_L g3866 ( 
.A1(n_3663),
.A2(n_3251),
.B1(n_3269),
.B2(n_3263),
.Y(n_3866)
);

AND2x2_ASAP7_75t_L g3867 ( 
.A(n_3429),
.B(n_3271),
.Y(n_3867)
);

HB1xp67_ASAP7_75t_L g3868 ( 
.A(n_3530),
.Y(n_3868)
);

BUFx5_ASAP7_75t_L g3869 ( 
.A(n_3691),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_3459),
.B(n_3273),
.Y(n_3870)
);

BUFx2_ASAP7_75t_L g3871 ( 
.A(n_3637),
.Y(n_3871)
);

INVx3_ASAP7_75t_L g3872 ( 
.A(n_3693),
.Y(n_3872)
);

INVx4_ASAP7_75t_L g3873 ( 
.A(n_3508),
.Y(n_3873)
);

AND2x4_ASAP7_75t_L g3874 ( 
.A(n_3464),
.B(n_3066),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3443),
.B(n_3141),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3584),
.Y(n_3876)
);

BUFx12f_ASAP7_75t_L g3877 ( 
.A(n_3503),
.Y(n_3877)
);

INVx2_ASAP7_75t_SL g3878 ( 
.A(n_3454),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3596),
.Y(n_3879)
);

INVx4_ASAP7_75t_L g3880 ( 
.A(n_3508),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3597),
.Y(n_3881)
);

INVx5_ASAP7_75t_L g3882 ( 
.A(n_3693),
.Y(n_3882)
);

O2A1O1Ixp33_ASAP7_75t_L g3883 ( 
.A1(n_3488),
.A2(n_3277),
.B(n_3085),
.C(n_3152),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3441),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_3430),
.B(n_3039),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3613),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3614),
.Y(n_3887)
);

NOR2xp33_ASAP7_75t_R g3888 ( 
.A(n_3789),
.B(n_3295),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3481),
.B(n_3147),
.Y(n_3889)
);

BUFx3_ASAP7_75t_L g3890 ( 
.A(n_3640),
.Y(n_3890)
);

BUFx3_ASAP7_75t_L g3891 ( 
.A(n_3648),
.Y(n_3891)
);

AND2x6_ASAP7_75t_SL g3892 ( 
.A(n_3539),
.B(n_3256),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3444),
.Y(n_3893)
);

NOR2xp33_ASAP7_75t_L g3894 ( 
.A(n_3440),
.B(n_3325),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3615),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3484),
.B(n_3159),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3622),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3579),
.B(n_3171),
.Y(n_3898)
);

OR2x6_ASAP7_75t_L g3899 ( 
.A(n_3506),
.B(n_3171),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3493),
.B(n_3162),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3627),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3632),
.Y(n_3902)
);

OR2x6_ASAP7_75t_L g3903 ( 
.A(n_3506),
.B(n_3080),
.Y(n_3903)
);

BUFx3_ASAP7_75t_L g3904 ( 
.A(n_3453),
.Y(n_3904)
);

INVx4_ASAP7_75t_L g3905 ( 
.A(n_3729),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3469),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3658),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3497),
.B(n_3164),
.Y(n_3908)
);

INVxp67_ASAP7_75t_L g3909 ( 
.A(n_3483),
.Y(n_3909)
);

AOI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3542),
.A2(n_3124),
.B1(n_3166),
.B2(n_3126),
.Y(n_3910)
);

AOI22xp33_ASAP7_75t_L g3911 ( 
.A1(n_3689),
.A2(n_3124),
.B1(n_3166),
.B2(n_3126),
.Y(n_3911)
);

INVx2_ASAP7_75t_SL g3912 ( 
.A(n_3523),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3666),
.Y(n_3913)
);

BUFx3_ASAP7_75t_L g3914 ( 
.A(n_3806),
.Y(n_3914)
);

AND2x4_ASAP7_75t_L g3915 ( 
.A(n_3464),
.B(n_3080),
.Y(n_3915)
);

AND2x4_ASAP7_75t_L g3916 ( 
.A(n_3758),
.B(n_3285),
.Y(n_3916)
);

AND2x4_ASAP7_75t_L g3917 ( 
.A(n_3439),
.B(n_3285),
.Y(n_3917)
);

INVx5_ASAP7_75t_L g3918 ( 
.A(n_3729),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_3592),
.Y(n_3919)
);

AND2x4_ASAP7_75t_L g3920 ( 
.A(n_3506),
.B(n_3039),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3706),
.Y(n_3921)
);

HB1xp67_ASAP7_75t_L g3922 ( 
.A(n_3639),
.Y(n_3922)
);

OR2x2_ASAP7_75t_SL g3923 ( 
.A(n_3688),
.B(n_1661),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3474),
.Y(n_3924)
);

INVx2_ASAP7_75t_L g3925 ( 
.A(n_3482),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3711),
.Y(n_3926)
);

CKINVDCx5p33_ASAP7_75t_R g3927 ( 
.A(n_3565),
.Y(n_3927)
);

AND2x4_ASAP7_75t_L g3928 ( 
.A(n_3629),
.B(n_3059),
.Y(n_3928)
);

OAI22xp33_ASAP7_75t_L g3929 ( 
.A1(n_3716),
.A2(n_3173),
.B1(n_3182),
.B2(n_3072),
.Y(n_3929)
);

CKINVDCx20_ASAP7_75t_R g3930 ( 
.A(n_3565),
.Y(n_3930)
);

INVx4_ASAP7_75t_L g3931 ( 
.A(n_3729),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3491),
.Y(n_3932)
);

INVx5_ASAP7_75t_L g3933 ( 
.A(n_3773),
.Y(n_3933)
);

CKINVDCx8_ASAP7_75t_R g3934 ( 
.A(n_3733),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3537),
.B(n_3167),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3712),
.Y(n_3936)
);

INVx3_ASAP7_75t_L g3937 ( 
.A(n_3773),
.Y(n_3937)
);

BUFx6f_ASAP7_75t_L g3938 ( 
.A(n_3514),
.Y(n_3938)
);

BUFx3_ASAP7_75t_L g3939 ( 
.A(n_3470),
.Y(n_3939)
);

INVx4_ASAP7_75t_L g3940 ( 
.A(n_3773),
.Y(n_3940)
);

BUFx6f_ASAP7_75t_L g3941 ( 
.A(n_3514),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3537),
.B(n_3169),
.Y(n_3942)
);

CKINVDCx20_ASAP7_75t_R g3943 ( 
.A(n_3807),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3513),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3471),
.B(n_3170),
.Y(n_3945)
);

BUFx2_ASAP7_75t_L g3946 ( 
.A(n_3524),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3718),
.Y(n_3947)
);

INVx2_ASAP7_75t_SL g3948 ( 
.A(n_3485),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3518),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3522),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3529),
.Y(n_3951)
);

CKINVDCx5p33_ASAP7_75t_R g3952 ( 
.A(n_3783),
.Y(n_3952)
);

INVx4_ASAP7_75t_L g3953 ( 
.A(n_3801),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3656),
.B(n_3264),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3550),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3557),
.Y(n_3956)
);

BUFx6f_ASAP7_75t_L g3957 ( 
.A(n_3649),
.Y(n_3957)
);

BUFx6f_ASAP7_75t_L g3958 ( 
.A(n_3649),
.Y(n_3958)
);

BUFx6f_ASAP7_75t_L g3959 ( 
.A(n_3649),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3719),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3478),
.B(n_3655),
.Y(n_3961)
);

OR2x6_ASAP7_75t_L g3962 ( 
.A(n_3629),
.B(n_3059),
.Y(n_3962)
);

NAND2x1p5_ASAP7_75t_L g3963 ( 
.A(n_3801),
.B(n_3060),
.Y(n_3963)
);

BUFx6f_ASAP7_75t_L g3964 ( 
.A(n_3676),
.Y(n_3964)
);

BUFx2_ASAP7_75t_L g3965 ( 
.A(n_3558),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_SL g3966 ( 
.A(n_3494),
.B(n_3060),
.Y(n_3966)
);

INVx4_ASAP7_75t_L g3967 ( 
.A(n_3801),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3721),
.Y(n_3968)
);

BUFx2_ASAP7_75t_L g3969 ( 
.A(n_3671),
.Y(n_3969)
);

INVx5_ASAP7_75t_L g3970 ( 
.A(n_3608),
.Y(n_3970)
);

INVx2_ASAP7_75t_SL g3971 ( 
.A(n_3800),
.Y(n_3971)
);

HB1xp67_ASAP7_75t_L g3972 ( 
.A(n_3684),
.Y(n_3972)
);

NOR2xp33_ASAP7_75t_L g3973 ( 
.A(n_3475),
.B(n_3120),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3703),
.B(n_3174),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3717),
.Y(n_3975)
);

INVx2_ASAP7_75t_L g3976 ( 
.A(n_3599),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3755),
.B(n_3299),
.Y(n_3977)
);

NOR2xp33_ASAP7_75t_L g3978 ( 
.A(n_3480),
.B(n_3120),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_SL g3979 ( 
.A(n_3490),
.B(n_3072),
.Y(n_3979)
);

AOI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3507),
.A2(n_3089),
.B1(n_3187),
.B2(n_3144),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_3600),
.Y(n_3981)
);

NOR2xp33_ASAP7_75t_L g3982 ( 
.A(n_3456),
.B(n_3702),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3670),
.Y(n_3983)
);

BUFx2_ASAP7_75t_L g3984 ( 
.A(n_3709),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3724),
.Y(n_3985)
);

INVx3_ASAP7_75t_L g3986 ( 
.A(n_3654),
.Y(n_3986)
);

INVx2_ASAP7_75t_L g3987 ( 
.A(n_3690),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3727),
.Y(n_3988)
);

INVx1_ASAP7_75t_SL g3989 ( 
.A(n_3788),
.Y(n_3989)
);

AND2x4_ASAP7_75t_L g3990 ( 
.A(n_3629),
.B(n_3129),
.Y(n_3990)
);

BUFx3_ASAP7_75t_L g3991 ( 
.A(n_3725),
.Y(n_3991)
);

BUFx6f_ASAP7_75t_L g3992 ( 
.A(n_3676),
.Y(n_3992)
);

AND3x2_ASAP7_75t_SL g3993 ( 
.A(n_3681),
.B(n_3300),
.C(n_1722),
.Y(n_3993)
);

AOI221xp5_ASAP7_75t_L g3994 ( 
.A1(n_3804),
.A2(n_3445),
.B1(n_3560),
.B2(n_3762),
.C(n_3661),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3512),
.B(n_3186),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3703),
.B(n_3191),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3742),
.Y(n_3997)
);

INVx4_ASAP7_75t_L g3998 ( 
.A(n_3676),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3698),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3717),
.Y(n_4000)
);

INVx3_ASAP7_75t_L g4001 ( 
.A(n_3654),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3753),
.Y(n_4002)
);

BUFx3_ASAP7_75t_L g4003 ( 
.A(n_3752),
.Y(n_4003)
);

INVx3_ASAP7_75t_L g4004 ( 
.A(n_3680),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3606),
.B(n_3274),
.Y(n_4005)
);

BUFx3_ASAP7_75t_L g4006 ( 
.A(n_3540),
.Y(n_4006)
);

INVx5_ASAP7_75t_L g4007 ( 
.A(n_3608),
.Y(n_4007)
);

NOR2xp67_ASAP7_75t_L g4008 ( 
.A(n_3777),
.B(n_3072),
.Y(n_4008)
);

NOR2xp33_ASAP7_75t_L g4009 ( 
.A(n_3462),
.B(n_3129),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3759),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3786),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3790),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3701),
.Y(n_4013)
);

INVx3_ASAP7_75t_L g4014 ( 
.A(n_3680),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3795),
.Y(n_4015)
);

OR2x6_ASAP7_75t_L g4016 ( 
.A(n_3704),
.B(n_3099),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3479),
.B(n_3275),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3595),
.B(n_3283),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3708),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3616),
.B(n_3284),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3498),
.B(n_3294),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3594),
.B(n_3301),
.Y(n_4022)
);

BUFx6f_ASAP7_75t_L g4023 ( 
.A(n_3685),
.Y(n_4023)
);

AO22x1_ASAP7_75t_L g4024 ( 
.A1(n_3623),
.A2(n_3533),
.B1(n_3511),
.B2(n_3793),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3551),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3552),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3715),
.Y(n_4027)
);

AND2x4_ASAP7_75t_L g4028 ( 
.A(n_3667),
.B(n_3144),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3553),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3476),
.B(n_3387),
.Y(n_4030)
);

OAI21x1_ASAP7_75t_L g4031 ( 
.A1(n_3489),
.A2(n_3368),
.B(n_3355),
.Y(n_4031)
);

NOR2xp67_ASAP7_75t_L g4032 ( 
.A(n_3510),
.B(n_3173),
.Y(n_4032)
);

INVx1_ASAP7_75t_SL g4033 ( 
.A(n_3788),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3536),
.B(n_3387),
.Y(n_4034)
);

BUFx3_ASAP7_75t_L g4035 ( 
.A(n_3687),
.Y(n_4035)
);

INVx3_ASAP7_75t_SL g4036 ( 
.A(n_3732),
.Y(n_4036)
);

BUFx6f_ASAP7_75t_L g4037 ( 
.A(n_3685),
.Y(n_4037)
);

AOI22xp5_ASAP7_75t_L g4038 ( 
.A1(n_3737),
.A2(n_3238),
.B1(n_3267),
.B2(n_3117),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3562),
.Y(n_4039)
);

BUFx2_ASAP7_75t_L g4040 ( 
.A(n_3704),
.Y(n_4040)
);

BUFx2_ASAP7_75t_L g4041 ( 
.A(n_3704),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3726),
.Y(n_4042)
);

BUFx6f_ASAP7_75t_L g4043 ( 
.A(n_3685),
.Y(n_4043)
);

AND2x4_ASAP7_75t_L g4044 ( 
.A(n_3556),
.B(n_3150),
.Y(n_4044)
);

INVx2_ASAP7_75t_L g4045 ( 
.A(n_3731),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_SL g4046 ( 
.A(n_3716),
.B(n_3173),
.Y(n_4046)
);

AND2x4_ASAP7_75t_L g4047 ( 
.A(n_3636),
.B(n_3150),
.Y(n_4047)
);

AND2x4_ASAP7_75t_L g4048 ( 
.A(n_3573),
.B(n_3189),
.Y(n_4048)
);

HB1xp67_ASAP7_75t_L g4049 ( 
.A(n_3678),
.Y(n_4049)
);

AND2x2_ASAP7_75t_SL g4050 ( 
.A(n_3766),
.B(n_3125),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3536),
.B(n_3603),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3603),
.B(n_3400),
.Y(n_4052)
);

AND3x1_ASAP7_75t_SL g4053 ( 
.A(n_3772),
.B(n_1665),
.C(n_1662),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3499),
.B(n_3400),
.Y(n_4054)
);

BUFx6f_ASAP7_75t_L g4055 ( 
.A(n_3767),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3768),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3509),
.B(n_3189),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_3769),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3776),
.Y(n_4059)
);

AOI22xp33_ASAP7_75t_L g4060 ( 
.A1(n_3757),
.A2(n_3187),
.B1(n_3089),
.B2(n_3268),
.Y(n_4060)
);

NOR2xp33_ASAP7_75t_L g4061 ( 
.A(n_3625),
.B(n_3268),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3781),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_3808),
.B(n_1667),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3541),
.B(n_3515),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3782),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3796),
.Y(n_4066)
);

INVx2_ASAP7_75t_L g4067 ( 
.A(n_3798),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3805),
.Y(n_4068)
);

BUFx6f_ASAP7_75t_L g4069 ( 
.A(n_3767),
.Y(n_4069)
);

BUFx3_ASAP7_75t_L g4070 ( 
.A(n_3544),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3541),
.B(n_3310),
.Y(n_4071)
);

BUFx6f_ASAP7_75t_L g4072 ( 
.A(n_3767),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_SL g4073 ( 
.A(n_3766),
.B(n_3182),
.Y(n_4073)
);

BUFx6f_ASAP7_75t_L g4074 ( 
.A(n_3799),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3794),
.Y(n_4075)
);

BUFx6f_ASAP7_75t_L g4076 ( 
.A(n_3799),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_3628),
.B(n_3310),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3692),
.Y(n_4078)
);

INVx4_ASAP7_75t_L g4079 ( 
.A(n_3799),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3500),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3634),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_3765),
.B(n_1668),
.Y(n_4082)
);

INVxp67_ASAP7_75t_SL g4083 ( 
.A(n_3791),
.Y(n_4083)
);

BUFx4f_ASAP7_75t_L g4084 ( 
.A(n_3714),
.Y(n_4084)
);

INVx2_ASAP7_75t_SL g4085 ( 
.A(n_3714),
.Y(n_4085)
);

AOI22xp5_ASAP7_75t_L g4086 ( 
.A1(n_3739),
.A2(n_3182),
.B1(n_3361),
.B2(n_3320),
.Y(n_4086)
);

INVxp67_ASAP7_75t_L g4087 ( 
.A(n_3723),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3672),
.Y(n_4088)
);

INVx3_ASAP7_75t_L g4089 ( 
.A(n_3713),
.Y(n_4089)
);

AND2x2_ASAP7_75t_SL g4090 ( 
.A(n_3696),
.B(n_3336),
.Y(n_4090)
);

BUFx6f_ASAP7_75t_L g4091 ( 
.A(n_3571),
.Y(n_4091)
);

INVx2_ASAP7_75t_SL g4092 ( 
.A(n_3714),
.Y(n_4092)
);

BUFx6f_ASAP7_75t_L g4093 ( 
.A(n_3571),
.Y(n_4093)
);

INVx2_ASAP7_75t_L g4094 ( 
.A(n_3683),
.Y(n_4094)
);

BUFx2_ASAP7_75t_L g4095 ( 
.A(n_3458),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_SL g4096 ( 
.A(n_3495),
.B(n_3423),
.Y(n_4096)
);

BUFx4f_ASAP7_75t_L g4097 ( 
.A(n_3458),
.Y(n_4097)
);

AOI22xp5_ASAP7_75t_L g4098 ( 
.A1(n_3748),
.A2(n_3320),
.B1(n_3371),
.B2(n_3361),
.Y(n_4098)
);

BUFx12f_ASAP7_75t_SL g4099 ( 
.A(n_3783),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_SL g4100 ( 
.A(n_3696),
.B(n_3423),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_3774),
.Y(n_4101)
);

HB1xp67_ASAP7_75t_L g4102 ( 
.A(n_3868),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3839),
.Y(n_4103)
);

INVx3_ASAP7_75t_L g4104 ( 
.A(n_3904),
.Y(n_4104)
);

NOR2x1_ASAP7_75t_L g4105 ( 
.A(n_4070),
.B(n_3451),
.Y(n_4105)
);

NOR2xp33_ASAP7_75t_R g4106 ( 
.A(n_3810),
.B(n_3733),
.Y(n_4106)
);

BUFx4f_ASAP7_75t_L g4107 ( 
.A(n_3877),
.Y(n_4107)
);

BUFx6f_ASAP7_75t_SL g4108 ( 
.A(n_3860),
.Y(n_4108)
);

HB1xp67_ASAP7_75t_L g4109 ( 
.A(n_3815),
.Y(n_4109)
);

INVxp67_ASAP7_75t_L g4110 ( 
.A(n_3871),
.Y(n_4110)
);

BUFx6f_ASAP7_75t_L g4111 ( 
.A(n_3814),
.Y(n_4111)
);

BUFx6f_ASAP7_75t_L g4112 ( 
.A(n_3814),
.Y(n_4112)
);

A2O1A1Ixp33_ASAP7_75t_L g4113 ( 
.A1(n_3982),
.A2(n_3496),
.B(n_3487),
.C(n_3461),
.Y(n_4113)
);

AOI21x1_ASAP7_75t_L g4114 ( 
.A1(n_4024),
.A2(n_3461),
.B(n_3602),
.Y(n_4114)
);

OAI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3829),
.A2(n_3501),
.B1(n_3591),
.B2(n_3438),
.Y(n_4115)
);

INVx3_ASAP7_75t_L g4116 ( 
.A(n_3939),
.Y(n_4116)
);

AOI21xp5_ASAP7_75t_L g4117 ( 
.A1(n_4034),
.A2(n_3465),
.B(n_3433),
.Y(n_4117)
);

OAI21xp33_ASAP7_75t_L g4118 ( 
.A1(n_3823),
.A2(n_3682),
.B(n_3720),
.Y(n_4118)
);

OAI22xp5_ASAP7_75t_L g4119 ( 
.A1(n_4087),
.A2(n_3651),
.B1(n_3605),
.B2(n_3610),
.Y(n_4119)
);

AOI21xp5_ASAP7_75t_L g4120 ( 
.A1(n_4083),
.A2(n_3525),
.B(n_3528),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_SL g4121 ( 
.A1(n_3816),
.A2(n_3644),
.B1(n_3517),
.B2(n_3468),
.Y(n_4121)
);

AOI22x1_ASAP7_75t_L g4122 ( 
.A1(n_4082),
.A2(n_3626),
.B1(n_3705),
.B2(n_3700),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_SL g4123 ( 
.A(n_3961),
.B(n_3619),
.Y(n_4123)
);

AOI21xp5_ASAP7_75t_L g4124 ( 
.A1(n_3935),
.A2(n_3631),
.B(n_3583),
.Y(n_4124)
);

A2O1A1Ixp33_ASAP7_75t_L g4125 ( 
.A1(n_3994),
.A2(n_3545),
.B(n_3740),
.C(n_3549),
.Y(n_4125)
);

O2A1O1Ixp33_ASAP7_75t_L g4126 ( 
.A1(n_3966),
.A2(n_3754),
.B(n_3644),
.C(n_3780),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3954),
.B(n_3707),
.Y(n_4127)
);

A2O1A1Ixp33_ASAP7_75t_L g4128 ( 
.A1(n_3826),
.A2(n_3740),
.B(n_3638),
.C(n_3548),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3852),
.Y(n_4129)
);

NOR2xp33_ASAP7_75t_L g4130 ( 
.A(n_3811),
.B(n_3468),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3856),
.B(n_3519),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_4025),
.B(n_3519),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_3977),
.B(n_3604),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_3812),
.B(n_3635),
.Y(n_4134)
);

AOI21xp5_ASAP7_75t_L g4135 ( 
.A1(n_3942),
.A2(n_3586),
.B(n_3582),
.Y(n_4135)
);

BUFx3_ASAP7_75t_L g4136 ( 
.A(n_3862),
.Y(n_4136)
);

NOR2xp33_ASAP7_75t_L g4137 ( 
.A(n_3831),
.B(n_3527),
.Y(n_4137)
);

BUFx6f_ASAP7_75t_L g4138 ( 
.A(n_3814),
.Y(n_4138)
);

NOR3xp33_ASAP7_75t_SL g4139 ( 
.A(n_3952),
.B(n_3660),
.C(n_3659),
.Y(n_4139)
);

NOR2xp33_ASAP7_75t_L g4140 ( 
.A(n_3946),
.B(n_3617),
.Y(n_4140)
);

BUFx6f_ASAP7_75t_L g4141 ( 
.A(n_3820),
.Y(n_4141)
);

INVx2_ASAP7_75t_SL g4142 ( 
.A(n_3830),
.Y(n_4142)
);

INVx2_ASAP7_75t_SL g4143 ( 
.A(n_3809),
.Y(n_4143)
);

A2O1A1Ixp33_ASAP7_75t_SL g4144 ( 
.A1(n_3973),
.A2(n_3738),
.B(n_3679),
.C(n_3460),
.Y(n_4144)
);

AOI21xp5_ASAP7_75t_L g4145 ( 
.A1(n_4054),
.A2(n_4021),
.B(n_3996),
.Y(n_4145)
);

BUFx6f_ASAP7_75t_L g4146 ( 
.A(n_3820),
.Y(n_4146)
);

A2O1A1Ixp33_ASAP7_75t_L g4147 ( 
.A1(n_4061),
.A2(n_3883),
.B(n_3822),
.C(n_3978),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_4026),
.B(n_3450),
.Y(n_4148)
);

O2A1O1Ixp5_ASAP7_75t_L g4149 ( 
.A1(n_4024),
.A2(n_3531),
.B(n_3734),
.C(n_3526),
.Y(n_4149)
);

A2O1A1Ixp33_ASAP7_75t_SL g4150 ( 
.A1(n_4009),
.A2(n_3848),
.B(n_3894),
.C(n_4060),
.Y(n_4150)
);

BUFx3_ASAP7_75t_L g4151 ( 
.A(n_3914),
.Y(n_4151)
);

NOR2xp33_ASAP7_75t_SL g4152 ( 
.A(n_3845),
.B(n_3713),
.Y(n_4152)
);

INVx3_ASAP7_75t_L g4153 ( 
.A(n_4035),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_4029),
.B(n_3761),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_L g4155 ( 
.A(n_4075),
.B(n_4078),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3818),
.Y(n_4156)
);

OAI21x1_ASAP7_75t_L g4157 ( 
.A1(n_4031),
.A2(n_3679),
.B(n_3521),
.Y(n_4157)
);

BUFx5_ASAP7_75t_L g4158 ( 
.A(n_3975),
.Y(n_4158)
);

HB1xp67_ASAP7_75t_L g4159 ( 
.A(n_3919),
.Y(n_4159)
);

AOI21xp5_ASAP7_75t_L g4160 ( 
.A1(n_3974),
.A2(n_3589),
.B(n_3532),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_3867),
.B(n_3995),
.Y(n_4161)
);

OAI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_3824),
.A2(n_3546),
.B(n_3775),
.Y(n_4162)
);

CKINVDCx5p33_ASAP7_75t_R g4163 ( 
.A(n_3847),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_4088),
.B(n_3764),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_4094),
.B(n_3607),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_3870),
.B(n_3564),
.Y(n_4166)
);

BUFx12f_ASAP7_75t_L g4167 ( 
.A(n_3927),
.Y(n_4167)
);

INVx4_ASAP7_75t_L g4168 ( 
.A(n_3817),
.Y(n_4168)
);

AND2x2_ASAP7_75t_L g4169 ( 
.A(n_4063),
.B(n_3535),
.Y(n_4169)
);

NOR2xp33_ASAP7_75t_L g4170 ( 
.A(n_3840),
.B(n_3535),
.Y(n_4170)
);

AOI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_3898),
.A2(n_3590),
.B1(n_3585),
.B2(n_3534),
.Y(n_4171)
);

O2A1O1Ixp33_ASAP7_75t_L g4172 ( 
.A1(n_3885),
.A2(n_3563),
.B(n_1672),
.C(n_1674),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3819),
.Y(n_4173)
);

AOI21xp5_ASAP7_75t_L g4174 ( 
.A1(n_3889),
.A2(n_3580),
.B(n_3442),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3821),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_SL g4176 ( 
.A(n_3838),
.B(n_3841),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_3849),
.B(n_3697),
.Y(n_4177)
);

OAI22xp5_ASAP7_75t_L g4178 ( 
.A1(n_3909),
.A2(n_3516),
.B1(n_3630),
.B2(n_3652),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_3851),
.B(n_3699),
.Y(n_4179)
);

A2O1A1Ixp33_ASAP7_75t_L g4180 ( 
.A1(n_4038),
.A2(n_3621),
.B(n_3633),
.C(n_3526),
.Y(n_4180)
);

OAI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_3911),
.A2(n_3694),
.B1(n_3574),
.B2(n_3609),
.Y(n_4181)
);

INVx6_ASAP7_75t_L g4182 ( 
.A(n_3865),
.Y(n_4182)
);

OR2x6_ASAP7_75t_L g4183 ( 
.A(n_3899),
.B(n_3763),
.Y(n_4183)
);

AOI22xp5_ASAP7_75t_L g4184 ( 
.A1(n_4006),
.A2(n_3749),
.B1(n_3618),
.B2(n_3691),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3859),
.Y(n_4185)
);

O2A1O1Ixp5_ASAP7_75t_SL g4186 ( 
.A1(n_3979),
.A2(n_3543),
.B(n_3576),
.C(n_1676),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3833),
.Y(n_4187)
);

O2A1O1Ixp33_ASAP7_75t_SL g4188 ( 
.A1(n_4100),
.A2(n_3929),
.B(n_4073),
.C(n_4046),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_3835),
.Y(n_4189)
);

AOI21xp5_ASAP7_75t_L g4190 ( 
.A1(n_3896),
.A2(n_3442),
.B(n_3642),
.Y(n_4190)
);

AO32x2_ASAP7_75t_L g4191 ( 
.A1(n_4085),
.A2(n_3543),
.A3(n_3576),
.B1(n_3394),
.B2(n_3376),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3837),
.Y(n_4192)
);

INVx11_ASAP7_75t_L g4193 ( 
.A(n_4097),
.Y(n_4193)
);

NOR2xp33_ASAP7_75t_R g4194 ( 
.A(n_3853),
.B(n_3624),
.Y(n_4194)
);

OAI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_3866),
.A2(n_3601),
.B1(n_3744),
.B2(n_3642),
.Y(n_4195)
);

AOI21xp5_ASAP7_75t_L g4196 ( 
.A1(n_3900),
.A2(n_3657),
.B(n_3653),
.Y(n_4196)
);

INVxp67_ASAP7_75t_L g4197 ( 
.A(n_3922),
.Y(n_4197)
);

AOI21xp5_ASAP7_75t_L g4198 ( 
.A1(n_4051),
.A2(n_3657),
.B(n_3653),
.Y(n_4198)
);

AOI21xp5_ASAP7_75t_L g4199 ( 
.A1(n_4052),
.A2(n_3908),
.B(n_4064),
.Y(n_4199)
);

AOI21xp5_ASAP7_75t_L g4200 ( 
.A1(n_4071),
.A2(n_3423),
.B(n_3668),
.Y(n_4200)
);

NOR2x1_ASAP7_75t_L g4201 ( 
.A(n_3817),
.B(n_3624),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_3861),
.B(n_3728),
.Y(n_4202)
);

INVx5_ASAP7_75t_L g4203 ( 
.A(n_3970),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_4039),
.B(n_3730),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_4049),
.B(n_3735),
.Y(n_4205)
);

A2O1A1Ixp33_ASAP7_75t_L g4206 ( 
.A1(n_4080),
.A2(n_3588),
.B(n_3289),
.C(n_3741),
.Y(n_4206)
);

OAI22xp5_ASAP7_75t_L g4207 ( 
.A1(n_3850),
.A2(n_3792),
.B1(n_3803),
.B2(n_3797),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_4081),
.B(n_3743),
.Y(n_4208)
);

BUFx6f_ASAP7_75t_L g4209 ( 
.A(n_3820),
.Y(n_4209)
);

AOI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_3975),
.A2(n_3336),
.B(n_3662),
.Y(n_4210)
);

O2A1O1Ixp33_ASAP7_75t_L g4211 ( 
.A1(n_4096),
.A2(n_1670),
.B(n_3554),
.C(n_3746),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_4000),
.A2(n_3664),
.B(n_3662),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_3916),
.B(n_3763),
.Y(n_4213)
);

A2O1A1Ixp33_ASAP7_75t_L g4214 ( 
.A1(n_4077),
.A2(n_3289),
.B(n_3750),
.C(n_3747),
.Y(n_4214)
);

AOI33xp33_ASAP7_75t_L g4215 ( 
.A1(n_3989),
.A2(n_1157),
.A3(n_1152),
.B1(n_1158),
.B2(n_1153),
.B3(n_1150),
.Y(n_4215)
);

NOR2xp33_ASAP7_75t_L g4216 ( 
.A(n_4033),
.B(n_3641),
.Y(n_4216)
);

OAI22xp5_ASAP7_75t_L g4217 ( 
.A1(n_3910),
.A2(n_3756),
.B1(n_3391),
.B2(n_3770),
.Y(n_4217)
);

BUFx3_ASAP7_75t_L g4218 ( 
.A(n_3890),
.Y(n_4218)
);

AND2x2_ASAP7_75t_L g4219 ( 
.A(n_3836),
.B(n_3641),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_3828),
.B(n_3646),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_3875),
.B(n_3646),
.Y(n_4221)
);

OR2x2_ASAP7_75t_L g4222 ( 
.A(n_3854),
.B(n_3643),
.Y(n_4222)
);

A2O1A1Ixp33_ASAP7_75t_L g4223 ( 
.A1(n_4008),
.A2(n_3643),
.B(n_3645),
.C(n_3143),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_3864),
.Y(n_4224)
);

INVx4_ASAP7_75t_L g4225 ( 
.A(n_3873),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4090),
.B(n_1894),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_SL g4227 ( 
.A(n_3916),
.B(n_3645),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_4000),
.A2(n_3686),
.B(n_3664),
.Y(n_4228)
);

BUFx6f_ASAP7_75t_L g4229 ( 
.A(n_3832),
.Y(n_4229)
);

O2A1O1Ixp33_ASAP7_75t_L g4230 ( 
.A1(n_4018),
.A2(n_3650),
.B(n_3669),
.C(n_3779),
.Y(n_4230)
);

INVx2_ASAP7_75t_L g4231 ( 
.A(n_3884),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_3846),
.Y(n_4232)
);

OAI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_4020),
.A2(n_3650),
.B(n_3143),
.Y(n_4233)
);

NOR2x1_ASAP7_75t_R g4234 ( 
.A(n_3891),
.B(n_1158),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_3984),
.B(n_1894),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_3945),
.B(n_3686),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_3893),
.B(n_1907),
.Y(n_4237)
);

NAND2xp5_ASAP7_75t_L g4238 ( 
.A(n_4022),
.B(n_3371),
.Y(n_4238)
);

AOI21xp33_ASAP7_75t_L g4239 ( 
.A1(n_4057),
.A2(n_3785),
.B(n_3784),
.Y(n_4239)
);

NOR2xp33_ASAP7_75t_L g4240 ( 
.A(n_3834),
.B(n_3388),
.Y(n_4240)
);

NOR2xp33_ASAP7_75t_L g4241 ( 
.A(n_3969),
.B(n_3388),
.Y(n_4241)
);

AND2x4_ASAP7_75t_L g4242 ( 
.A(n_3827),
.B(n_3357),
.Y(n_4242)
);

A2O1A1Ixp33_ASAP7_75t_L g4243 ( 
.A1(n_4047),
.A2(n_3771),
.B(n_3207),
.C(n_3710),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4005),
.B(n_1157),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_L g4245 ( 
.A(n_3965),
.B(n_1026),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_3906),
.Y(n_4246)
);

BUFx6f_ASAP7_75t_L g4247 ( 
.A(n_3832),
.Y(n_4247)
);

INVx4_ASAP7_75t_L g4248 ( 
.A(n_3873),
.Y(n_4248)
);

AOI21xp5_ASAP7_75t_L g4249 ( 
.A1(n_4017),
.A2(n_3022),
.B(n_2994),
.Y(n_4249)
);

BUFx2_ASAP7_75t_L g4250 ( 
.A(n_3878),
.Y(n_4250)
);

A2O1A1Ixp33_ASAP7_75t_L g4251 ( 
.A1(n_4047),
.A2(n_3199),
.B(n_3228),
.C(n_3224),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_3924),
.Y(n_4252)
);

AOI21xp5_ASAP7_75t_L g4253 ( 
.A1(n_4030),
.A2(n_3022),
.B(n_2994),
.Y(n_4253)
);

AND2x4_ASAP7_75t_L g4254 ( 
.A(n_3844),
.B(n_3357),
.Y(n_4254)
);

NOR2xp33_ASAP7_75t_L g4255 ( 
.A(n_3972),
.B(n_1027),
.Y(n_4255)
);

OR2x6_ASAP7_75t_L g4256 ( 
.A(n_3899),
.B(n_3695),
.Y(n_4256)
);

NOR2xp33_ASAP7_75t_L g4257 ( 
.A(n_3912),
.B(n_1028),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_3970),
.A2(n_4007),
.B(n_4050),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_3925),
.Y(n_4259)
);

HB1xp67_ASAP7_75t_L g4260 ( 
.A(n_3948),
.Y(n_4260)
);

OAI22xp5_ASAP7_75t_L g4261 ( 
.A1(n_4016),
.A2(n_3337),
.B1(n_3097),
.B2(n_3091),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_3825),
.B(n_1159),
.Y(n_4262)
);

NAND2xp5_ASAP7_75t_L g4263 ( 
.A(n_4101),
.B(n_1159),
.Y(n_4263)
);

HB1xp67_ASAP7_75t_L g4264 ( 
.A(n_3991),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_3932),
.B(n_1162),
.Y(n_4265)
);

NOR2xp33_ASAP7_75t_L g4266 ( 
.A(n_4036),
.B(n_1029),
.Y(n_4266)
);

AOI21xp5_ASAP7_75t_L g4267 ( 
.A1(n_3970),
.A2(n_3000),
.B(n_2992),
.Y(n_4267)
);

BUFx6f_ASAP7_75t_L g4268 ( 
.A(n_3832),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_3858),
.Y(n_4269)
);

AOI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_4007),
.A2(n_3000),
.B(n_2992),
.Y(n_4270)
);

AND2x2_ASAP7_75t_L g4271 ( 
.A(n_3944),
.B(n_1907),
.Y(n_4271)
);

NOR2xp33_ASAP7_75t_L g4272 ( 
.A(n_3923),
.B(n_1034),
.Y(n_4272)
);

O2A1O1Ixp33_ASAP7_75t_L g4273 ( 
.A1(n_4092),
.A2(n_3787),
.B(n_3802),
.C(n_3674),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_SL g4274 ( 
.A(n_4084),
.B(n_3099),
.Y(n_4274)
);

A2O1A1Ixp33_ASAP7_75t_L g4275 ( 
.A1(n_4098),
.A2(n_3677),
.B(n_3722),
.C(n_3665),
.Y(n_4275)
);

OAI222xp33_ASAP7_75t_L g4276 ( 
.A1(n_3934),
.A2(n_1169),
.B1(n_1167),
.B2(n_1170),
.C1(n_1168),
.C2(n_1163),
.Y(n_4276)
);

BUFx3_ASAP7_75t_L g4277 ( 
.A(n_4003),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_SL g4278 ( 
.A(n_4044),
.B(n_3099),
.Y(n_4278)
);

AOI21xp5_ASAP7_75t_L g4279 ( 
.A1(n_4007),
.A2(n_3027),
.B(n_3278),
.Y(n_4279)
);

AOI21xp33_ASAP7_75t_L g4280 ( 
.A1(n_4044),
.A2(n_3368),
.B(n_3355),
.Y(n_4280)
);

HB1xp67_ASAP7_75t_L g4281 ( 
.A(n_4095),
.Y(n_4281)
);

AOI22xp33_ASAP7_75t_L g4282 ( 
.A1(n_4040),
.A2(n_3691),
.B1(n_3369),
.B2(n_3367),
.Y(n_4282)
);

OAI22xp5_ASAP7_75t_L g4283 ( 
.A1(n_4016),
.A2(n_3411),
.B1(n_3376),
.B2(n_3127),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3876),
.Y(n_4284)
);

NOR2xp33_ASAP7_75t_L g4285 ( 
.A(n_4028),
.B(n_4041),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_3879),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_3949),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3950),
.B(n_1163),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_3951),
.B(n_1167),
.Y(n_4289)
);

AOI21xp5_ASAP7_75t_L g4290 ( 
.A1(n_3980),
.A2(n_3027),
.B(n_3278),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_3881),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_SL g4292 ( 
.A(n_3990),
.B(n_3127),
.Y(n_4292)
);

AOI21xp5_ASAP7_75t_L g4293 ( 
.A1(n_4086),
.A2(n_3318),
.B(n_3290),
.Y(n_4293)
);

OR2x6_ASAP7_75t_SL g4294 ( 
.A(n_3993),
.B(n_1168),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_3955),
.B(n_1169),
.Y(n_4295)
);

AOI21xp5_ASAP7_75t_L g4296 ( 
.A1(n_3962),
.A2(n_3318),
.B(n_3290),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_3956),
.B(n_1170),
.Y(n_4297)
);

AOI21xp5_ASAP7_75t_L g4298 ( 
.A1(n_3962),
.A2(n_3381),
.B(n_3375),
.Y(n_4298)
);

NOR2xp33_ASAP7_75t_L g4299 ( 
.A(n_4028),
.B(n_1035),
.Y(n_4299)
);

AOI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_3953),
.A2(n_3381),
.B(n_3375),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_3976),
.B(n_1172),
.Y(n_4301)
);

INVx3_ASAP7_75t_L g4302 ( 
.A(n_4091),
.Y(n_4302)
);

OAI21x1_ASAP7_75t_SL g4303 ( 
.A1(n_3905),
.A2(n_3411),
.B(n_3608),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_3981),
.Y(n_4304)
);

A2O1A1Ixp33_ASAP7_75t_L g4305 ( 
.A1(n_4032),
.A2(n_3745),
.B(n_3760),
.C(n_3736),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_3983),
.B(n_1172),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_3987),
.B(n_1174),
.Y(n_4307)
);

AOI22xp5_ASAP7_75t_L g4308 ( 
.A1(n_3844),
.A2(n_3691),
.B1(n_1037),
.B2(n_1039),
.Y(n_4308)
);

NOR2x1_ASAP7_75t_L g4309 ( 
.A(n_3880),
.B(n_3778),
.Y(n_4309)
);

A2O1A1Ixp33_ASAP7_75t_L g4310 ( 
.A1(n_3886),
.A2(n_3130),
.B(n_3181),
.C(n_3127),
.Y(n_4310)
);

HB1xp67_ASAP7_75t_L g4311 ( 
.A(n_3971),
.Y(n_4311)
);

NOR2xp33_ASAP7_75t_L g4312 ( 
.A(n_3990),
.B(n_1036),
.Y(n_4312)
);

INVx1_ASAP7_75t_SL g4313 ( 
.A(n_3813),
.Y(n_4313)
);

O2A1O1Ixp33_ASAP7_75t_L g4314 ( 
.A1(n_3887),
.A2(n_1968),
.B(n_1962),
.C(n_3695),
.Y(n_4314)
);

A2O1A1Ixp33_ASAP7_75t_L g4315 ( 
.A1(n_3895),
.A2(n_3181),
.B(n_3184),
.C(n_3130),
.Y(n_4315)
);

AOI21xp5_ASAP7_75t_L g4316 ( 
.A1(n_3953),
.A2(n_3181),
.B(n_3130),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_3897),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_3999),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_3901),
.Y(n_4319)
);

AOI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_3967),
.A2(n_3221),
.B(n_3184),
.Y(n_4320)
);

AOI21xp5_ASAP7_75t_L g4321 ( 
.A1(n_3967),
.A2(n_3221),
.B(n_3184),
.Y(n_4321)
);

BUFx6f_ASAP7_75t_L g4322 ( 
.A(n_3842),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_3903),
.A2(n_3241),
.B(n_3221),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4013),
.B(n_1962),
.Y(n_4324)
);

BUFx12f_ASAP7_75t_L g4325 ( 
.A(n_3857),
.Y(n_4325)
);

AO21x1_ASAP7_75t_L g4326 ( 
.A1(n_3902),
.A2(n_3369),
.B(n_3367),
.Y(n_4326)
);

A2O1A1Ixp33_ASAP7_75t_L g4327 ( 
.A1(n_3907),
.A2(n_3244),
.B(n_3252),
.C(n_3241),
.Y(n_4327)
);

A2O1A1Ixp33_ASAP7_75t_L g4328 ( 
.A1(n_3913),
.A2(n_3244),
.B(n_3252),
.C(n_3241),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3921),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4019),
.B(n_1968),
.Y(n_4330)
);

OAI21x1_ASAP7_75t_L g4331 ( 
.A1(n_3843),
.A2(n_2439),
.B(n_2391),
.Y(n_4331)
);

OR2x6_ASAP7_75t_L g4332 ( 
.A(n_3903),
.B(n_3244),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_3926),
.Y(n_4333)
);

NAND3xp33_ASAP7_75t_L g4334 ( 
.A(n_4056),
.B(n_1175),
.C(n_1174),
.Y(n_4334)
);

AOI21xp5_ASAP7_75t_L g4335 ( 
.A1(n_3986),
.A2(n_3258),
.B(n_3252),
.Y(n_4335)
);

AOI21xp5_ASAP7_75t_L g4336 ( 
.A1(n_3986),
.A2(n_4004),
.B(n_4001),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_3936),
.Y(n_4337)
);

O2A1O1Ixp33_ASAP7_75t_L g4338 ( 
.A1(n_3947),
.A2(n_2391),
.B(n_2449),
.C(n_2439),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_4001),
.A2(n_4014),
.B(n_4004),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_SL g4340 ( 
.A(n_3920),
.B(n_3258),
.Y(n_4340)
);

CKINVDCx5p33_ASAP7_75t_R g4341 ( 
.A(n_3888),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_4027),
.B(n_1175),
.Y(n_4342)
);

HB1xp67_ASAP7_75t_L g4343 ( 
.A(n_3960),
.Y(n_4343)
);

AND2x4_ASAP7_75t_L g4344 ( 
.A(n_3855),
.B(n_3258),
.Y(n_4344)
);

OAI22xp5_ASAP7_75t_L g4345 ( 
.A1(n_3968),
.A2(n_3265),
.B1(n_3280),
.B2(n_3261),
.Y(n_4345)
);

A2O1A1Ixp33_ASAP7_75t_L g4346 ( 
.A1(n_3985),
.A2(n_3265),
.B(n_3280),
.C(n_3261),
.Y(n_4346)
);

AOI21xp5_ASAP7_75t_L g4347 ( 
.A1(n_4014),
.A2(n_3265),
.B(n_3261),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4042),
.B(n_1176),
.Y(n_4348)
);

AOI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_4089),
.A2(n_3288),
.B(n_3280),
.Y(n_4349)
);

NOR2xp33_ASAP7_75t_R g4350 ( 
.A(n_4099),
.B(n_3608),
.Y(n_4350)
);

AOI21x1_ASAP7_75t_L g4351 ( 
.A1(n_3988),
.A2(n_3369),
.B(n_3367),
.Y(n_4351)
);

A2O1A1Ixp33_ASAP7_75t_L g4352 ( 
.A1(n_3997),
.A2(n_3351),
.B(n_3360),
.C(n_3288),
.Y(n_4352)
);

NOR3xp33_ASAP7_75t_SL g4353 ( 
.A(n_3863),
.B(n_1178),
.C(n_1176),
.Y(n_4353)
);

NOR2xp33_ASAP7_75t_L g4354 ( 
.A(n_4045),
.B(n_1040),
.Y(n_4354)
);

NAND2x1p5_ASAP7_75t_L g4355 ( 
.A(n_3882),
.B(n_3288),
.Y(n_4355)
);

NAND2xp5_ASAP7_75t_L g4356 ( 
.A(n_4058),
.B(n_1178),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_SL g4357 ( 
.A(n_3920),
.B(n_3360),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4002),
.Y(n_4358)
);

AND2x4_ASAP7_75t_L g4359 ( 
.A(n_3855),
.B(n_3351),
.Y(n_4359)
);

INVx4_ASAP7_75t_L g4360 ( 
.A(n_3880),
.Y(n_4360)
);

INVx2_ASAP7_75t_L g4361 ( 
.A(n_4065),
.Y(n_4361)
);

O2A1O1Ixp33_ASAP7_75t_L g4362 ( 
.A1(n_4010),
.A2(n_2391),
.B(n_2449),
.C(n_2439),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4067),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_L g4364 ( 
.A(n_4059),
.B(n_1179),
.Y(n_4364)
);

BUFx4f_ASAP7_75t_SL g4365 ( 
.A(n_3930),
.Y(n_4365)
);

AOI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_4089),
.A2(n_3360),
.B(n_3351),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4062),
.B(n_1179),
.Y(n_4367)
);

O2A1O1Ixp33_ASAP7_75t_L g4368 ( 
.A1(n_4011),
.A2(n_2463),
.B(n_2464),
.C(n_2449),
.Y(n_4368)
);

OR2x6_ASAP7_75t_L g4369 ( 
.A(n_3905),
.B(n_3931),
.Y(n_4369)
);

AND2x2_ASAP7_75t_L g4370 ( 
.A(n_4066),
.B(n_2017),
.Y(n_4370)
);

BUFx2_ASAP7_75t_L g4371 ( 
.A(n_4158),
.Y(n_4371)
);

OR2x6_ASAP7_75t_L g4372 ( 
.A(n_4258),
.B(n_3931),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4176),
.B(n_4012),
.Y(n_4373)
);

BUFx2_ASAP7_75t_L g4374 ( 
.A(n_4158),
.Y(n_4374)
);

OAI221xp5_ASAP7_75t_L g4375 ( 
.A1(n_4118),
.A2(n_1193),
.B1(n_1194),
.B2(n_1188),
.C(n_1184),
.Y(n_4375)
);

AND2x4_ASAP7_75t_L g4376 ( 
.A(n_4183),
.B(n_4256),
.Y(n_4376)
);

INVx2_ASAP7_75t_SL g4377 ( 
.A(n_4182),
.Y(n_4377)
);

BUFx6f_ASAP7_75t_L g4378 ( 
.A(n_4182),
.Y(n_4378)
);

AOI22xp33_ASAP7_75t_L g4379 ( 
.A1(n_4272),
.A2(n_3928),
.B1(n_4068),
.B2(n_3915),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4343),
.Y(n_4380)
);

INVxp67_ASAP7_75t_L g4381 ( 
.A(n_4102),
.Y(n_4381)
);

NAND3xp33_ASAP7_75t_L g4382 ( 
.A(n_4126),
.B(n_1188),
.C(n_1184),
.Y(n_4382)
);

BUFx2_ASAP7_75t_L g4383 ( 
.A(n_4158),
.Y(n_4383)
);

AOI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_4123),
.A2(n_3928),
.B1(n_3915),
.B2(n_3874),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4185),
.Y(n_4385)
);

OR2x2_ASAP7_75t_L g4386 ( 
.A(n_4222),
.B(n_4015),
.Y(n_4386)
);

INVx2_ASAP7_75t_L g4387 ( 
.A(n_4224),
.Y(n_4387)
);

INVx2_ASAP7_75t_L g4388 ( 
.A(n_4231),
.Y(n_4388)
);

AOI22xp5_ASAP7_75t_L g4389 ( 
.A1(n_4137),
.A2(n_4053),
.B1(n_3943),
.B2(n_3874),
.Y(n_4389)
);

NOR2xp33_ASAP7_75t_L g4390 ( 
.A(n_4127),
.B(n_3892),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4246),
.Y(n_4391)
);

AO22x1_ASAP7_75t_L g4392 ( 
.A1(n_4130),
.A2(n_3918),
.B1(n_3933),
.B2(n_3882),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4156),
.Y(n_4393)
);

AOI22xp33_ASAP7_75t_L g4394 ( 
.A1(n_4115),
.A2(n_1194),
.B1(n_1201),
.B2(n_1193),
.Y(n_4394)
);

BUFx2_ASAP7_75t_L g4395 ( 
.A(n_4158),
.Y(n_4395)
);

INVx4_ASAP7_75t_L g4396 ( 
.A(n_4193),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_4252),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_SL g4398 ( 
.A(n_4105),
.B(n_4048),
.Y(n_4398)
);

NOR2xp33_ASAP7_75t_L g4399 ( 
.A(n_4313),
.B(n_4048),
.Y(n_4399)
);

INVxp67_ASAP7_75t_SL g4400 ( 
.A(n_4109),
.Y(n_4400)
);

BUFx12f_ASAP7_75t_L g4401 ( 
.A(n_4163),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4173),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4175),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4187),
.Y(n_4404)
);

BUFx2_ASAP7_75t_L g4405 ( 
.A(n_4191),
.Y(n_4405)
);

CKINVDCx5p33_ASAP7_75t_R g4406 ( 
.A(n_4341),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4259),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_4189),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4192),
.Y(n_4409)
);

INVx2_ASAP7_75t_SL g4410 ( 
.A(n_4218),
.Y(n_4410)
);

AND2x2_ASAP7_75t_L g4411 ( 
.A(n_4161),
.B(n_3842),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_4165),
.B(n_3842),
.Y(n_4412)
);

AOI22xp33_ASAP7_75t_L g4413 ( 
.A1(n_4121),
.A2(n_4325),
.B1(n_4226),
.B2(n_4299),
.Y(n_4413)
);

OR2x2_ASAP7_75t_L g4414 ( 
.A(n_4155),
.B(n_3938),
.Y(n_4414)
);

BUFx2_ASAP7_75t_L g4415 ( 
.A(n_4191),
.Y(n_4415)
);

OAI22xp5_ASAP7_75t_L g4416 ( 
.A1(n_4171),
.A2(n_3918),
.B1(n_3933),
.B2(n_3882),
.Y(n_4416)
);

INVx6_ASAP7_75t_L g4417 ( 
.A(n_4151),
.Y(n_4417)
);

AOI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_4196),
.A2(n_3933),
.B(n_3918),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4232),
.Y(n_4419)
);

INVx4_ASAP7_75t_L g4420 ( 
.A(n_4108),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4269),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4133),
.B(n_3938),
.Y(n_4422)
);

OR2x6_ASAP7_75t_L g4423 ( 
.A(n_4183),
.B(n_3940),
.Y(n_4423)
);

INVx4_ASAP7_75t_L g4424 ( 
.A(n_4104),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4284),
.Y(n_4425)
);

AOI22xp5_ASAP7_75t_L g4426 ( 
.A1(n_4266),
.A2(n_3917),
.B1(n_1042),
.B2(n_1044),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_4287),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_4199),
.B(n_3938),
.Y(n_4428)
);

BUFx6f_ASAP7_75t_L g4429 ( 
.A(n_4111),
.Y(n_4429)
);

AOI21xp5_ASAP7_75t_L g4430 ( 
.A1(n_4145),
.A2(n_3963),
.B(n_3380),
.Y(n_4430)
);

INVx5_ASAP7_75t_L g4431 ( 
.A(n_4203),
.Y(n_4431)
);

INVx2_ASAP7_75t_SL g4432 ( 
.A(n_4277),
.Y(n_4432)
);

HB1xp67_ASAP7_75t_L g4433 ( 
.A(n_4281),
.Y(n_4433)
);

INVx2_ASAP7_75t_L g4434 ( 
.A(n_4304),
.Y(n_4434)
);

AOI21xp5_ASAP7_75t_L g4435 ( 
.A1(n_4198),
.A2(n_3380),
.B(n_3362),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_4286),
.Y(n_4436)
);

OR2x6_ASAP7_75t_L g4437 ( 
.A(n_4369),
.B(n_3940),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4177),
.B(n_3941),
.Y(n_4438)
);

BUFx3_ASAP7_75t_L g4439 ( 
.A(n_4136),
.Y(n_4439)
);

BUFx3_ASAP7_75t_L g4440 ( 
.A(n_4116),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4318),
.Y(n_4441)
);

NOR2xp33_ASAP7_75t_L g4442 ( 
.A(n_4110),
.B(n_3941),
.Y(n_4442)
);

HB1xp67_ASAP7_75t_L g4443 ( 
.A(n_4159),
.Y(n_4443)
);

AOI22xp33_ASAP7_75t_L g4444 ( 
.A1(n_4162),
.A2(n_1201),
.B1(n_1202),
.B2(n_1195),
.Y(n_4444)
);

A2O1A1Ixp33_ASAP7_75t_L g4445 ( 
.A1(n_4113),
.A2(n_3872),
.B(n_3937),
.C(n_3843),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4361),
.Y(n_4446)
);

CKINVDCx5p33_ASAP7_75t_R g4447 ( 
.A(n_4194),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4363),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4219),
.B(n_3941),
.Y(n_4449)
);

OR2x6_ASAP7_75t_L g4450 ( 
.A(n_4369),
.B(n_3872),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4103),
.Y(n_4451)
);

BUFx4f_ASAP7_75t_L g4452 ( 
.A(n_4167),
.Y(n_4452)
);

AOI21xp5_ASAP7_75t_L g4453 ( 
.A1(n_4212),
.A2(n_3380),
.B(n_3362),
.Y(n_4453)
);

BUFx3_ASAP7_75t_L g4454 ( 
.A(n_4153),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4129),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_4169),
.B(n_3957),
.Y(n_4456)
);

HB1xp67_ASAP7_75t_L g4457 ( 
.A(n_4220),
.Y(n_4457)
);

BUFx6f_ASAP7_75t_L g4458 ( 
.A(n_4111),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4291),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4317),
.Y(n_4460)
);

AOI21xp33_ASAP7_75t_L g4461 ( 
.A1(n_4150),
.A2(n_3937),
.B(n_3917),
.Y(n_4461)
);

BUFx6f_ASAP7_75t_L g4462 ( 
.A(n_4111),
.Y(n_4462)
);

INVx3_ASAP7_75t_L g4463 ( 
.A(n_4302),
.Y(n_4463)
);

CKINVDCx6p67_ASAP7_75t_R g4464 ( 
.A(n_4203),
.Y(n_4464)
);

BUFx3_ASAP7_75t_L g4465 ( 
.A(n_4250),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4319),
.Y(n_4466)
);

BUFx12f_ASAP7_75t_L g4467 ( 
.A(n_4142),
.Y(n_4467)
);

INVx2_ASAP7_75t_SL g4468 ( 
.A(n_4143),
.Y(n_4468)
);

CKINVDCx11_ASAP7_75t_R g4469 ( 
.A(n_4294),
.Y(n_4469)
);

INVx1_ASAP7_75t_SL g4470 ( 
.A(n_4260),
.Y(n_4470)
);

AOI21xp5_ASAP7_75t_L g4471 ( 
.A1(n_4228),
.A2(n_3404),
.B(n_3362),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_4179),
.B(n_3957),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4170),
.B(n_3957),
.Y(n_4473)
);

BUFx6f_ASAP7_75t_L g4474 ( 
.A(n_4112),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4329),
.Y(n_4475)
);

AOI22xp5_ASAP7_75t_L g4476 ( 
.A1(n_4140),
.A2(n_1046),
.B1(n_1049),
.B2(n_1041),
.Y(n_4476)
);

AOI22xp5_ASAP7_75t_L g4477 ( 
.A1(n_4308),
.A2(n_1051),
.B1(n_1053),
.B2(n_1050),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_4333),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4202),
.B(n_3958),
.Y(n_4479)
);

BUFx2_ASAP7_75t_L g4480 ( 
.A(n_4191),
.Y(n_4480)
);

AND2x2_ASAP7_75t_L g4481 ( 
.A(n_4353),
.B(n_3958),
.Y(n_4481)
);

INVx8_ASAP7_75t_L g4482 ( 
.A(n_4203),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4205),
.B(n_3958),
.Y(n_4483)
);

BUFx6f_ASAP7_75t_L g4484 ( 
.A(n_4112),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_4154),
.B(n_3959),
.Y(n_4485)
);

AOI22xp33_ASAP7_75t_L g4486 ( 
.A1(n_4312),
.A2(n_1202),
.B1(n_1204),
.B2(n_1195),
.Y(n_4486)
);

INVx2_ASAP7_75t_SL g4487 ( 
.A(n_4311),
.Y(n_4487)
);

A2O1A1Ixp33_ASAP7_75t_SL g4488 ( 
.A1(n_4245),
.A2(n_2464),
.B(n_2471),
.C(n_2463),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_4337),
.Y(n_4489)
);

AND2x4_ASAP7_75t_L g4490 ( 
.A(n_4256),
.B(n_3998),
.Y(n_4490)
);

BUFx2_ASAP7_75t_L g4491 ( 
.A(n_4358),
.Y(n_4491)
);

HB1xp67_ASAP7_75t_L g4492 ( 
.A(n_4197),
.Y(n_4492)
);

AND2x2_ASAP7_75t_L g4493 ( 
.A(n_4285),
.B(n_3959),
.Y(n_4493)
);

INVx4_ASAP7_75t_L g4494 ( 
.A(n_4112),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4237),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_4204),
.B(n_4208),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_SL g4497 ( 
.A(n_4152),
.B(n_3869),
.Y(n_4497)
);

HB1xp67_ASAP7_75t_L g4498 ( 
.A(n_4221),
.Y(n_4498)
);

NAND3xp33_ASAP7_75t_L g4499 ( 
.A(n_4147),
.B(n_1204),
.C(n_1203),
.Y(n_4499)
);

O2A1O1Ixp5_ASAP7_75t_SL g4500 ( 
.A1(n_4278),
.A2(n_2464),
.B(n_2471),
.C(n_2463),
.Y(n_4500)
);

BUFx6f_ASAP7_75t_L g4501 ( 
.A(n_4138),
.Y(n_4501)
);

HB1xp67_ASAP7_75t_L g4502 ( 
.A(n_4264),
.Y(n_4502)
);

OR2x2_ASAP7_75t_L g4503 ( 
.A(n_4131),
.B(n_3959),
.Y(n_4503)
);

CKINVDCx20_ASAP7_75t_R g4504 ( 
.A(n_4365),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4132),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4114),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4164),
.Y(n_4507)
);

BUFx6f_ASAP7_75t_L g4508 ( 
.A(n_4138),
.Y(n_4508)
);

AOI21xp5_ASAP7_75t_L g4509 ( 
.A1(n_4117),
.A2(n_4120),
.B(n_4236),
.Y(n_4509)
);

BUFx3_ASAP7_75t_L g4510 ( 
.A(n_4138),
.Y(n_4510)
);

CKINVDCx5p33_ASAP7_75t_R g4511 ( 
.A(n_4107),
.Y(n_4511)
);

OR2x2_ASAP7_75t_SL g4512 ( 
.A(n_4334),
.B(n_4091),
.Y(n_4512)
);

INVx3_ASAP7_75t_L g4513 ( 
.A(n_4242),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4166),
.Y(n_4514)
);

AOI21x1_ASAP7_75t_L g4515 ( 
.A1(n_4351),
.A2(n_3869),
.B(n_3369),
.Y(n_4515)
);

AND2x4_ASAP7_75t_L g4516 ( 
.A(n_4332),
.B(n_3998),
.Y(n_4516)
);

AOI22xp33_ASAP7_75t_L g4517 ( 
.A1(n_4148),
.A2(n_1205),
.B1(n_1211),
.B2(n_1203),
.Y(n_4517)
);

AND2x2_ASAP7_75t_SL g4518 ( 
.A(n_4282),
.B(n_4091),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4227),
.Y(n_4519)
);

OAI21x1_ASAP7_75t_L g4520 ( 
.A1(n_4157),
.A2(n_2473),
.B(n_2471),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4271),
.Y(n_4521)
);

OAI22xp5_ASAP7_75t_L g4522 ( 
.A1(n_4139),
.A2(n_4093),
.B1(n_4079),
.B2(n_3992),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_4324),
.Y(n_4523)
);

AOI21xp5_ASAP7_75t_L g4524 ( 
.A1(n_4124),
.A2(n_3404),
.B(n_3869),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_4134),
.B(n_3964),
.Y(n_4525)
);

INVx4_ASAP7_75t_L g4526 ( 
.A(n_4141),
.Y(n_4526)
);

NOR2x1_ASAP7_75t_SL g4527 ( 
.A(n_4332),
.B(n_4345),
.Y(n_4527)
);

OR2x2_ASAP7_75t_L g4528 ( 
.A(n_4262),
.B(n_3964),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4128),
.Y(n_4529)
);

OR2x6_ASAP7_75t_L g4530 ( 
.A(n_4323),
.B(n_4093),
.Y(n_4530)
);

CKINVDCx11_ASAP7_75t_R g4531 ( 
.A(n_4141),
.Y(n_4531)
);

AND2x4_ASAP7_75t_L g4532 ( 
.A(n_4340),
.B(n_4079),
.Y(n_4532)
);

BUFx6f_ASAP7_75t_SL g4533 ( 
.A(n_4254),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_4330),
.Y(n_4534)
);

CKINVDCx5p33_ASAP7_75t_R g4535 ( 
.A(n_4106),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4238),
.Y(n_4536)
);

INVx2_ASAP7_75t_SL g4537 ( 
.A(n_4141),
.Y(n_4537)
);

AOI21xp5_ASAP7_75t_L g4538 ( 
.A1(n_4174),
.A2(n_3404),
.B(n_3869),
.Y(n_4538)
);

BUFx6f_ASAP7_75t_L g4539 ( 
.A(n_4146),
.Y(n_4539)
);

BUFx6f_ASAP7_75t_L g4540 ( 
.A(n_4146),
.Y(n_4540)
);

OAI22xp5_ASAP7_75t_L g4541 ( 
.A1(n_4184),
.A2(n_4093),
.B1(n_3992),
.B2(n_4023),
.Y(n_4541)
);

BUFx2_ASAP7_75t_L g4542 ( 
.A(n_4326),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4235),
.Y(n_4543)
);

OR2x6_ASAP7_75t_L g4544 ( 
.A(n_4355),
.B(n_3964),
.Y(n_4544)
);

AOI21xp5_ASAP7_75t_L g4545 ( 
.A1(n_4210),
.A2(n_3040),
.B(n_3992),
.Y(n_4545)
);

BUFx2_ASAP7_75t_L g4546 ( 
.A(n_4310),
.Y(n_4546)
);

BUFx6f_ASAP7_75t_L g4547 ( 
.A(n_4146),
.Y(n_4547)
);

HB1xp67_ASAP7_75t_L g4548 ( 
.A(n_4241),
.Y(n_4548)
);

AOI21xp33_ASAP7_75t_L g4549 ( 
.A1(n_4144),
.A2(n_4037),
.B(n_4023),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4315),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4327),
.Y(n_4551)
);

INVx3_ASAP7_75t_L g4552 ( 
.A(n_4209),
.Y(n_4552)
);

INVx2_ASAP7_75t_L g4553 ( 
.A(n_4370),
.Y(n_4553)
);

BUFx6f_ASAP7_75t_L g4554 ( 
.A(n_4209),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4328),
.Y(n_4555)
);

AND2x4_ASAP7_75t_L g4556 ( 
.A(n_4357),
.B(n_4023),
.Y(n_4556)
);

INVx1_ASAP7_75t_SL g4557 ( 
.A(n_4216),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4244),
.B(n_4037),
.Y(n_4558)
);

HB1xp67_ASAP7_75t_L g4559 ( 
.A(n_4292),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4346),
.Y(n_4560)
);

INVx3_ASAP7_75t_L g4561 ( 
.A(n_4209),
.Y(n_4561)
);

OAI22xp5_ASAP7_75t_L g4562 ( 
.A1(n_4119),
.A2(n_4274),
.B1(n_4125),
.B2(n_4263),
.Y(n_4562)
);

CKINVDCx5p33_ASAP7_75t_R g4563 ( 
.A(n_4350),
.Y(n_4563)
);

INVx6_ASAP7_75t_SL g4564 ( 
.A(n_4344),
.Y(n_4564)
);

INVx4_ASAP7_75t_L g4565 ( 
.A(n_4229),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4352),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4229),
.Y(n_4567)
);

BUFx3_ASAP7_75t_L g4568 ( 
.A(n_4229),
.Y(n_4568)
);

AOI22xp33_ASAP7_75t_L g4569 ( 
.A1(n_4178),
.A2(n_1208),
.B1(n_1214),
.B2(n_1205),
.Y(n_4569)
);

BUFx3_ASAP7_75t_L g4570 ( 
.A(n_4247),
.Y(n_4570)
);

AOI221xp5_ASAP7_75t_L g4571 ( 
.A1(n_4276),
.A2(n_1057),
.B1(n_1058),
.B2(n_1056),
.C(n_1054),
.Y(n_4571)
);

HAxp5_ASAP7_75t_L g4572 ( 
.A(n_4215),
.B(n_1208),
.CON(n_4572),
.SN(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_4135),
.A2(n_3040),
.B(n_4037),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4253),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4233),
.Y(n_4575)
);

AOI21xp5_ASAP7_75t_L g4576 ( 
.A1(n_4298),
.A2(n_4300),
.B(n_4190),
.Y(n_4576)
);

OAI22xp5_ASAP7_75t_L g4577 ( 
.A1(n_4180),
.A2(n_4055),
.B1(n_4069),
.B2(n_4043),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4188),
.Y(n_4578)
);

BUFx6f_ASAP7_75t_L g4579 ( 
.A(n_4247),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_4160),
.B(n_4043),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4364),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4247),
.Y(n_4582)
);

OAI21x1_ASAP7_75t_L g4583 ( 
.A1(n_4331),
.A2(n_2473),
.B(n_2423),
.Y(n_4583)
);

INVx3_ASAP7_75t_L g4584 ( 
.A(n_4268),
.Y(n_4584)
);

BUFx3_ASAP7_75t_L g4585 ( 
.A(n_4268),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4367),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4230),
.Y(n_4587)
);

INVx2_ASAP7_75t_L g4588 ( 
.A(n_4268),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4265),
.Y(n_4589)
);

INVx2_ASAP7_75t_SL g4590 ( 
.A(n_4322),
.Y(n_4590)
);

CKINVDCx20_ASAP7_75t_R g4591 ( 
.A(n_4257),
.Y(n_4591)
);

BUFx6f_ASAP7_75t_L g4592 ( 
.A(n_4322),
.Y(n_4592)
);

BUFx6f_ASAP7_75t_L g4593 ( 
.A(n_4322),
.Y(n_4593)
);

CKINVDCx11_ASAP7_75t_R g4594 ( 
.A(n_4359),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4288),
.Y(n_4595)
);

INVx3_ASAP7_75t_L g4596 ( 
.A(n_4168),
.Y(n_4596)
);

INVx2_ASAP7_75t_SL g4597 ( 
.A(n_4225),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4354),
.B(n_4043),
.Y(n_4598)
);

NAND2xp33_ASAP7_75t_L g4599 ( 
.A(n_4275),
.B(n_4309),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4201),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4214),
.B(n_4055),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4255),
.B(n_4055),
.Y(n_4602)
);

AOI22xp5_ASAP7_75t_L g4603 ( 
.A1(n_4181),
.A2(n_1062),
.B1(n_1063),
.B2(n_1059),
.Y(n_4603)
);

NAND2xp5_ASAP7_75t_SL g4604 ( 
.A(n_4280),
.B(n_4069),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4289),
.Y(n_4605)
);

OAI22xp5_ASAP7_75t_L g4606 ( 
.A1(n_4251),
.A2(n_4072),
.B1(n_4074),
.B2(n_4069),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4295),
.Y(n_4607)
);

INVxp67_ASAP7_75t_L g4608 ( 
.A(n_4240),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4297),
.Y(n_4609)
);

INVx3_ASAP7_75t_SL g4610 ( 
.A(n_4248),
.Y(n_4610)
);

BUFx3_ASAP7_75t_L g4611 ( 
.A(n_4360),
.Y(n_4611)
);

A2O1A1Ixp33_ASAP7_75t_L g4612 ( 
.A1(n_4172),
.A2(n_1214),
.B(n_1217),
.C(n_1211),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4301),
.Y(n_4613)
);

BUFx3_ASAP7_75t_L g4614 ( 
.A(n_4303),
.Y(n_4614)
);

AOI22xp33_ASAP7_75t_L g4615 ( 
.A1(n_4195),
.A2(n_1219),
.B1(n_1221),
.B2(n_1217),
.Y(n_4615)
);

OAI22xp33_ASAP7_75t_SL g4616 ( 
.A1(n_4213),
.A2(n_4122),
.B1(n_1219),
.B2(n_1221),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4306),
.Y(n_4617)
);

BUFx3_ASAP7_75t_L g4618 ( 
.A(n_4307),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_4342),
.B(n_4072),
.Y(n_4619)
);

INVxp67_ASAP7_75t_SL g4620 ( 
.A(n_4296),
.Y(n_4620)
);

OAI22xp5_ASAP7_75t_L g4621 ( 
.A1(n_4305),
.A2(n_4074),
.B1(n_4076),
.B2(n_4072),
.Y(n_4621)
);

BUFx3_ASAP7_75t_L g4622 ( 
.A(n_4348),
.Y(n_4622)
);

INVx8_ASAP7_75t_L g4623 ( 
.A(n_4234),
.Y(n_4623)
);

INVx6_ASAP7_75t_SL g4624 ( 
.A(n_4283),
.Y(n_4624)
);

INVx4_ASAP7_75t_L g4625 ( 
.A(n_4316),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4356),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4206),
.Y(n_4627)
);

OR2x6_ASAP7_75t_SL g4628 ( 
.A(n_4261),
.B(n_1218),
.Y(n_4628)
);

NOR2xp67_ASAP7_75t_L g4629 ( 
.A(n_4336),
.B(n_4339),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4200),
.B(n_4074),
.Y(n_4630)
);

OAI22xp5_ASAP7_75t_SL g4631 ( 
.A1(n_4207),
.A2(n_1226),
.B1(n_1227),
.B2(n_1218),
.Y(n_4631)
);

HB1xp67_ASAP7_75t_L g4632 ( 
.A(n_4217),
.Y(n_4632)
);

NOR2xp67_ASAP7_75t_SL g4633 ( 
.A(n_4267),
.B(n_4076),
.Y(n_4633)
);

HB1xp67_ASAP7_75t_L g4634 ( 
.A(n_4223),
.Y(n_4634)
);

BUFx6f_ASAP7_75t_L g4635 ( 
.A(n_4320),
.Y(n_4635)
);

INVx4_ASAP7_75t_L g4636 ( 
.A(n_4321),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4239),
.B(n_4076),
.Y(n_4637)
);

INVx4_ASAP7_75t_L g4638 ( 
.A(n_4335),
.Y(n_4638)
);

O2A1O1Ixp33_ASAP7_75t_L g4639 ( 
.A1(n_4562),
.A2(n_4243),
.B(n_4273),
.C(n_4211),
.Y(n_4639)
);

A2O1A1Ixp33_ASAP7_75t_L g4640 ( 
.A1(n_4499),
.A2(n_4149),
.B(n_4314),
.C(n_4338),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4451),
.Y(n_4641)
);

OR2x2_ASAP7_75t_L g4642 ( 
.A(n_4380),
.B(n_4249),
.Y(n_4642)
);

AOI21xp5_ASAP7_75t_L g4643 ( 
.A1(n_4576),
.A2(n_4290),
.B(n_4293),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4449),
.B(n_4186),
.Y(n_4644)
);

INVx2_ASAP7_75t_SL g4645 ( 
.A(n_4417),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4491),
.Y(n_4646)
);

NAND2xp5_ASAP7_75t_L g4647 ( 
.A(n_4457),
.B(n_1065),
.Y(n_4647)
);

INVx2_ASAP7_75t_SL g4648 ( 
.A(n_4417),
.Y(n_4648)
);

O2A1O1Ixp33_ASAP7_75t_SL g4649 ( 
.A1(n_4398),
.A2(n_4347),
.B(n_4366),
.C(n_4349),
.Y(n_4649)
);

AOI21xp5_ASAP7_75t_L g4650 ( 
.A1(n_4509),
.A2(n_4270),
.B(n_4279),
.Y(n_4650)
);

A2O1A1Ixp33_ASAP7_75t_L g4651 ( 
.A1(n_4382),
.A2(n_4368),
.B(n_4362),
.C(n_1241),
.Y(n_4651)
);

INVx5_ASAP7_75t_L g4652 ( 
.A(n_4482),
.Y(n_4652)
);

AOI221xp5_ASAP7_75t_SL g4653 ( 
.A1(n_4631),
.A2(n_1227),
.B1(n_1228),
.B2(n_1226),
.C(n_1222),
.Y(n_4653)
);

AO31x2_ASAP7_75t_L g4654 ( 
.A1(n_4506),
.A2(n_3367),
.A3(n_3179),
.B(n_3064),
.Y(n_4654)
);

AO31x2_ASAP7_75t_L g4655 ( 
.A1(n_4542),
.A2(n_3179),
.A3(n_3064),
.B(n_2142),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4491),
.Y(n_4656)
);

BUFx2_ASAP7_75t_L g4657 ( 
.A(n_4502),
.Y(n_4657)
);

NOR2xp33_ASAP7_75t_L g4658 ( 
.A(n_4557),
.B(n_1066),
.Y(n_4658)
);

OAI21x1_ASAP7_75t_L g4659 ( 
.A1(n_4520),
.A2(n_2473),
.B(n_2423),
.Y(n_4659)
);

O2A1O1Ixp33_ASAP7_75t_SL g4660 ( 
.A1(n_4578),
.A2(n_13),
.B(n_24),
.C(n_5),
.Y(n_4660)
);

AOI21xp5_ASAP7_75t_L g4661 ( 
.A1(n_4599),
.A2(n_4620),
.B(n_4418),
.Y(n_4661)
);

BUFx12f_ASAP7_75t_L g4662 ( 
.A(n_4511),
.Y(n_4662)
);

BUFx8_ASAP7_75t_SL g4663 ( 
.A(n_4504),
.Y(n_4663)
);

NAND2x1p5_ASAP7_75t_L g4664 ( 
.A(n_4431),
.B(n_2528),
.Y(n_4664)
);

A2O1A1Ixp33_ASAP7_75t_L g4665 ( 
.A1(n_4394),
.A2(n_1255),
.B(n_1273),
.C(n_1238),
.Y(n_4665)
);

BUFx12f_ASAP7_75t_L g4666 ( 
.A(n_4406),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4393),
.Y(n_4667)
);

NOR2xp33_ASAP7_75t_SL g4668 ( 
.A(n_4447),
.B(n_1222),
.Y(n_4668)
);

INVx3_ASAP7_75t_L g4669 ( 
.A(n_4378),
.Y(n_4669)
);

O2A1O1Ixp33_ASAP7_75t_SL g4670 ( 
.A1(n_4497),
.A2(n_15),
.B(n_26),
.C(n_5),
.Y(n_4670)
);

A2O1A1Ixp33_ASAP7_75t_L g4671 ( 
.A1(n_4529),
.A2(n_1263),
.B(n_1280),
.C(n_1240),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4455),
.Y(n_4672)
);

HB1xp67_ASAP7_75t_L g4673 ( 
.A(n_4443),
.Y(n_4673)
);

NAND2xp33_ASAP7_75t_L g4674 ( 
.A(n_4615),
.B(n_1228),
.Y(n_4674)
);

OR2x2_ASAP7_75t_L g4675 ( 
.A(n_4498),
.B(n_2017),
.Y(n_4675)
);

OAI21x1_ASAP7_75t_L g4676 ( 
.A1(n_4524),
.A2(n_2483),
.B(n_2184),
.Y(n_4676)
);

OAI22xp5_ASAP7_75t_L g4677 ( 
.A1(n_4628),
.A2(n_1236),
.B1(n_1237),
.B2(n_1235),
.Y(n_4677)
);

INVx1_ASAP7_75t_SL g4678 ( 
.A(n_4548),
.Y(n_4678)
);

OAI21xp5_ASAP7_75t_L g4679 ( 
.A1(n_4603),
.A2(n_1236),
.B(n_1235),
.Y(n_4679)
);

BUFx3_ASAP7_75t_L g4680 ( 
.A(n_4378),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4536),
.B(n_1067),
.Y(n_4681)
);

A2O1A1Ixp33_ASAP7_75t_L g4682 ( 
.A1(n_4612),
.A2(n_1269),
.B(n_1286),
.C(n_1247),
.Y(n_4682)
);

AO221x2_ASAP7_75t_L g4683 ( 
.A1(n_4587),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_4683)
);

AOI221xp5_ASAP7_75t_L g4684 ( 
.A1(n_4569),
.A2(n_1239),
.B1(n_1240),
.B2(n_1238),
.C(n_1237),
.Y(n_4684)
);

O2A1O1Ixp33_ASAP7_75t_L g4685 ( 
.A1(n_4375),
.A2(n_1244),
.B(n_1245),
.C(n_1239),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4496),
.B(n_1068),
.Y(n_4686)
);

A2O1A1Ixp33_ASAP7_75t_L g4687 ( 
.A1(n_4634),
.A2(n_1268),
.B(n_1285),
.C(n_1245),
.Y(n_4687)
);

AO21x2_ASAP7_75t_L g4688 ( 
.A1(n_4574),
.A2(n_3179),
.B(n_3064),
.Y(n_4688)
);

AO31x2_ASAP7_75t_L g4689 ( 
.A1(n_4542),
.A2(n_3179),
.A3(n_3064),
.B(n_2142),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4402),
.Y(n_4690)
);

INVx2_ASAP7_75t_SL g4691 ( 
.A(n_4378),
.Y(n_4691)
);

OAI21x1_ASAP7_75t_SL g4692 ( 
.A1(n_4527),
.A2(n_7),
.B(n_8),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4507),
.B(n_1071),
.Y(n_4693)
);

INVx5_ASAP7_75t_L g4694 ( 
.A(n_4482),
.Y(n_4694)
);

OAI21xp5_ASAP7_75t_L g4695 ( 
.A1(n_4444),
.A2(n_1244),
.B(n_1241),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4514),
.B(n_1074),
.Y(n_4696)
);

O2A1O1Ixp33_ASAP7_75t_L g4697 ( 
.A1(n_4616),
.A2(n_1251),
.B(n_1255),
.C(n_1247),
.Y(n_4697)
);

A2O1A1Ixp33_ASAP7_75t_L g4698 ( 
.A1(n_4389),
.A2(n_1286),
.B(n_1269),
.C(n_1261),
.Y(n_4698)
);

OAI21x1_ASAP7_75t_L g4699 ( 
.A1(n_4515),
.A2(n_2483),
.B(n_2184),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4403),
.Y(n_4700)
);

A2O1A1Ixp33_ASAP7_75t_L g4701 ( 
.A1(n_4413),
.A2(n_1270),
.B(n_1261),
.C(n_1263),
.Y(n_4701)
);

AO31x2_ASAP7_75t_L g4702 ( 
.A1(n_4546),
.A2(n_2142),
.A3(n_2263),
.B(n_2123),
.Y(n_4702)
);

OR2x2_ASAP7_75t_L g4703 ( 
.A(n_4400),
.B(n_2017),
.Y(n_4703)
);

NOR2x1_ASAP7_75t_SL g4704 ( 
.A(n_4372),
.B(n_2021),
.Y(n_4704)
);

CKINVDCx11_ASAP7_75t_R g4705 ( 
.A(n_4401),
.Y(n_4705)
);

NOR2xp67_ASAP7_75t_L g4706 ( 
.A(n_4424),
.B(n_10),
.Y(n_4706)
);

CKINVDCx20_ASAP7_75t_R g4707 ( 
.A(n_4591),
.Y(n_4707)
);

AOI21xp5_ASAP7_75t_L g4708 ( 
.A1(n_4430),
.A2(n_2535),
.B(n_2528),
.Y(n_4708)
);

BUFx4f_ASAP7_75t_SL g4709 ( 
.A(n_4467),
.Y(n_4709)
);

AOI21xp5_ASAP7_75t_L g4710 ( 
.A1(n_4538),
.A2(n_4573),
.B(n_4580),
.Y(n_4710)
);

INVx4_ASAP7_75t_L g4711 ( 
.A(n_4531),
.Y(n_4711)
);

AOI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4428),
.A2(n_2535),
.B(n_2528),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4404),
.Y(n_4713)
);

OAI21x1_ASAP7_75t_L g4714 ( 
.A1(n_4515),
.A2(n_2023),
.B(n_2021),
.Y(n_4714)
);

INVx3_ASAP7_75t_L g4715 ( 
.A(n_4440),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_SL g4716 ( 
.A(n_4384),
.B(n_2021),
.Y(n_4716)
);

BUFx2_ASAP7_75t_L g4717 ( 
.A(n_4376),
.Y(n_4717)
);

AOI22xp33_ASAP7_75t_L g4718 ( 
.A1(n_4632),
.A2(n_1264),
.B1(n_1266),
.B2(n_1251),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4408),
.Y(n_4719)
);

BUFx3_ASAP7_75t_L g4720 ( 
.A(n_4454),
.Y(n_4720)
);

AOI22xp33_ASAP7_75t_L g4721 ( 
.A1(n_4575),
.A2(n_1266),
.B1(n_1268),
.B2(n_1264),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4409),
.Y(n_4722)
);

INVx4_ASAP7_75t_L g4723 ( 
.A(n_4429),
.Y(n_4723)
);

AOI21xp5_ASAP7_75t_L g4724 ( 
.A1(n_4545),
.A2(n_2540),
.B(n_2492),
.Y(n_4724)
);

NOR2xp33_ASAP7_75t_L g4725 ( 
.A(n_4399),
.B(n_1077),
.Y(n_4725)
);

OAI21x1_ASAP7_75t_L g4726 ( 
.A1(n_4583),
.A2(n_2023),
.B(n_2021),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4419),
.Y(n_4727)
);

OAI22xp5_ASAP7_75t_L g4728 ( 
.A1(n_4379),
.A2(n_4512),
.B1(n_4518),
.B2(n_4517),
.Y(n_4728)
);

OAI21x1_ASAP7_75t_L g4729 ( 
.A1(n_4500),
.A2(n_2044),
.B(n_2023),
.Y(n_4729)
);

AO31x2_ASAP7_75t_L g4730 ( 
.A1(n_4546),
.A2(n_2263),
.A3(n_2441),
.B(n_2123),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4505),
.B(n_1081),
.Y(n_4731)
);

AO32x2_ASAP7_75t_L g4732 ( 
.A1(n_4416),
.A2(n_1276),
.A3(n_1280),
.B1(n_1273),
.B2(n_1270),
.Y(n_4732)
);

INVxp67_ASAP7_75t_L g4733 ( 
.A(n_4433),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4421),
.Y(n_4734)
);

O2A1O1Ixp33_ASAP7_75t_L g4735 ( 
.A1(n_4461),
.A2(n_4445),
.B(n_4572),
.C(n_4581),
.Y(n_4735)
);

AO32x2_ASAP7_75t_L g4736 ( 
.A1(n_4487),
.A2(n_1284),
.A3(n_1285),
.B1(n_1282),
.B2(n_1276),
.Y(n_4736)
);

NOR4xp25_ASAP7_75t_L g4737 ( 
.A(n_4627),
.B(n_1284),
.C(n_1287),
.D(n_1282),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4425),
.Y(n_4738)
);

BUFx12f_ASAP7_75t_L g4739 ( 
.A(n_4535),
.Y(n_4739)
);

INVx2_ASAP7_75t_SL g4740 ( 
.A(n_4439),
.Y(n_4740)
);

AOI21xp5_ASAP7_75t_L g4741 ( 
.A1(n_4435),
.A2(n_2540),
.B(n_2492),
.Y(n_4741)
);

O2A1O1Ixp33_ASAP7_75t_L g4742 ( 
.A1(n_4586),
.A2(n_1287),
.B(n_1091),
.C(n_1092),
.Y(n_4742)
);

INVx2_ASAP7_75t_L g4743 ( 
.A(n_4478),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4381),
.B(n_1084),
.Y(n_4744)
);

BUFx10_ASAP7_75t_L g4745 ( 
.A(n_4377),
.Y(n_4745)
);

OAI22xp5_ASAP7_75t_L g4746 ( 
.A1(n_4618),
.A2(n_4622),
.B1(n_4608),
.B2(n_4426),
.Y(n_4746)
);

OAI21x1_ASAP7_75t_L g4747 ( 
.A1(n_4453),
.A2(n_2044),
.B(n_2023),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4436),
.Y(n_4748)
);

AOI21xp5_ASAP7_75t_L g4749 ( 
.A1(n_4471),
.A2(n_2540),
.B(n_2492),
.Y(n_4749)
);

AO31x2_ASAP7_75t_L g4750 ( 
.A1(n_4371),
.A2(n_2263),
.A3(n_2441),
.B(n_2123),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4473),
.B(n_11),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4519),
.B(n_1100),
.Y(n_4752)
);

AOI221x1_ASAP7_75t_L g4753 ( 
.A1(n_4549),
.A2(n_2058),
.B1(n_2069),
.B2(n_2049),
.C(n_2044),
.Y(n_4753)
);

AOI22xp5_ASAP7_75t_L g4754 ( 
.A1(n_4390),
.A2(n_1107),
.B1(n_1109),
.B2(n_1104),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4459),
.Y(n_4755)
);

INVx3_ASAP7_75t_L g4756 ( 
.A(n_4494),
.Y(n_4756)
);

BUFx2_ASAP7_75t_L g4757 ( 
.A(n_4376),
.Y(n_4757)
);

NOR2xp67_ASAP7_75t_L g4758 ( 
.A(n_4420),
.B(n_11),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4460),
.Y(n_4759)
);

AOI221xp5_ASAP7_75t_L g4760 ( 
.A1(n_4571),
.A2(n_1118),
.B1(n_1121),
.B2(n_1117),
.C(n_1111),
.Y(n_4760)
);

O2A1O1Ixp33_ASAP7_75t_SL g4761 ( 
.A1(n_4522),
.A2(n_25),
.B(n_33),
.C(n_12),
.Y(n_4761)
);

AO31x2_ASAP7_75t_L g4762 ( 
.A1(n_4371),
.A2(n_2509),
.A3(n_2441),
.B(n_16),
.Y(n_4762)
);

INVx2_ASAP7_75t_L g4763 ( 
.A(n_4489),
.Y(n_4763)
);

AOI22xp33_ASAP7_75t_L g4764 ( 
.A1(n_4469),
.A2(n_4543),
.B1(n_4595),
.B2(n_4589),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4386),
.B(n_1122),
.Y(n_4765)
);

OAI21x1_ASAP7_75t_L g4766 ( 
.A1(n_4630),
.A2(n_2049),
.B(n_2044),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_SL g4767 ( 
.A(n_4495),
.B(n_2049),
.Y(n_4767)
);

NAND2x1_ASAP7_75t_L g4768 ( 
.A(n_4372),
.B(n_2049),
.Y(n_4768)
);

O2A1O1Ixp33_ASAP7_75t_SL g4769 ( 
.A1(n_4601),
.A2(n_26),
.B(n_34),
.C(n_12),
.Y(n_4769)
);

AO31x2_ASAP7_75t_L g4770 ( 
.A1(n_4374),
.A2(n_2509),
.A3(n_19),
.B(n_15),
.Y(n_4770)
);

OAI21xp5_ASAP7_75t_L g4771 ( 
.A1(n_4477),
.A2(n_1124),
.B(n_1123),
.Y(n_4771)
);

OAI211xp5_ASAP7_75t_L g4772 ( 
.A1(n_4486),
.A2(n_1131),
.B(n_1132),
.C(n_1125),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4466),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4475),
.Y(n_4774)
);

AOI21xp5_ASAP7_75t_L g4775 ( 
.A1(n_4431),
.A2(n_2540),
.B(n_2202),
.Y(n_4775)
);

OAI21xp5_ASAP7_75t_L g4776 ( 
.A1(n_4476),
.A2(n_1137),
.B(n_1133),
.Y(n_4776)
);

OAI22xp5_ASAP7_75t_L g4777 ( 
.A1(n_4598),
.A2(n_1143),
.B1(n_1140),
.B2(n_2058),
.Y(n_4777)
);

HB1xp67_ASAP7_75t_L g4778 ( 
.A(n_4559),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4373),
.Y(n_4779)
);

INVx3_ASAP7_75t_L g4780 ( 
.A(n_4526),
.Y(n_4780)
);

A2O1A1Ixp33_ASAP7_75t_L g4781 ( 
.A1(n_4605),
.A2(n_2069),
.B(n_2077),
.C(n_2058),
.Y(n_4781)
);

A2O1A1Ixp33_ASAP7_75t_L g4782 ( 
.A1(n_4607),
.A2(n_2069),
.B(n_2077),
.C(n_2058),
.Y(n_4782)
);

AOI22xp5_ASAP7_75t_L g4783 ( 
.A1(n_4609),
.A2(n_4617),
.B1(n_4626),
.B2(n_4613),
.Y(n_4783)
);

BUFx2_ASAP7_75t_L g4784 ( 
.A(n_4465),
.Y(n_4784)
);

HB1xp67_ASAP7_75t_L g4785 ( 
.A(n_4637),
.Y(n_4785)
);

AND2x4_ASAP7_75t_L g4786 ( 
.A(n_4493),
.B(n_636),
.Y(n_4786)
);

INVx2_ASAP7_75t_L g4787 ( 
.A(n_4385),
.Y(n_4787)
);

AO31x2_ASAP7_75t_L g4788 ( 
.A1(n_4374),
.A2(n_2509),
.A3(n_20),
.B(n_17),
.Y(n_4788)
);

OAI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4604),
.A2(n_1921),
.B(n_1900),
.Y(n_4789)
);

AOI221xp5_ASAP7_75t_SL g4790 ( 
.A1(n_4481),
.A2(n_2085),
.B1(n_2089),
.B2(n_2077),
.C(n_2069),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4383),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4383),
.Y(n_4792)
);

BUFx3_ASAP7_75t_L g4793 ( 
.A(n_4410),
.Y(n_4793)
);

CKINVDCx5p33_ASAP7_75t_R g4794 ( 
.A(n_4563),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4395),
.Y(n_4795)
);

BUFx8_ASAP7_75t_L g4796 ( 
.A(n_4533),
.Y(n_4796)
);

OAI21xp5_ASAP7_75t_L g4797 ( 
.A1(n_4629),
.A2(n_1921),
.B(n_1900),
.Y(n_4797)
);

AOI21xp5_ASAP7_75t_L g4798 ( 
.A1(n_4431),
.A2(n_2202),
.B(n_2189),
.Y(n_4798)
);

AOI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4488),
.A2(n_2202),
.B(n_2189),
.Y(n_4799)
);

INVx3_ASAP7_75t_L g4800 ( 
.A(n_4565),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4438),
.B(n_2077),
.Y(n_4801)
);

AOI21x1_ASAP7_75t_L g4802 ( 
.A1(n_4633),
.A2(n_2089),
.B(n_2085),
.Y(n_4802)
);

AOI22xp33_ASAP7_75t_L g4803 ( 
.A1(n_4521),
.A2(n_2089),
.B1(n_2093),
.B2(n_2085),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4395),
.Y(n_4804)
);

AOI21xp5_ASAP7_75t_L g4805 ( 
.A1(n_4392),
.A2(n_2202),
.B(n_2189),
.Y(n_4805)
);

O2A1O1Ixp33_ASAP7_75t_L g4806 ( 
.A1(n_4577),
.A2(n_22),
.B(n_17),
.C(n_19),
.Y(n_4806)
);

OAI21x1_ASAP7_75t_L g4807 ( 
.A1(n_4550),
.A2(n_2089),
.B(n_2085),
.Y(n_4807)
);

A2O1A1Ixp33_ASAP7_75t_L g4808 ( 
.A1(n_4405),
.A2(n_2114),
.B(n_2093),
.C(n_25),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4387),
.Y(n_4809)
);

AOI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4625),
.A2(n_2206),
.B(n_2189),
.Y(n_4810)
);

OAI21xp5_ASAP7_75t_L g4811 ( 
.A1(n_4621),
.A2(n_1921),
.B(n_1900),
.Y(n_4811)
);

INVx3_ASAP7_75t_L g4812 ( 
.A(n_4429),
.Y(n_4812)
);

AOI22xp33_ASAP7_75t_SL g4813 ( 
.A1(n_4405),
.A2(n_2114),
.B1(n_2093),
.B2(n_27),
.Y(n_4813)
);

HB1xp67_ASAP7_75t_L g4814 ( 
.A(n_4503),
.Y(n_4814)
);

AOI22xp5_ASAP7_75t_L g4815 ( 
.A1(n_4423),
.A2(n_4534),
.B1(n_4523),
.B2(n_4490),
.Y(n_4815)
);

O2A1O1Ixp33_ASAP7_75t_L g4816 ( 
.A1(n_4558),
.A2(n_28),
.B(n_22),
.C(n_23),
.Y(n_4816)
);

OAI22xp5_ASAP7_75t_L g4817 ( 
.A1(n_4624),
.A2(n_2114),
.B1(n_2093),
.B2(n_2206),
.Y(n_4817)
);

INVx1_ASAP7_75t_L g4818 ( 
.A(n_4388),
.Y(n_4818)
);

OAI21xp5_ASAP7_75t_L g4819 ( 
.A1(n_4606),
.A2(n_1921),
.B(n_1900),
.Y(n_4819)
);

A2O1A1Ixp33_ASAP7_75t_L g4820 ( 
.A1(n_4415),
.A2(n_2114),
.B(n_30),
.C(n_28),
.Y(n_4820)
);

O2A1O1Ixp33_ASAP7_75t_L g4821 ( 
.A1(n_4619),
.A2(n_32),
.B(n_29),
.C(n_31),
.Y(n_4821)
);

O2A1O1Ixp33_ASAP7_75t_SL g4822 ( 
.A1(n_4525),
.A2(n_4597),
.B(n_4470),
.C(n_4602),
.Y(n_4822)
);

OAI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_4624),
.A2(n_2215),
.B1(n_2230),
.B2(n_2206),
.Y(n_4823)
);

AO31x2_ASAP7_75t_L g4824 ( 
.A1(n_4415),
.A2(n_33),
.A3(n_31),
.B(n_32),
.Y(n_4824)
);

AOI22xp5_ASAP7_75t_L g4825 ( 
.A1(n_4423),
.A2(n_4490),
.B1(n_4432),
.B2(n_4636),
.Y(n_4825)
);

AND2x2_ASAP7_75t_L g4826 ( 
.A(n_4411),
.B(n_34),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4391),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_4472),
.B(n_4479),
.Y(n_4828)
);

BUFx2_ASAP7_75t_L g4829 ( 
.A(n_4492),
.Y(n_4829)
);

O2A1O1Ixp33_ASAP7_75t_SL g4830 ( 
.A1(n_4485),
.A2(n_47),
.B(n_58),
.C(n_35),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4483),
.B(n_35),
.Y(n_4831)
);

AOI21xp5_ASAP7_75t_L g4832 ( 
.A1(n_4437),
.A2(n_2215),
.B(n_2206),
.Y(n_4832)
);

AOI22xp5_ASAP7_75t_L g4833 ( 
.A1(n_4437),
.A2(n_1924),
.B1(n_2230),
.B2(n_2215),
.Y(n_4833)
);

OR2x6_ASAP7_75t_L g4834 ( 
.A(n_4450),
.B(n_2215),
.Y(n_4834)
);

AOI22xp33_ASAP7_75t_L g4835 ( 
.A1(n_4553),
.A2(n_1924),
.B1(n_2239),
.B2(n_2230),
.Y(n_4835)
);

AOI21xp5_ASAP7_75t_L g4836 ( 
.A1(n_4450),
.A2(n_2239),
.B(n_2230),
.Y(n_4836)
);

OAI21x1_ASAP7_75t_L g4837 ( 
.A1(n_4551),
.A2(n_4560),
.B(n_4555),
.Y(n_4837)
);

NOR2x1_ASAP7_75t_SL g4838 ( 
.A(n_4530),
.B(n_2239),
.Y(n_4838)
);

OAI21x1_ASAP7_75t_L g4839 ( 
.A1(n_4566),
.A2(n_640),
.B(n_637),
.Y(n_4839)
);

NAND2xp33_ASAP7_75t_SL g4840 ( 
.A(n_4610),
.B(n_36),
.Y(n_4840)
);

AOI21xp5_ASAP7_75t_L g4841 ( 
.A1(n_4638),
.A2(n_2243),
.B(n_2239),
.Y(n_4841)
);

BUFx4f_ASAP7_75t_L g4842 ( 
.A(n_4623),
.Y(n_4842)
);

AOI221xp5_ASAP7_75t_L g4843 ( 
.A1(n_4480),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.C(n_41),
.Y(n_4843)
);

INVx3_ASAP7_75t_SL g4844 ( 
.A(n_4623),
.Y(n_4844)
);

AOI22xp5_ASAP7_75t_L g4845 ( 
.A1(n_4442),
.A2(n_1924),
.B1(n_2247),
.B2(n_2243),
.Y(n_4845)
);

A2O1A1Ixp33_ASAP7_75t_L g4846 ( 
.A1(n_4480),
.A2(n_45),
.B(n_39),
.C(n_42),
.Y(n_4846)
);

AOI22xp33_ASAP7_75t_L g4847 ( 
.A1(n_4528),
.A2(n_1924),
.B1(n_2247),
.B2(n_2243),
.Y(n_4847)
);

O2A1O1Ixp33_ASAP7_75t_SL g4848 ( 
.A1(n_4468),
.A2(n_55),
.B(n_67),
.C(n_42),
.Y(n_4848)
);

AO32x2_ASAP7_75t_L g4849 ( 
.A1(n_4541),
.A2(n_48),
.A3(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_4849)
);

A2O1A1Ixp33_ASAP7_75t_L g4850 ( 
.A1(n_4614),
.A2(n_52),
.B(n_46),
.C(n_50),
.Y(n_4850)
);

INVx2_ASAP7_75t_SL g4851 ( 
.A(n_4458),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4397),
.Y(n_4852)
);

INVx2_ASAP7_75t_SL g4853 ( 
.A(n_4458),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4456),
.B(n_4422),
.Y(n_4854)
);

INVx2_ASAP7_75t_L g4855 ( 
.A(n_4407),
.Y(n_4855)
);

AOI22xp5_ASAP7_75t_L g4856 ( 
.A1(n_4516),
.A2(n_4635),
.B1(n_4513),
.B2(n_4594),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4412),
.B(n_53),
.Y(n_4857)
);

AO32x2_ASAP7_75t_L g4858 ( 
.A1(n_4537),
.A2(n_57),
.A3(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_4858)
);

AND2x4_ASAP7_75t_L g4859 ( 
.A(n_4414),
.B(n_642),
.Y(n_4859)
);

O2A1O1Ixp33_ASAP7_75t_L g4860 ( 
.A1(n_4530),
.A2(n_4600),
.B(n_4532),
.C(n_4463),
.Y(n_4860)
);

O2A1O1Ixp33_ASAP7_75t_SL g4861 ( 
.A1(n_4590),
.A2(n_69),
.B(n_79),
.C(n_54),
.Y(n_4861)
);

NOR2xp33_ASAP7_75t_L g4862 ( 
.A(n_4396),
.B(n_59),
.Y(n_4862)
);

OAI21xp5_ASAP7_75t_L g4863 ( 
.A1(n_4633),
.A2(n_645),
.B(n_644),
.Y(n_4863)
);

AOI21xp5_ASAP7_75t_L g4864 ( 
.A1(n_4635),
.A2(n_2247),
.B(n_2243),
.Y(n_4864)
);

AOI21xp5_ASAP7_75t_L g4865 ( 
.A1(n_4544),
.A2(n_2253),
.B(n_2247),
.Y(n_4865)
);

AOI21xp5_ASAP7_75t_L g4866 ( 
.A1(n_4544),
.A2(n_2276),
.B(n_2253),
.Y(n_4866)
);

INVx1_ASAP7_75t_SL g4867 ( 
.A(n_4510),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_L g4868 ( 
.A(n_4427),
.B(n_61),
.Y(n_4868)
);

AOI22xp5_ASAP7_75t_L g4869 ( 
.A1(n_4516),
.A2(n_2276),
.B1(n_2289),
.B2(n_2253),
.Y(n_4869)
);

INVx2_ASAP7_75t_L g4870 ( 
.A(n_4434),
.Y(n_4870)
);

INVx3_ASAP7_75t_L g4871 ( 
.A(n_4539),
.Y(n_4871)
);

O2A1O1Ixp33_ASAP7_75t_SL g4872 ( 
.A1(n_4596),
.A2(n_71),
.B(n_81),
.C(n_61),
.Y(n_4872)
);

A2O1A1Ixp33_ASAP7_75t_L g4873 ( 
.A1(n_4611),
.A2(n_65),
.B(n_62),
.C(n_64),
.Y(n_4873)
);

AND2x2_ASAP7_75t_L g4874 ( 
.A(n_4567),
.B(n_64),
.Y(n_4874)
);

OAI22xp5_ASAP7_75t_L g4875 ( 
.A1(n_4564),
.A2(n_2276),
.B1(n_2289),
.B2(n_2253),
.Y(n_4875)
);

OAI22x1_ASAP7_75t_L g4876 ( 
.A1(n_4556),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_L g4877 ( 
.A(n_4441),
.B(n_70),
.Y(n_4877)
);

AOI22xp5_ASAP7_75t_L g4878 ( 
.A1(n_4532),
.A2(n_2289),
.B1(n_2292),
.B2(n_2276),
.Y(n_4878)
);

O2A1O1Ixp33_ASAP7_75t_SL g4879 ( 
.A1(n_4582),
.A2(n_87),
.B(n_97),
.C(n_72),
.Y(n_4879)
);

OAI22x1_ASAP7_75t_L g4880 ( 
.A1(n_4556),
.A2(n_77),
.B1(n_73),
.B2(n_75),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4446),
.Y(n_4881)
);

AND2x4_ASAP7_75t_L g4882 ( 
.A(n_4568),
.B(n_648),
.Y(n_4882)
);

AOI21xp5_ASAP7_75t_L g4883 ( 
.A1(n_4448),
.A2(n_2292),
.B(n_2289),
.Y(n_4883)
);

CKINVDCx11_ASAP7_75t_R g4884 ( 
.A(n_4539),
.Y(n_4884)
);

AOI22xp33_ASAP7_75t_L g4885 ( 
.A1(n_4452),
.A2(n_4464),
.B1(n_4564),
.B2(n_4588),
.Y(n_4885)
);

INVx2_ASAP7_75t_L g4886 ( 
.A(n_4552),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4561),
.B(n_73),
.Y(n_4887)
);

INVx3_ASAP7_75t_L g4888 ( 
.A(n_4547),
.Y(n_4888)
);

NOR4xp25_ASAP7_75t_L g4889 ( 
.A(n_4584),
.B(n_79),
.C(n_75),
.D(n_78),
.Y(n_4889)
);

BUFx8_ASAP7_75t_L g4890 ( 
.A(n_4547),
.Y(n_4890)
);

NOR2xp33_ASAP7_75t_L g4891 ( 
.A(n_4570),
.B(n_80),
.Y(n_4891)
);

AOI21xp5_ASAP7_75t_L g4892 ( 
.A1(n_4458),
.A2(n_2299),
.B(n_2292),
.Y(n_4892)
);

A2O1A1Ixp33_ASAP7_75t_L g4893 ( 
.A1(n_4585),
.A2(n_88),
.B(n_80),
.C(n_83),
.Y(n_4893)
);

AO31x2_ASAP7_75t_L g4894 ( 
.A1(n_4462),
.A2(n_93),
.A3(n_89),
.B(n_92),
.Y(n_4894)
);

O2A1O1Ixp33_ASAP7_75t_SL g4895 ( 
.A1(n_4462),
.A2(n_101),
.B(n_109),
.C(n_89),
.Y(n_4895)
);

AOI21xp5_ASAP7_75t_L g4896 ( 
.A1(n_4462),
.A2(n_2299),
.B(n_2292),
.Y(n_4896)
);

AO32x2_ASAP7_75t_L g4897 ( 
.A1(n_4474),
.A2(n_95),
.A3(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_4897)
);

AOI21xp5_ASAP7_75t_L g4898 ( 
.A1(n_4474),
.A2(n_2307),
.B(n_2299),
.Y(n_4898)
);

NOR2xp33_ASAP7_75t_SL g4899 ( 
.A(n_4474),
.B(n_2299),
.Y(n_4899)
);

NOR2xp33_ASAP7_75t_L g4900 ( 
.A(n_4484),
.B(n_94),
.Y(n_4900)
);

AOI21xp5_ASAP7_75t_L g4901 ( 
.A1(n_4484),
.A2(n_2309),
.B(n_2307),
.Y(n_4901)
);

OAI21x1_ASAP7_75t_L g4902 ( 
.A1(n_4484),
.A2(n_652),
.B(n_649),
.Y(n_4902)
);

INVx2_ASAP7_75t_L g4903 ( 
.A(n_4743),
.Y(n_4903)
);

OAI21x1_ASAP7_75t_L g4904 ( 
.A1(n_4661),
.A2(n_4508),
.B(n_4501),
.Y(n_4904)
);

INVx2_ASAP7_75t_L g4905 ( 
.A(n_4763),
.Y(n_4905)
);

OAI22xp5_ASAP7_75t_L g4906 ( 
.A1(n_4698),
.A2(n_4508),
.B1(n_4540),
.B2(n_4501),
.Y(n_4906)
);

OR2x2_ASAP7_75t_L g4907 ( 
.A(n_4814),
.B(n_4501),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4785),
.B(n_4508),
.Y(n_4908)
);

AOI22xp33_ASAP7_75t_L g4909 ( 
.A1(n_4683),
.A2(n_4554),
.B1(n_4579),
.B2(n_4540),
.Y(n_4909)
);

INVx2_ASAP7_75t_L g4910 ( 
.A(n_4667),
.Y(n_4910)
);

AOI22xp33_ASAP7_75t_SL g4911 ( 
.A1(n_4683),
.A2(n_4728),
.B1(n_4863),
.B2(n_4692),
.Y(n_4911)
);

BUFx3_ASAP7_75t_L g4912 ( 
.A(n_4662),
.Y(n_4912)
);

CKINVDCx20_ASAP7_75t_R g4913 ( 
.A(n_4663),
.Y(n_4913)
);

INVx2_ASAP7_75t_L g4914 ( 
.A(n_4690),
.Y(n_4914)
);

NOR2x1_ASAP7_75t_SL g4915 ( 
.A(n_4642),
.B(n_4540),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4717),
.B(n_4554),
.Y(n_4916)
);

INVx1_ASAP7_75t_L g4917 ( 
.A(n_4700),
.Y(n_4917)
);

AND2x2_ASAP7_75t_L g4918 ( 
.A(n_4757),
.B(n_4554),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_4779),
.B(n_4579),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4713),
.Y(n_4920)
);

INVx6_ASAP7_75t_L g4921 ( 
.A(n_4796),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4719),
.Y(n_4922)
);

OAI22xp5_ASAP7_75t_L g4923 ( 
.A1(n_4850),
.A2(n_4592),
.B1(n_4593),
.B2(n_4579),
.Y(n_4923)
);

AOI22xp33_ASAP7_75t_L g4924 ( 
.A1(n_4843),
.A2(n_4593),
.B1(n_4592),
.B2(n_2309),
.Y(n_4924)
);

AOI221xp5_ASAP7_75t_L g4925 ( 
.A1(n_4737),
.A2(n_4889),
.B1(n_4816),
.B2(n_4821),
.C(n_4848),
.Y(n_4925)
);

BUFx3_ASAP7_75t_L g4926 ( 
.A(n_4680),
.Y(n_4926)
);

INVx2_ASAP7_75t_L g4927 ( 
.A(n_4722),
.Y(n_4927)
);

INVx2_ASAP7_75t_L g4928 ( 
.A(n_4727),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4734),
.Y(n_4929)
);

CKINVDCx11_ASAP7_75t_R g4930 ( 
.A(n_4707),
.Y(n_4930)
);

BUFx2_ASAP7_75t_L g4931 ( 
.A(n_4657),
.Y(n_4931)
);

OAI22xp5_ASAP7_75t_L g4932 ( 
.A1(n_4701),
.A2(n_4593),
.B1(n_4592),
.B2(n_99),
.Y(n_4932)
);

OAI22xp5_ASAP7_75t_L g4933 ( 
.A1(n_4764),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_4933)
);

AOI22xp5_ASAP7_75t_L g4934 ( 
.A1(n_4716),
.A2(n_2309),
.B1(n_2369),
.B2(n_2307),
.Y(n_4934)
);

INVx4_ASAP7_75t_L g4935 ( 
.A(n_4652),
.Y(n_4935)
);

OR2x2_ASAP7_75t_L g4936 ( 
.A(n_4646),
.B(n_100),
.Y(n_4936)
);

INVx2_ASAP7_75t_SL g4937 ( 
.A(n_4720),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4738),
.Y(n_4938)
);

CKINVDCx5p33_ASAP7_75t_R g4939 ( 
.A(n_4666),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_4673),
.B(n_101),
.Y(n_4940)
);

OAI22xp5_ASAP7_75t_L g4941 ( 
.A1(n_4873),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_4748),
.Y(n_4942)
);

AND2x4_ASAP7_75t_L g4943 ( 
.A(n_4791),
.B(n_102),
.Y(n_4943)
);

OR2x2_ASAP7_75t_L g4944 ( 
.A(n_4656),
.B(n_4733),
.Y(n_4944)
);

AOI22xp33_ASAP7_75t_L g4945 ( 
.A1(n_4840),
.A2(n_2309),
.B1(n_2369),
.B2(n_2307),
.Y(n_4945)
);

AOI222xp33_ASAP7_75t_L g4946 ( 
.A1(n_4674),
.A2(n_107),
.B1(n_109),
.B2(n_105),
.C1(n_106),
.C2(n_108),
.Y(n_4946)
);

INVx3_ASAP7_75t_L g4947 ( 
.A(n_4652),
.Y(n_4947)
);

AOI22xp33_ASAP7_75t_L g4948 ( 
.A1(n_4746),
.A2(n_4813),
.B1(n_4644),
.B2(n_4725),
.Y(n_4948)
);

INVx11_ASAP7_75t_L g4949 ( 
.A(n_4890),
.Y(n_4949)
);

AND2x2_ASAP7_75t_L g4950 ( 
.A(n_4829),
.B(n_106),
.Y(n_4950)
);

BUFx2_ASAP7_75t_L g4951 ( 
.A(n_4778),
.Y(n_4951)
);

OAI22xp5_ASAP7_75t_L g4952 ( 
.A1(n_4893),
.A2(n_114),
.B1(n_110),
.B2(n_112),
.Y(n_4952)
);

NOR2xp67_ASAP7_75t_L g4953 ( 
.A(n_4783),
.B(n_112),
.Y(n_4953)
);

AOI21xp5_ASAP7_75t_L g4954 ( 
.A1(n_4643),
.A2(n_2385),
.B(n_2369),
.Y(n_4954)
);

INVx8_ASAP7_75t_L g4955 ( 
.A(n_4739),
.Y(n_4955)
);

AOI22xp33_ASAP7_75t_L g4956 ( 
.A1(n_4679),
.A2(n_2385),
.B1(n_2395),
.B2(n_2369),
.Y(n_4956)
);

OAI22xp33_ASAP7_75t_SL g4957 ( 
.A1(n_4825),
.A2(n_118),
.B1(n_114),
.B2(n_117),
.Y(n_4957)
);

INVx1_ASAP7_75t_SL g4958 ( 
.A(n_4678),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4828),
.B(n_4641),
.Y(n_4959)
);

A2O1A1Ixp33_ASAP7_75t_L g4960 ( 
.A1(n_4639),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4672),
.B(n_119),
.Y(n_4961)
);

AND2x2_ASAP7_75t_L g4962 ( 
.A(n_4854),
.B(n_121),
.Y(n_4962)
);

AOI222xp33_ASAP7_75t_L g4963 ( 
.A1(n_4695),
.A2(n_125),
.B1(n_127),
.B2(n_121),
.C1(n_124),
.C2(n_126),
.Y(n_4963)
);

OAI22xp5_ASAP7_75t_L g4964 ( 
.A1(n_4820),
.A2(n_4846),
.B1(n_4808),
.B2(n_4885),
.Y(n_4964)
);

AOI21xp33_ASAP7_75t_L g4965 ( 
.A1(n_4735),
.A2(n_124),
.B(n_127),
.Y(n_4965)
);

INVx2_ASAP7_75t_L g4966 ( 
.A(n_4755),
.Y(n_4966)
);

NAND2x1_ASAP7_75t_L g4967 ( 
.A(n_4792),
.B(n_2442),
.Y(n_4967)
);

A2O1A1Ixp33_ASAP7_75t_L g4968 ( 
.A1(n_4806),
.A2(n_4685),
.B(n_4697),
.C(n_4671),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4759),
.Y(n_4969)
);

BUFx2_ASAP7_75t_L g4970 ( 
.A(n_4784),
.Y(n_4970)
);

AOI22xp33_ASAP7_75t_L g4971 ( 
.A1(n_4876),
.A2(n_2395),
.B1(n_2398),
.B2(n_2385),
.Y(n_4971)
);

BUFx10_ASAP7_75t_L g4972 ( 
.A(n_4658),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4773),
.Y(n_4973)
);

HB1xp67_ASAP7_75t_L g4974 ( 
.A(n_4795),
.Y(n_4974)
);

OR2x6_ASAP7_75t_L g4975 ( 
.A(n_4860),
.B(n_2385),
.Y(n_4975)
);

BUFx6f_ASAP7_75t_L g4976 ( 
.A(n_4884),
.Y(n_4976)
);

AOI22xp33_ASAP7_75t_SL g4977 ( 
.A1(n_4704),
.A2(n_133),
.B1(n_128),
.B2(n_132),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4774),
.Y(n_4978)
);

A2O1A1Ixp33_ASAP7_75t_L g4979 ( 
.A1(n_4653),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_4979)
);

NOR2xp67_ASAP7_75t_L g4980 ( 
.A(n_4652),
.B(n_4694),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4804),
.Y(n_4981)
);

AOI221xp5_ASAP7_75t_L g4982 ( 
.A1(n_4880),
.A2(n_137),
.B1(n_135),
.B2(n_136),
.C(n_138),
.Y(n_4982)
);

INVx2_ASAP7_75t_L g4983 ( 
.A(n_4809),
.Y(n_4983)
);

AOI22xp33_ASAP7_75t_L g4984 ( 
.A1(n_4771),
.A2(n_2398),
.B1(n_2412),
.B2(n_2395),
.Y(n_4984)
);

AO21x1_ASAP7_75t_L g4985 ( 
.A1(n_4897),
.A2(n_135),
.B(n_136),
.Y(n_4985)
);

OAI22xp5_ASAP7_75t_L g4986 ( 
.A1(n_4856),
.A2(n_141),
.B1(n_137),
.B2(n_139),
.Y(n_4986)
);

CKINVDCx5p33_ASAP7_75t_R g4987 ( 
.A(n_4705),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4818),
.Y(n_4988)
);

AOI22xp33_ASAP7_75t_L g4989 ( 
.A1(n_4862),
.A2(n_2398),
.B1(n_2412),
.B2(n_2395),
.Y(n_4989)
);

INVx4_ASAP7_75t_L g4990 ( 
.A(n_4694),
.Y(n_4990)
);

CKINVDCx5p33_ASAP7_75t_R g4991 ( 
.A(n_4794),
.Y(n_4991)
);

AOI22xp33_ASAP7_75t_L g4992 ( 
.A1(n_4758),
.A2(n_2412),
.B1(n_2417),
.B2(n_2398),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4881),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4787),
.Y(n_4994)
);

OAI22xp33_ASAP7_75t_L g4995 ( 
.A1(n_4815),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4827),
.Y(n_4996)
);

INVx2_ASAP7_75t_L g4997 ( 
.A(n_4852),
.Y(n_4997)
);

O2A1O1Ixp33_ASAP7_75t_L g4998 ( 
.A1(n_4687),
.A2(n_146),
.B(n_142),
.C(n_145),
.Y(n_4998)
);

INVxp67_ASAP7_75t_L g4999 ( 
.A(n_4647),
.Y(n_4999)
);

INVx2_ASAP7_75t_L g5000 ( 
.A(n_4855),
.Y(n_5000)
);

O2A1O1Ixp33_ASAP7_75t_L g5001 ( 
.A1(n_4761),
.A2(n_149),
.B(n_145),
.C(n_148),
.Y(n_5001)
);

AOI22xp5_ASAP7_75t_L g5002 ( 
.A1(n_4706),
.A2(n_2442),
.B1(n_2417),
.B2(n_2424),
.Y(n_5002)
);

INVx2_ASAP7_75t_SL g5003 ( 
.A(n_4793),
.Y(n_5003)
);

O2A1O1Ixp5_ASAP7_75t_L g5004 ( 
.A1(n_4710),
.A2(n_4768),
.B(n_4640),
.C(n_4900),
.Y(n_5004)
);

INVx2_ASAP7_75t_L g5005 ( 
.A(n_4870),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4824),
.Y(n_5006)
);

OAI22xp33_ASAP7_75t_L g5007 ( 
.A1(n_4833),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_5007)
);

OAI22xp5_ASAP7_75t_L g5008 ( 
.A1(n_4682),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_5008)
);

INVx8_ASAP7_75t_L g5009 ( 
.A(n_4786),
.Y(n_5009)
);

AOI221xp5_ASAP7_75t_L g5010 ( 
.A1(n_4677),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.C(n_158),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4824),
.Y(n_5011)
);

OAI22xp5_ASAP7_75t_L g5012 ( 
.A1(n_4754),
.A2(n_159),
.B1(n_155),
.B2(n_156),
.Y(n_5012)
);

AOI22xp5_ASAP7_75t_L g5013 ( 
.A1(n_4740),
.A2(n_2442),
.B1(n_2417),
.B2(n_2424),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4675),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_4703),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4837),
.Y(n_5016)
);

A2O1A1Ixp33_ASAP7_75t_L g5017 ( 
.A1(n_4742),
.A2(n_168),
.B(n_162),
.C(n_164),
.Y(n_5017)
);

INVx2_ASAP7_75t_L g5018 ( 
.A(n_4886),
.Y(n_5018)
);

INVx1_ASAP7_75t_SL g5019 ( 
.A(n_4867),
.Y(n_5019)
);

NAND2x1p5_ASAP7_75t_L g5020 ( 
.A(n_4694),
.B(n_2412),
.Y(n_5020)
);

OAI21xp5_ASAP7_75t_L g5021 ( 
.A1(n_4776),
.A2(n_162),
.B(n_168),
.Y(n_5021)
);

AOI22xp33_ASAP7_75t_SL g5022 ( 
.A1(n_4819),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_5022)
);

OAI211xp5_ASAP7_75t_L g5023 ( 
.A1(n_4872),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_4897),
.Y(n_5024)
);

INVx4_ASAP7_75t_L g5025 ( 
.A(n_4715),
.Y(n_5025)
);

OR2x2_ASAP7_75t_L g5026 ( 
.A(n_4831),
.B(n_172),
.Y(n_5026)
);

BUFx3_ASAP7_75t_L g5027 ( 
.A(n_4645),
.Y(n_5027)
);

OAI22xp5_ASAP7_75t_L g5028 ( 
.A1(n_4718),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_5028)
);

NAND2xp5_ASAP7_75t_L g5029 ( 
.A(n_4857),
.B(n_4686),
.Y(n_5029)
);

NAND2x1p5_ASAP7_75t_L g5030 ( 
.A(n_4711),
.B(n_2417),
.Y(n_5030)
);

BUFx2_ASAP7_75t_L g5031 ( 
.A(n_4669),
.Y(n_5031)
);

OAI222xp33_ASAP7_75t_L g5032 ( 
.A1(n_4801),
.A2(n_178),
.B1(n_180),
.B2(n_174),
.C1(n_175),
.C2(n_179),
.Y(n_5032)
);

AND2x4_ASAP7_75t_L g5033 ( 
.A(n_4851),
.B(n_178),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_L g5034 ( 
.A(n_4765),
.B(n_181),
.Y(n_5034)
);

INVx2_ASAP7_75t_L g5035 ( 
.A(n_4853),
.Y(n_5035)
);

AOI22xp33_ASAP7_75t_L g5036 ( 
.A1(n_4859),
.A2(n_2427),
.B1(n_2442),
.B2(n_2424),
.Y(n_5036)
);

INVx2_ASAP7_75t_L g5037 ( 
.A(n_4762),
.Y(n_5037)
);

BUFx6f_ASAP7_75t_L g5038 ( 
.A(n_4745),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_SL g5039 ( 
.A(n_4756),
.B(n_2424),
.Y(n_5039)
);

CKINVDCx20_ASAP7_75t_R g5040 ( 
.A(n_4709),
.Y(n_5040)
);

AOI22xp33_ASAP7_75t_L g5041 ( 
.A1(n_4760),
.A2(n_2427),
.B1(n_186),
.B2(n_184),
.Y(n_5041)
);

AOI22xp5_ASAP7_75t_L g5042 ( 
.A1(n_4648),
.A2(n_2427),
.B1(n_188),
.B2(n_185),
.Y(n_5042)
);

AND2x2_ASAP7_75t_L g5043 ( 
.A(n_4751),
.B(n_185),
.Y(n_5043)
);

OR2x6_ASAP7_75t_L g5044 ( 
.A(n_4834),
.B(n_2427),
.Y(n_5044)
);

HB1xp67_ASAP7_75t_L g5045 ( 
.A(n_4770),
.Y(n_5045)
);

BUFx2_ASAP7_75t_L g5046 ( 
.A(n_4780),
.Y(n_5046)
);

OAI221xp5_ASAP7_75t_L g5047 ( 
.A1(n_4721),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_5047)
);

NAND2xp5_ASAP7_75t_L g5048 ( 
.A(n_4752),
.B(n_187),
.Y(n_5048)
);

AOI221xp5_ASAP7_75t_L g5049 ( 
.A1(n_4769),
.A2(n_4861),
.B1(n_4830),
.B2(n_4879),
.C(n_4660),
.Y(n_5049)
);

NAND3xp33_ASAP7_75t_L g5050 ( 
.A(n_4777),
.B(n_192),
.C(n_193),
.Y(n_5050)
);

OAI22xp5_ASAP7_75t_L g5051 ( 
.A1(n_4665),
.A2(n_4845),
.B1(n_4651),
.B2(n_4731),
.Y(n_5051)
);

CKINVDCx5p33_ASAP7_75t_R g5052 ( 
.A(n_4842),
.Y(n_5052)
);

OAI22xp5_ASAP7_75t_L g5053 ( 
.A1(n_4696),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_5053)
);

INVx3_ASAP7_75t_L g5054 ( 
.A(n_4723),
.Y(n_5054)
);

NOR2xp33_ASAP7_75t_L g5055 ( 
.A(n_4681),
.B(n_195),
.Y(n_5055)
);

AOI22xp33_ASAP7_75t_L g5056 ( 
.A1(n_4684),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_5056)
);

OAI22xp5_ASAP7_75t_L g5057 ( 
.A1(n_4691),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_5057)
);

AND2x2_ASAP7_75t_L g5058 ( 
.A(n_4826),
.B(n_199),
.Y(n_5058)
);

AOI22xp33_ASAP7_75t_L g5059 ( 
.A1(n_4891),
.A2(n_205),
.B1(n_201),
.B2(n_203),
.Y(n_5059)
);

AOI22xp33_ASAP7_75t_L g5060 ( 
.A1(n_4767),
.A2(n_207),
.B1(n_203),
.B2(n_206),
.Y(n_5060)
);

AOI221x1_ASAP7_75t_SL g5061 ( 
.A1(n_4736),
.A2(n_209),
.B1(n_206),
.B2(n_208),
.C(n_210),
.Y(n_5061)
);

INVx1_ASAP7_75t_SL g5062 ( 
.A(n_4812),
.Y(n_5062)
);

O2A1O1Ixp33_ASAP7_75t_L g5063 ( 
.A1(n_4895),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_5063)
);

CKINVDCx5p33_ASAP7_75t_R g5064 ( 
.A(n_4844),
.Y(n_5064)
);

AOI22xp33_ASAP7_75t_L g5065 ( 
.A1(n_4693),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_5065)
);

OAI211xp5_ASAP7_75t_SL g5066 ( 
.A1(n_4772),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_5066)
);

OAI21x1_ASAP7_75t_L g5067 ( 
.A1(n_4650),
.A2(n_659),
.B(n_653),
.Y(n_5067)
);

AOI22xp33_ASAP7_75t_SL g5068 ( 
.A1(n_4811),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_5068)
);

AOI22xp5_ASAP7_75t_L g5069 ( 
.A1(n_4668),
.A2(n_220),
.B1(n_217),
.B2(n_218),
.Y(n_5069)
);

INVx2_ASAP7_75t_L g5070 ( 
.A(n_4762),
.Y(n_5070)
);

AOI22xp33_ASAP7_75t_SL g5071 ( 
.A1(n_4838),
.A2(n_223),
.B1(n_220),
.B2(n_222),
.Y(n_5071)
);

INVx3_ASAP7_75t_L g5072 ( 
.A(n_4800),
.Y(n_5072)
);

AO21x2_ASAP7_75t_L g5073 ( 
.A1(n_4712),
.A2(n_222),
.B(n_223),
.Y(n_5073)
);

INVx2_ASAP7_75t_L g5074 ( 
.A(n_4894),
.Y(n_5074)
);

INVx3_ASAP7_75t_L g5075 ( 
.A(n_4871),
.Y(n_5075)
);

AOI22xp33_ASAP7_75t_L g5076 ( 
.A1(n_4744),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_5076)
);

INVx2_ASAP7_75t_L g5077 ( 
.A(n_4894),
.Y(n_5077)
);

BUFx12f_ASAP7_75t_L g5078 ( 
.A(n_4882),
.Y(n_5078)
);

HB1xp67_ASAP7_75t_L g5079 ( 
.A(n_4770),
.Y(n_5079)
);

OAI22xp5_ASAP7_75t_L g5080 ( 
.A1(n_4834),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_5080)
);

AND2x4_ASAP7_75t_L g5081 ( 
.A(n_4888),
.B(n_228),
.Y(n_5081)
);

AOI22xp33_ASAP7_75t_L g5082 ( 
.A1(n_4817),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_5082)
);

INVx1_ASAP7_75t_L g5083 ( 
.A(n_4897),
.Y(n_5083)
);

OAI22xp5_ASAP7_75t_L g5084 ( 
.A1(n_4847),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_4788),
.Y(n_5085)
);

AOI22xp33_ASAP7_75t_L g5086 ( 
.A1(n_4789),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4788),
.Y(n_5087)
);

AND2x2_ASAP7_75t_L g5088 ( 
.A(n_4874),
.B(n_232),
.Y(n_5088)
);

NAND2x1_ASAP7_75t_L g5089 ( 
.A(n_4724),
.B(n_233),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4868),
.Y(n_5090)
);

OAI22xp5_ASAP7_75t_L g5091 ( 
.A1(n_4878),
.A2(n_4869),
.B1(n_4835),
.B2(n_4803),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4877),
.Y(n_5092)
);

INVxp67_ASAP7_75t_L g5093 ( 
.A(n_4887),
.Y(n_5093)
);

AOI22xp33_ASAP7_75t_L g5094 ( 
.A1(n_4797),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_L g5095 ( 
.A(n_4822),
.B(n_235),
.Y(n_5095)
);

AND2x4_ASAP7_75t_L g5096 ( 
.A(n_4766),
.B(n_236),
.Y(n_5096)
);

AOI22xp33_ASAP7_75t_L g5097 ( 
.A1(n_4839),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_5097)
);

BUFx6f_ASAP7_75t_L g5098 ( 
.A(n_4664),
.Y(n_5098)
);

AND2x2_ASAP7_75t_L g5099 ( 
.A(n_4688),
.B(n_240),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4849),
.Y(n_5100)
);

NAND2xp5_ASAP7_75t_L g5101 ( 
.A(n_4670),
.B(n_241),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_4849),
.Y(n_5102)
);

BUFx12f_ASAP7_75t_L g5103 ( 
.A(n_4899),
.Y(n_5103)
);

AOI21xp5_ASAP7_75t_L g5104 ( 
.A1(n_4649),
.A2(n_2037),
.B(n_1793),
.Y(n_5104)
);

NOR2xp33_ASAP7_75t_L g5105 ( 
.A(n_4999),
.B(n_4781),
.Y(n_5105)
);

INVx2_ASAP7_75t_L g5106 ( 
.A(n_4951),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_4917),
.Y(n_5107)
);

INVx2_ASAP7_75t_L g5108 ( 
.A(n_4981),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_4910),
.Y(n_5109)
);

CKINVDCx20_ASAP7_75t_R g5110 ( 
.A(n_4913),
.Y(n_5110)
);

INVx3_ASAP7_75t_L g5111 ( 
.A(n_4947),
.Y(n_5111)
);

INVx3_ASAP7_75t_L g5112 ( 
.A(n_4947),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4920),
.Y(n_5113)
);

OR2x2_ASAP7_75t_L g5114 ( 
.A(n_4944),
.B(n_4702),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4922),
.Y(n_5115)
);

INVx2_ASAP7_75t_L g5116 ( 
.A(n_4914),
.Y(n_5116)
);

OAI21x1_ASAP7_75t_L g5117 ( 
.A1(n_5037),
.A2(n_4708),
.B(n_4714),
.Y(n_5117)
);

INVx2_ASAP7_75t_L g5118 ( 
.A(n_4927),
.Y(n_5118)
);

INVx2_ASAP7_75t_L g5119 ( 
.A(n_4928),
.Y(n_5119)
);

HB1xp67_ASAP7_75t_L g5120 ( 
.A(n_4974),
.Y(n_5120)
);

INVx1_ASAP7_75t_L g5121 ( 
.A(n_4929),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4938),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_4969),
.Y(n_5123)
);

INVx1_ASAP7_75t_L g5124 ( 
.A(n_4973),
.Y(n_5124)
);

INVx2_ASAP7_75t_L g5125 ( 
.A(n_4942),
.Y(n_5125)
);

INVx1_ASAP7_75t_L g5126 ( 
.A(n_4978),
.Y(n_5126)
);

OAI22xp5_ASAP7_75t_L g5127 ( 
.A1(n_4911),
.A2(n_4858),
.B1(n_4849),
.B2(n_4736),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_4988),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_4988),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_4966),
.Y(n_5130)
);

INVx2_ASAP7_75t_L g5131 ( 
.A(n_4983),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_5102),
.B(n_4790),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_4993),
.Y(n_5133)
);

AOI21xp5_ASAP7_75t_L g5134 ( 
.A1(n_4954),
.A2(n_4753),
.B(n_4782),
.Y(n_5134)
);

OAI21xp5_ASAP7_75t_L g5135 ( 
.A1(n_4953),
.A2(n_4902),
.B(n_4832),
.Y(n_5135)
);

INVx2_ASAP7_75t_L g5136 ( 
.A(n_4903),
.Y(n_5136)
);

INVx3_ASAP7_75t_L g5137 ( 
.A(n_5025),
.Y(n_5137)
);

INVx2_ASAP7_75t_L g5138 ( 
.A(n_4905),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_4994),
.Y(n_5139)
);

INVx2_ASAP7_75t_L g5140 ( 
.A(n_4997),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_4996),
.Y(n_5141)
);

INVx2_ASAP7_75t_L g5142 ( 
.A(n_4931),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_5000),
.Y(n_5143)
);

INVx2_ASAP7_75t_L g5144 ( 
.A(n_4907),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_5005),
.Y(n_5145)
);

INVx3_ASAP7_75t_L g5146 ( 
.A(n_5025),
.Y(n_5146)
);

INVx1_ASAP7_75t_L g5147 ( 
.A(n_5014),
.Y(n_5147)
);

INVx4_ASAP7_75t_L g5148 ( 
.A(n_4976),
.Y(n_5148)
);

BUFx6f_ASAP7_75t_L g5149 ( 
.A(n_4976),
.Y(n_5149)
);

BUFx6f_ASAP7_75t_L g5150 ( 
.A(n_4976),
.Y(n_5150)
);

INVx3_ASAP7_75t_L g5151 ( 
.A(n_5072),
.Y(n_5151)
);

INVx1_ASAP7_75t_L g5152 ( 
.A(n_5015),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_5006),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5011),
.Y(n_5154)
);

INVx3_ASAP7_75t_L g5155 ( 
.A(n_5072),
.Y(n_5155)
);

AND2x4_ASAP7_75t_L g5156 ( 
.A(n_4970),
.B(n_4836),
.Y(n_5156)
);

INVx1_ASAP7_75t_L g5157 ( 
.A(n_4959),
.Y(n_5157)
);

AND2x2_ASAP7_75t_L g5158 ( 
.A(n_4916),
.B(n_4732),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_5018),
.Y(n_5159)
);

NOR2xp33_ASAP7_75t_L g5160 ( 
.A(n_5090),
.B(n_4823),
.Y(n_5160)
);

INVx2_ASAP7_75t_L g5161 ( 
.A(n_5035),
.Y(n_5161)
);

INVx2_ASAP7_75t_L g5162 ( 
.A(n_5031),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_5085),
.Y(n_5163)
);

INVx2_ASAP7_75t_L g5164 ( 
.A(n_4918),
.Y(n_5164)
);

INVx1_ASAP7_75t_SL g5165 ( 
.A(n_4958),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_L g5166 ( 
.A(n_5102),
.B(n_4741),
.Y(n_5166)
);

AND2x2_ASAP7_75t_L g5167 ( 
.A(n_5046),
.B(n_4732),
.Y(n_5167)
);

NAND2xp5_ASAP7_75t_L g5168 ( 
.A(n_5024),
.B(n_5083),
.Y(n_5168)
);

INVx2_ASAP7_75t_SL g5169 ( 
.A(n_5038),
.Y(n_5169)
);

OR2x2_ASAP7_75t_L g5170 ( 
.A(n_4908),
.B(n_4702),
.Y(n_5170)
);

INVx4_ASAP7_75t_SL g5171 ( 
.A(n_4921),
.Y(n_5171)
);

OAI21x1_ASAP7_75t_L g5172 ( 
.A1(n_5070),
.A2(n_4807),
.B(n_4841),
.Y(n_5172)
);

INVx2_ASAP7_75t_L g5173 ( 
.A(n_5074),
.Y(n_5173)
);

INVxp67_ASAP7_75t_L g5174 ( 
.A(n_5045),
.Y(n_5174)
);

INVx2_ASAP7_75t_L g5175 ( 
.A(n_5077),
.Y(n_5175)
);

AND2x2_ASAP7_75t_L g5176 ( 
.A(n_5093),
.B(n_4732),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_4919),
.Y(n_5177)
);

INVx3_ASAP7_75t_L g5178 ( 
.A(n_4935),
.Y(n_5178)
);

BUFx2_ASAP7_75t_L g5179 ( 
.A(n_5075),
.Y(n_5179)
);

INVx2_ASAP7_75t_L g5180 ( 
.A(n_5016),
.Y(n_5180)
);

NOR2x1_ASAP7_75t_L g5181 ( 
.A(n_4980),
.B(n_4805),
.Y(n_5181)
);

INVx2_ASAP7_75t_L g5182 ( 
.A(n_4915),
.Y(n_5182)
);

BUFx2_ASAP7_75t_L g5183 ( 
.A(n_5075),
.Y(n_5183)
);

INVx2_ASAP7_75t_L g5184 ( 
.A(n_4915),
.Y(n_5184)
);

AND2x2_ASAP7_75t_L g5185 ( 
.A(n_5019),
.B(n_4654),
.Y(n_5185)
);

INVx3_ASAP7_75t_L g5186 ( 
.A(n_4935),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_5087),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_5092),
.Y(n_5188)
);

OAI21x1_ASAP7_75t_L g5189 ( 
.A1(n_4967),
.A2(n_4810),
.B(n_4749),
.Y(n_5189)
);

BUFx2_ASAP7_75t_L g5190 ( 
.A(n_5054),
.Y(n_5190)
);

INVx2_ASAP7_75t_L g5191 ( 
.A(n_4904),
.Y(n_5191)
);

INVx2_ASAP7_75t_L g5192 ( 
.A(n_4926),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_5079),
.Y(n_5193)
);

INVx4_ASAP7_75t_L g5194 ( 
.A(n_4949),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_L g5195 ( 
.A(n_5100),
.B(n_4654),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_4936),
.Y(n_5196)
);

OR2x6_ASAP7_75t_L g5197 ( 
.A(n_4975),
.B(n_4883),
.Y(n_5197)
);

INVx2_ASAP7_75t_L g5198 ( 
.A(n_5062),
.Y(n_5198)
);

INVx2_ASAP7_75t_L g5199 ( 
.A(n_5003),
.Y(n_5199)
);

INVx3_ASAP7_75t_L g5200 ( 
.A(n_4990),
.Y(n_5200)
);

INVx2_ASAP7_75t_SL g5201 ( 
.A(n_5038),
.Y(n_5201)
);

AO21x2_ASAP7_75t_L g5202 ( 
.A1(n_4985),
.A2(n_4659),
.B(n_4726),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_4961),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_4940),
.Y(n_5204)
);

INVx2_ASAP7_75t_L g5205 ( 
.A(n_5096),
.Y(n_5205)
);

BUFx6f_ASAP7_75t_L g5206 ( 
.A(n_5038),
.Y(n_5206)
);

INVxp33_ASAP7_75t_L g5207 ( 
.A(n_4930),
.Y(n_5207)
);

INVx3_ASAP7_75t_L g5208 ( 
.A(n_4990),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_4937),
.B(n_4750),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_4943),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_4943),
.Y(n_5211)
);

BUFx2_ASAP7_75t_L g5212 ( 
.A(n_5054),
.Y(n_5212)
);

OAI21x1_ASAP7_75t_L g5213 ( 
.A1(n_5004),
.A2(n_4699),
.B(n_4747),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_4950),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_4975),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_5096),
.Y(n_5216)
);

CKINVDCx11_ASAP7_75t_R g5217 ( 
.A(n_5040),
.Y(n_5217)
);

BUFx6f_ASAP7_75t_L g5218 ( 
.A(n_4921),
.Y(n_5218)
);

OAI21x1_ASAP7_75t_L g5219 ( 
.A1(n_5067),
.A2(n_4802),
.B(n_4676),
.Y(n_5219)
);

INVx2_ASAP7_75t_L g5220 ( 
.A(n_5027),
.Y(n_5220)
);

OAI21x1_ASAP7_75t_L g5221 ( 
.A1(n_5089),
.A2(n_4775),
.B(n_4798),
.Y(n_5221)
);

OR2x6_ASAP7_75t_L g5222 ( 
.A(n_4955),
.B(n_4865),
.Y(n_5222)
);

AND2x2_ASAP7_75t_L g5223 ( 
.A(n_4912),
.B(n_4750),
.Y(n_5223)
);

AND2x2_ASAP7_75t_L g5224 ( 
.A(n_4962),
.B(n_4655),
.Y(n_5224)
);

OA21x2_ASAP7_75t_L g5225 ( 
.A1(n_5095),
.A2(n_4729),
.B(n_4864),
.Y(n_5225)
);

INVx3_ASAP7_75t_L g5226 ( 
.A(n_5098),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_5029),
.B(n_4655),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5073),
.Y(n_5228)
);

OAI22xp5_ASAP7_75t_L g5229 ( 
.A1(n_4948),
.A2(n_4858),
.B1(n_4736),
.B2(n_4866),
.Y(n_5229)
);

BUFx2_ASAP7_75t_L g5230 ( 
.A(n_5064),
.Y(n_5230)
);

BUFx4f_ASAP7_75t_SL g5231 ( 
.A(n_5078),
.Y(n_5231)
);

HB1xp67_ASAP7_75t_L g5232 ( 
.A(n_5099),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5026),
.Y(n_5233)
);

OAI21x1_ASAP7_75t_L g5234 ( 
.A1(n_5104),
.A2(n_4799),
.B(n_4892),
.Y(n_5234)
);

BUFx3_ASAP7_75t_L g5235 ( 
.A(n_4955),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_5033),
.Y(n_5236)
);

BUFx2_ASAP7_75t_L g5237 ( 
.A(n_4987),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_5033),
.Y(n_5238)
);

BUFx2_ASAP7_75t_L g5239 ( 
.A(n_4939),
.Y(n_5239)
);

INVx2_ASAP7_75t_L g5240 ( 
.A(n_5081),
.Y(n_5240)
);

HB1xp67_ASAP7_75t_L g5241 ( 
.A(n_5081),
.Y(n_5241)
);

INVx3_ASAP7_75t_L g5242 ( 
.A(n_5098),
.Y(n_5242)
);

CKINVDCx20_ASAP7_75t_R g5243 ( 
.A(n_4991),
.Y(n_5243)
);

AND2x2_ASAP7_75t_L g5244 ( 
.A(n_4972),
.B(n_4689),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5048),
.Y(n_5245)
);

BUFx2_ASAP7_75t_SL g5246 ( 
.A(n_4972),
.Y(n_5246)
);

CKINVDCx9p33_ASAP7_75t_R g5247 ( 
.A(n_5101),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5034),
.Y(n_5248)
);

CKINVDCx16_ASAP7_75t_R g5249 ( 
.A(n_5043),
.Y(n_5249)
);

OAI21x1_ASAP7_75t_L g5250 ( 
.A1(n_5039),
.A2(n_4898),
.B(n_4896),
.Y(n_5250)
);

OA21x2_ASAP7_75t_L g5251 ( 
.A1(n_4965),
.A2(n_4901),
.B(n_4875),
.Y(n_5251)
);

OA21x2_ASAP7_75t_L g5252 ( 
.A1(n_4925),
.A2(n_4730),
.B(n_4689),
.Y(n_5252)
);

INVx1_ASAP7_75t_L g5253 ( 
.A(n_5098),
.Y(n_5253)
);

BUFx2_ASAP7_75t_SL g5254 ( 
.A(n_5088),
.Y(n_5254)
);

INVx2_ASAP7_75t_L g5255 ( 
.A(n_5044),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_5061),
.B(n_4730),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5044),
.Y(n_5257)
);

OAI21x1_ASAP7_75t_L g5258 ( 
.A1(n_5020),
.A2(n_243),
.B(n_244),
.Y(n_5258)
);

INVx3_ASAP7_75t_L g5259 ( 
.A(n_5009),
.Y(n_5259)
);

AND2x4_ASAP7_75t_L g5260 ( 
.A(n_4909),
.B(n_243),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_L g5261 ( 
.A(n_5055),
.B(n_244),
.Y(n_5261)
);

OAI22xp5_ASAP7_75t_L g5262 ( 
.A1(n_5127),
.A2(n_4964),
.B1(n_4960),
.B2(n_5049),
.Y(n_5262)
);

AOI22xp5_ASAP7_75t_L g5263 ( 
.A1(n_5127),
.A2(n_5229),
.B1(n_4963),
.B2(n_5105),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5163),
.Y(n_5264)
);

BUFx2_ASAP7_75t_L g5265 ( 
.A(n_5190),
.Y(n_5265)
);

AOI22xp5_ASAP7_75t_L g5266 ( 
.A1(n_5229),
.A2(n_4941),
.B1(n_4952),
.B2(n_4946),
.Y(n_5266)
);

AOI21xp5_ASAP7_75t_L g5267 ( 
.A1(n_5135),
.A2(n_5021),
.B(n_5001),
.Y(n_5267)
);

AOI22xp33_ASAP7_75t_L g5268 ( 
.A1(n_5232),
.A2(n_5050),
.B1(n_5066),
.B2(n_5047),
.Y(n_5268)
);

AOI22xp33_ASAP7_75t_L g5269 ( 
.A1(n_5232),
.A2(n_4933),
.B1(n_5051),
.B2(n_4982),
.Y(n_5269)
);

OR2x2_ASAP7_75t_L g5270 ( 
.A(n_5166),
.B(n_5058),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_L g5271 ( 
.A(n_5157),
.B(n_4957),
.Y(n_5271)
);

AOI22xp33_ASAP7_75t_SL g5272 ( 
.A1(n_5246),
.A2(n_5023),
.B1(n_4986),
.B2(n_5012),
.Y(n_5272)
);

NOR2x1_ASAP7_75t_L g5273 ( 
.A(n_5235),
.B(n_5063),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_5187),
.Y(n_5274)
);

AOI222xp33_ASAP7_75t_L g5275 ( 
.A1(n_5261),
.A2(n_5010),
.B1(n_5053),
.B2(n_5076),
.C1(n_5065),
.C2(n_5028),
.Y(n_5275)
);

AOI22xp33_ASAP7_75t_L g5276 ( 
.A1(n_5228),
.A2(n_5233),
.B1(n_5248),
.B2(n_5245),
.Y(n_5276)
);

AOI22xp33_ASAP7_75t_L g5277 ( 
.A1(n_5205),
.A2(n_5022),
.B1(n_5068),
.B2(n_5008),
.Y(n_5277)
);

INVx5_ASAP7_75t_SL g5278 ( 
.A(n_5149),
.Y(n_5278)
);

CKINVDCx5p33_ASAP7_75t_R g5279 ( 
.A(n_5217),
.Y(n_5279)
);

OAI221xp5_ASAP7_75t_L g5280 ( 
.A1(n_5261),
.A2(n_5059),
.B1(n_5069),
.B2(n_4968),
.C(n_4979),
.Y(n_5280)
);

AOI22xp33_ASAP7_75t_L g5281 ( 
.A1(n_5205),
.A2(n_5041),
.B1(n_4932),
.B2(n_5056),
.Y(n_5281)
);

BUFx6f_ASAP7_75t_L g5282 ( 
.A(n_5218),
.Y(n_5282)
);

OAI211xp5_ASAP7_75t_L g5283 ( 
.A1(n_5105),
.A2(n_5042),
.B(n_5017),
.C(n_4998),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_5153),
.Y(n_5284)
);

AND2x2_ASAP7_75t_L g5285 ( 
.A(n_5144),
.B(n_5216),
.Y(n_5285)
);

AND2x2_ASAP7_75t_L g5286 ( 
.A(n_5212),
.B(n_5052),
.Y(n_5286)
);

AOI22xp33_ASAP7_75t_L g5287 ( 
.A1(n_5260),
.A2(n_4995),
.B1(n_5094),
.B2(n_5097),
.Y(n_5287)
);

NAND2xp5_ASAP7_75t_L g5288 ( 
.A(n_5227),
.B(n_5091),
.Y(n_5288)
);

INVx5_ASAP7_75t_L g5289 ( 
.A(n_5218),
.Y(n_5289)
);

AOI22xp33_ASAP7_75t_L g5290 ( 
.A1(n_5260),
.A2(n_5007),
.B1(n_4984),
.B2(n_4924),
.Y(n_5290)
);

BUFx4f_ASAP7_75t_SL g5291 ( 
.A(n_5110),
.Y(n_5291)
);

AOI22xp33_ASAP7_75t_SL g5292 ( 
.A1(n_5254),
.A2(n_4923),
.B1(n_5080),
.B2(n_5009),
.Y(n_5292)
);

OAI211xp5_ASAP7_75t_L g5293 ( 
.A1(n_5256),
.A2(n_5071),
.B(n_4977),
.C(n_4971),
.Y(n_5293)
);

OAI22xp33_ASAP7_75t_L g5294 ( 
.A1(n_5256),
.A2(n_5002),
.B1(n_4934),
.B2(n_5103),
.Y(n_5294)
);

INVx1_ASAP7_75t_SL g5295 ( 
.A(n_5217),
.Y(n_5295)
);

AOI222xp33_ASAP7_75t_L g5296 ( 
.A1(n_5203),
.A2(n_5032),
.B1(n_5057),
.B2(n_5060),
.C1(n_5084),
.C2(n_5086),
.Y(n_5296)
);

OAI211xp5_ASAP7_75t_L g5297 ( 
.A1(n_5135),
.A2(n_5082),
.B(n_4945),
.C(n_4989),
.Y(n_5297)
);

AOI22xp5_ASAP7_75t_L g5298 ( 
.A1(n_5223),
.A2(n_4906),
.B1(n_4992),
.B2(n_5036),
.Y(n_5298)
);

AOI22xp33_ASAP7_75t_L g5299 ( 
.A1(n_5251),
.A2(n_4956),
.B1(n_5030),
.B2(n_5013),
.Y(n_5299)
);

INVx1_ASAP7_75t_L g5300 ( 
.A(n_5154),
.Y(n_5300)
);

OAI22xp5_ASAP7_75t_L g5301 ( 
.A1(n_5241),
.A2(n_249),
.B1(n_245),
.B2(n_248),
.Y(n_5301)
);

INVx2_ASAP7_75t_L g5302 ( 
.A(n_5131),
.Y(n_5302)
);

AOI221xp5_ASAP7_75t_L g5303 ( 
.A1(n_5227),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.C(n_251),
.Y(n_5303)
);

AOI22xp33_ASAP7_75t_SL g5304 ( 
.A1(n_5249),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_5304)
);

AOI22xp33_ASAP7_75t_L g5305 ( 
.A1(n_5251),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_5305)
);

AOI22xp33_ASAP7_75t_L g5306 ( 
.A1(n_5176),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_5306)
);

NAND2xp5_ASAP7_75t_L g5307 ( 
.A(n_5167),
.B(n_5158),
.Y(n_5307)
);

AOI221xp5_ASAP7_75t_L g5308 ( 
.A1(n_5160),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.C(n_262),
.Y(n_5308)
);

NAND2xp5_ASAP7_75t_L g5309 ( 
.A(n_5244),
.B(n_259),
.Y(n_5309)
);

INVx4_ASAP7_75t_SL g5310 ( 
.A(n_5218),
.Y(n_5310)
);

AND2x2_ASAP7_75t_L g5311 ( 
.A(n_5142),
.B(n_261),
.Y(n_5311)
);

OAI22xp5_ASAP7_75t_L g5312 ( 
.A1(n_5241),
.A2(n_267),
.B1(n_263),
.B2(n_264),
.Y(n_5312)
);

OAI211xp5_ASAP7_75t_L g5313 ( 
.A1(n_5166),
.A2(n_267),
.B(n_263),
.C(n_264),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_5131),
.Y(n_5314)
);

OR2x2_ASAP7_75t_L g5315 ( 
.A(n_5106),
.B(n_268),
.Y(n_5315)
);

OR2x2_ASAP7_75t_L g5316 ( 
.A(n_5195),
.B(n_270),
.Y(n_5316)
);

OAI22xp33_ASAP7_75t_L g5317 ( 
.A1(n_5222),
.A2(n_5197),
.B1(n_5132),
.B2(n_5165),
.Y(n_5317)
);

AOI22xp33_ASAP7_75t_L g5318 ( 
.A1(n_5210),
.A2(n_276),
.B1(n_273),
.B2(n_275),
.Y(n_5318)
);

OA21x2_ASAP7_75t_L g5319 ( 
.A1(n_5174),
.A2(n_5193),
.B(n_5175),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_5128),
.Y(n_5320)
);

INVx2_ASAP7_75t_L g5321 ( 
.A(n_5116),
.Y(n_5321)
);

AOI22xp33_ASAP7_75t_L g5322 ( 
.A1(n_5211),
.A2(n_276),
.B1(n_273),
.B2(n_275),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_5129),
.Y(n_5323)
);

OAI22xp5_ASAP7_75t_L g5324 ( 
.A1(n_5160),
.A2(n_281),
.B1(n_278),
.B2(n_280),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_5120),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_5185),
.B(n_278),
.Y(n_5326)
);

INVx3_ASAP7_75t_L g5327 ( 
.A(n_5111),
.Y(n_5327)
);

AOI22xp33_ASAP7_75t_L g5328 ( 
.A1(n_5224),
.A2(n_284),
.B1(n_280),
.B2(n_283),
.Y(n_5328)
);

AOI21xp5_ASAP7_75t_L g5329 ( 
.A1(n_5207),
.A2(n_284),
.B(n_285),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5120),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_5107),
.Y(n_5331)
);

AOI21x1_ASAP7_75t_L g5332 ( 
.A1(n_5230),
.A2(n_286),
.B(n_287),
.Y(n_5332)
);

INVx1_ASAP7_75t_L g5333 ( 
.A(n_5113),
.Y(n_5333)
);

OR2x2_ASAP7_75t_L g5334 ( 
.A(n_5195),
.B(n_287),
.Y(n_5334)
);

AOI22xp33_ASAP7_75t_L g5335 ( 
.A1(n_5215),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.Y(n_5335)
);

INVx2_ASAP7_75t_L g5336 ( 
.A(n_5116),
.Y(n_5336)
);

OAI22xp5_ASAP7_75t_L g5337 ( 
.A1(n_5222),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_5119),
.Y(n_5338)
);

OAI22xp5_ASAP7_75t_SL g5339 ( 
.A1(n_5231),
.A2(n_295),
.B1(n_291),
.B2(n_294),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5115),
.Y(n_5340)
);

AOI22xp33_ASAP7_75t_L g5341 ( 
.A1(n_5240),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_5188),
.B(n_296),
.Y(n_5342)
);

OAI31xp33_ASAP7_75t_L g5343 ( 
.A1(n_5207),
.A2(n_299),
.A3(n_297),
.B(n_298),
.Y(n_5343)
);

AOI22xp33_ASAP7_75t_L g5344 ( 
.A1(n_5196),
.A2(n_301),
.B1(n_298),
.B2(n_300),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_5121),
.Y(n_5345)
);

AOI221xp5_ASAP7_75t_L g5346 ( 
.A1(n_5174),
.A2(n_306),
.B1(n_302),
.B2(n_303),
.C(n_307),
.Y(n_5346)
);

AND2x2_ASAP7_75t_L g5347 ( 
.A(n_5162),
.B(n_302),
.Y(n_5347)
);

AOI22xp33_ASAP7_75t_L g5348 ( 
.A1(n_5214),
.A2(n_309),
.B1(n_306),
.B2(n_308),
.Y(n_5348)
);

AOI221xp5_ASAP7_75t_L g5349 ( 
.A1(n_5204),
.A2(n_312),
.B1(n_309),
.B2(n_310),
.C(n_313),
.Y(n_5349)
);

BUFx5_ASAP7_75t_L g5350 ( 
.A(n_5209),
.Y(n_5350)
);

HB1xp67_ASAP7_75t_L g5351 ( 
.A(n_5114),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5122),
.Y(n_5352)
);

AOI21xp5_ASAP7_75t_L g5353 ( 
.A1(n_5132),
.A2(n_310),
.B(n_312),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5123),
.Y(n_5354)
);

OR2x2_ASAP7_75t_L g5355 ( 
.A(n_5170),
.B(n_315),
.Y(n_5355)
);

AOI22xp33_ASAP7_75t_L g5356 ( 
.A1(n_5222),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_5356)
);

OAI22xp5_ASAP7_75t_L g5357 ( 
.A1(n_5165),
.A2(n_5236),
.B1(n_5238),
.B2(n_5197),
.Y(n_5357)
);

OAI211xp5_ASAP7_75t_L g5358 ( 
.A1(n_5247),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_5358)
);

NAND2xp5_ASAP7_75t_L g5359 ( 
.A(n_5177),
.B(n_319),
.Y(n_5359)
);

AOI22xp33_ASAP7_75t_L g5360 ( 
.A1(n_5197),
.A2(n_5235),
.B1(n_5198),
.B2(n_5192),
.Y(n_5360)
);

AOI22xp33_ASAP7_75t_SL g5361 ( 
.A1(n_5247),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_5361)
);

NAND2xp5_ASAP7_75t_L g5362 ( 
.A(n_5147),
.B(n_320),
.Y(n_5362)
);

OAI22xp5_ASAP7_75t_L g5363 ( 
.A1(n_5257),
.A2(n_5148),
.B1(n_5201),
.B2(n_5169),
.Y(n_5363)
);

AND2x4_ASAP7_75t_L g5364 ( 
.A(n_5156),
.B(n_321),
.Y(n_5364)
);

INVx2_ASAP7_75t_L g5365 ( 
.A(n_5119),
.Y(n_5365)
);

INVx1_ASAP7_75t_L g5366 ( 
.A(n_5124),
.Y(n_5366)
);

AOI22xp33_ASAP7_75t_L g5367 ( 
.A1(n_5148),
.A2(n_5252),
.B1(n_5156),
.B2(n_5184),
.Y(n_5367)
);

AOI22xp33_ASAP7_75t_L g5368 ( 
.A1(n_5252),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_5368)
);

AND2x2_ASAP7_75t_L g5369 ( 
.A(n_5164),
.B(n_325),
.Y(n_5369)
);

HB1xp67_ASAP7_75t_L g5370 ( 
.A(n_5136),
.Y(n_5370)
);

AOI221xp5_ASAP7_75t_L g5371 ( 
.A1(n_5168),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.C(n_329),
.Y(n_5371)
);

AOI221xp5_ASAP7_75t_L g5372 ( 
.A1(n_5168),
.A2(n_330),
.B1(n_326),
.B2(n_329),
.C(n_331),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_5139),
.B(n_330),
.Y(n_5373)
);

AOI22xp33_ASAP7_75t_L g5374 ( 
.A1(n_5182),
.A2(n_338),
.B1(n_332),
.B2(n_334),
.Y(n_5374)
);

INVx3_ASAP7_75t_L g5375 ( 
.A(n_5111),
.Y(n_5375)
);

OAI22xp5_ASAP7_75t_L g5376 ( 
.A1(n_5259),
.A2(n_340),
.B1(n_332),
.B2(n_338),
.Y(n_5376)
);

OAI22xp33_ASAP7_75t_L g5377 ( 
.A1(n_5149),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_5377)
);

OAI22xp5_ASAP7_75t_L g5378 ( 
.A1(n_5259),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_5378)
);

AOI22xp33_ASAP7_75t_L g5379 ( 
.A1(n_5220),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_5379)
);

BUFx2_ASAP7_75t_L g5380 ( 
.A(n_5179),
.Y(n_5380)
);

AOI22xp33_ASAP7_75t_L g5381 ( 
.A1(n_5199),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_5381)
);

HB1xp67_ASAP7_75t_L g5382 ( 
.A(n_5136),
.Y(n_5382)
);

AOI22xp33_ASAP7_75t_L g5383 ( 
.A1(n_5149),
.A2(n_351),
.B1(n_349),
.B2(n_350),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_5126),
.Y(n_5384)
);

NAND2xp5_ASAP7_75t_L g5385 ( 
.A(n_5141),
.B(n_352),
.Y(n_5385)
);

CKINVDCx5p33_ASAP7_75t_R g5386 ( 
.A(n_5110),
.Y(n_5386)
);

INVx5_ASAP7_75t_L g5387 ( 
.A(n_5150),
.Y(n_5387)
);

AOI22xp33_ASAP7_75t_L g5388 ( 
.A1(n_5150),
.A2(n_357),
.B1(n_353),
.B2(n_355),
.Y(n_5388)
);

AOI22xp33_ASAP7_75t_L g5389 ( 
.A1(n_5150),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_5389)
);

INVx4_ASAP7_75t_L g5390 ( 
.A(n_5171),
.Y(n_5390)
);

HB1xp67_ASAP7_75t_L g5391 ( 
.A(n_5138),
.Y(n_5391)
);

AOI22xp33_ASAP7_75t_L g5392 ( 
.A1(n_5206),
.A2(n_361),
.B1(n_358),
.B2(n_360),
.Y(n_5392)
);

OAI22xp5_ASAP7_75t_L g5393 ( 
.A1(n_5255),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_5393)
);

AOI22xp33_ASAP7_75t_L g5394 ( 
.A1(n_5206),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_5394)
);

OAI22xp5_ASAP7_75t_L g5395 ( 
.A1(n_5255),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_5395)
);

HB1xp67_ASAP7_75t_L g5396 ( 
.A(n_5138),
.Y(n_5396)
);

OAI22xp5_ASAP7_75t_L g5397 ( 
.A1(n_5206),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_5397)
);

OAI221xp5_ASAP7_75t_L g5398 ( 
.A1(n_5191),
.A2(n_372),
.B1(n_369),
.B2(n_371),
.C(n_373),
.Y(n_5398)
);

OAI22xp5_ASAP7_75t_L g5399 ( 
.A1(n_5181),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_5399)
);

AOI22xp33_ASAP7_75t_L g5400 ( 
.A1(n_5231),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_5400)
);

NAND2xp5_ASAP7_75t_L g5401 ( 
.A(n_5288),
.B(n_5133),
.Y(n_5401)
);

AND2x2_ASAP7_75t_L g5402 ( 
.A(n_5360),
.B(n_5137),
.Y(n_5402)
);

AND2x4_ASAP7_75t_L g5403 ( 
.A(n_5390),
.B(n_5171),
.Y(n_5403)
);

INVx2_ASAP7_75t_L g5404 ( 
.A(n_5350),
.Y(n_5404)
);

AND2x4_ASAP7_75t_SL g5405 ( 
.A(n_5390),
.B(n_5194),
.Y(n_5405)
);

AND2x2_ASAP7_75t_L g5406 ( 
.A(n_5285),
.B(n_5137),
.Y(n_5406)
);

AND2x2_ASAP7_75t_L g5407 ( 
.A(n_5265),
.B(n_5146),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5320),
.Y(n_5408)
);

AND2x4_ASAP7_75t_L g5409 ( 
.A(n_5325),
.B(n_5171),
.Y(n_5409)
);

AND2x2_ASAP7_75t_L g5410 ( 
.A(n_5380),
.B(n_5146),
.Y(n_5410)
);

AND2x4_ASAP7_75t_L g5411 ( 
.A(n_5330),
.B(n_5178),
.Y(n_5411)
);

NAND2xp5_ASAP7_75t_L g5412 ( 
.A(n_5263),
.B(n_5109),
.Y(n_5412)
);

AND2x2_ASAP7_75t_L g5413 ( 
.A(n_5286),
.B(n_5183),
.Y(n_5413)
);

AOI22xp5_ASAP7_75t_L g5414 ( 
.A1(n_5262),
.A2(n_5266),
.B1(n_5283),
.B2(n_5267),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5323),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5264),
.Y(n_5416)
);

OR2x2_ASAP7_75t_L g5417 ( 
.A(n_5270),
.B(n_5152),
.Y(n_5417)
);

AND2x2_ASAP7_75t_L g5418 ( 
.A(n_5367),
.B(n_5112),
.Y(n_5418)
);

INVx2_ASAP7_75t_L g5419 ( 
.A(n_5350),
.Y(n_5419)
);

AND2x2_ASAP7_75t_L g5420 ( 
.A(n_5363),
.B(n_5112),
.Y(n_5420)
);

AND2x2_ASAP7_75t_SL g5421 ( 
.A(n_5268),
.B(n_5194),
.Y(n_5421)
);

INVx2_ASAP7_75t_L g5422 ( 
.A(n_5319),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_5276),
.B(n_5118),
.Y(n_5423)
);

HB1xp67_ASAP7_75t_L g5424 ( 
.A(n_5319),
.Y(n_5424)
);

NOR2x1p5_ASAP7_75t_L g5425 ( 
.A(n_5279),
.B(n_5178),
.Y(n_5425)
);

INVx2_ASAP7_75t_L g5426 ( 
.A(n_5302),
.Y(n_5426)
);

AND2x2_ASAP7_75t_L g5427 ( 
.A(n_5357),
.B(n_5151),
.Y(n_5427)
);

AOI22xp33_ASAP7_75t_L g5428 ( 
.A1(n_5280),
.A2(n_5225),
.B1(n_5237),
.B2(n_5202),
.Y(n_5428)
);

INVx3_ASAP7_75t_L g5429 ( 
.A(n_5289),
.Y(n_5429)
);

BUFx2_ASAP7_75t_L g5430 ( 
.A(n_5289),
.Y(n_5430)
);

NAND2x1p5_ASAP7_75t_L g5431 ( 
.A(n_5387),
.B(n_5186),
.Y(n_5431)
);

INVx2_ASAP7_75t_L g5432 ( 
.A(n_5314),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_5274),
.Y(n_5433)
);

OR2x2_ASAP7_75t_L g5434 ( 
.A(n_5307),
.B(n_5159),
.Y(n_5434)
);

BUFx3_ASAP7_75t_L g5435 ( 
.A(n_5289),
.Y(n_5435)
);

HB1xp67_ASAP7_75t_L g5436 ( 
.A(n_5370),
.Y(n_5436)
);

NOR2xp33_ASAP7_75t_L g5437 ( 
.A(n_5295),
.B(n_5239),
.Y(n_5437)
);

AND2x2_ASAP7_75t_L g5438 ( 
.A(n_5351),
.B(n_5151),
.Y(n_5438)
);

INVx2_ASAP7_75t_L g5439 ( 
.A(n_5321),
.Y(n_5439)
);

AND2x2_ASAP7_75t_L g5440 ( 
.A(n_5364),
.B(n_5155),
.Y(n_5440)
);

NOR2xp33_ASAP7_75t_R g5441 ( 
.A(n_5332),
.B(n_5243),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_5284),
.Y(n_5442)
);

OR2x2_ASAP7_75t_L g5443 ( 
.A(n_5355),
.B(n_5271),
.Y(n_5443)
);

AND2x2_ASAP7_75t_L g5444 ( 
.A(n_5364),
.B(n_5155),
.Y(n_5444)
);

INVx3_ASAP7_75t_L g5445 ( 
.A(n_5282),
.Y(n_5445)
);

INVx2_ASAP7_75t_L g5446 ( 
.A(n_5350),
.Y(n_5446)
);

INVxp67_ASAP7_75t_SL g5447 ( 
.A(n_5273),
.Y(n_5447)
);

INVx2_ASAP7_75t_L g5448 ( 
.A(n_5350),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_5300),
.Y(n_5449)
);

NAND2xp5_ASAP7_75t_SL g5450 ( 
.A(n_5317),
.B(n_5186),
.Y(n_5450)
);

INVx2_ASAP7_75t_L g5451 ( 
.A(n_5350),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_L g5452 ( 
.A(n_5331),
.B(n_5125),
.Y(n_5452)
);

INVx4_ASAP7_75t_L g5453 ( 
.A(n_5387),
.Y(n_5453)
);

HB1xp67_ASAP7_75t_L g5454 ( 
.A(n_5382),
.Y(n_5454)
);

AND2x2_ASAP7_75t_L g5455 ( 
.A(n_5327),
.B(n_5200),
.Y(n_5455)
);

INVx3_ASAP7_75t_L g5456 ( 
.A(n_5282),
.Y(n_5456)
);

NAND2xp5_ASAP7_75t_L g5457 ( 
.A(n_5333),
.B(n_5130),
.Y(n_5457)
);

NAND2xp5_ASAP7_75t_L g5458 ( 
.A(n_5340),
.B(n_5143),
.Y(n_5458)
);

INVxp67_ASAP7_75t_L g5459 ( 
.A(n_5316),
.Y(n_5459)
);

AND2x2_ASAP7_75t_L g5460 ( 
.A(n_5327),
.B(n_5200),
.Y(n_5460)
);

INVx1_ASAP7_75t_SL g5461 ( 
.A(n_5291),
.Y(n_5461)
);

OR2x2_ASAP7_75t_L g5462 ( 
.A(n_5334),
.B(n_5145),
.Y(n_5462)
);

AND2x2_ASAP7_75t_L g5463 ( 
.A(n_5375),
.B(n_5208),
.Y(n_5463)
);

AND2x2_ASAP7_75t_L g5464 ( 
.A(n_5375),
.B(n_5208),
.Y(n_5464)
);

INVx2_ASAP7_75t_L g5465 ( 
.A(n_5336),
.Y(n_5465)
);

AND2x4_ASAP7_75t_L g5466 ( 
.A(n_5387),
.B(n_5253),
.Y(n_5466)
);

CKINVDCx20_ASAP7_75t_R g5467 ( 
.A(n_5386),
.Y(n_5467)
);

INVx2_ASAP7_75t_L g5468 ( 
.A(n_5282),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_5338),
.Y(n_5469)
);

AND2x2_ASAP7_75t_L g5470 ( 
.A(n_5278),
.B(n_5226),
.Y(n_5470)
);

NAND2xp5_ASAP7_75t_L g5471 ( 
.A(n_5345),
.B(n_5140),
.Y(n_5471)
);

INVx2_ASAP7_75t_SL g5472 ( 
.A(n_5310),
.Y(n_5472)
);

INVx2_ASAP7_75t_L g5473 ( 
.A(n_5365),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5352),
.Y(n_5474)
);

NAND2xp5_ASAP7_75t_L g5475 ( 
.A(n_5354),
.B(n_5140),
.Y(n_5475)
);

AND2x2_ASAP7_75t_L g5476 ( 
.A(n_5278),
.B(n_5226),
.Y(n_5476)
);

INVx2_ASAP7_75t_L g5477 ( 
.A(n_5366),
.Y(n_5477)
);

OR2x2_ASAP7_75t_L g5478 ( 
.A(n_5384),
.B(n_5161),
.Y(n_5478)
);

INVx2_ASAP7_75t_L g5479 ( 
.A(n_5391),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_5396),
.Y(n_5480)
);

INVx2_ASAP7_75t_L g5481 ( 
.A(n_5310),
.Y(n_5481)
);

OAI22xp33_ASAP7_75t_L g5482 ( 
.A1(n_5398),
.A2(n_5134),
.B1(n_5225),
.B2(n_5242),
.Y(n_5482)
);

HB1xp67_ASAP7_75t_L g5483 ( 
.A(n_5342),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_5373),
.Y(n_5484)
);

AND2x2_ASAP7_75t_L g5485 ( 
.A(n_5347),
.B(n_5242),
.Y(n_5485)
);

AND2x2_ASAP7_75t_L g5486 ( 
.A(n_5311),
.B(n_5108),
.Y(n_5486)
);

BUFx2_ASAP7_75t_L g5487 ( 
.A(n_5315),
.Y(n_5487)
);

AND2x4_ASAP7_75t_L g5488 ( 
.A(n_5369),
.B(n_5173),
.Y(n_5488)
);

INVx2_ASAP7_75t_L g5489 ( 
.A(n_5359),
.Y(n_5489)
);

OR2x2_ASAP7_75t_L g5490 ( 
.A(n_5326),
.B(n_5180),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5385),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5362),
.Y(n_5492)
);

NOR2xp33_ASAP7_75t_L g5493 ( 
.A(n_5358),
.B(n_5243),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_5309),
.Y(n_5494)
);

INVx2_ASAP7_75t_SL g5495 ( 
.A(n_5399),
.Y(n_5495)
);

OAI321xp33_ASAP7_75t_L g5496 ( 
.A1(n_5294),
.A2(n_5175),
.A3(n_5173),
.B1(n_5134),
.B2(n_5258),
.C(n_5221),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5298),
.Y(n_5497)
);

INVx2_ASAP7_75t_L g5498 ( 
.A(n_5337),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5305),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_5313),
.Y(n_5500)
);

INVx2_ASAP7_75t_L g5501 ( 
.A(n_5301),
.Y(n_5501)
);

OA21x2_ASAP7_75t_L g5502 ( 
.A1(n_5269),
.A2(n_5172),
.B(n_5117),
.Y(n_5502)
);

AOI221xp5_ASAP7_75t_L g5503 ( 
.A1(n_5308),
.A2(n_5202),
.B1(n_379),
.B2(n_377),
.C(n_378),
.Y(n_5503)
);

OR2x2_ASAP7_75t_L g5504 ( 
.A(n_5299),
.B(n_5353),
.Y(n_5504)
);

AOI22xp33_ASAP7_75t_L g5505 ( 
.A1(n_5272),
.A2(n_5213),
.B1(n_5234),
.B2(n_5250),
.Y(n_5505)
);

OR2x2_ASAP7_75t_L g5506 ( 
.A(n_5277),
.B(n_5189),
.Y(n_5506)
);

BUFx3_ASAP7_75t_L g5507 ( 
.A(n_5339),
.Y(n_5507)
);

NAND2xp5_ASAP7_75t_L g5508 ( 
.A(n_5303),
.B(n_5219),
.Y(n_5508)
);

INVx2_ASAP7_75t_L g5509 ( 
.A(n_5312),
.Y(n_5509)
);

AND2x2_ASAP7_75t_L g5510 ( 
.A(n_5292),
.B(n_378),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_5293),
.Y(n_5511)
);

INVx2_ASAP7_75t_L g5512 ( 
.A(n_5393),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_5395),
.Y(n_5513)
);

INVx2_ASAP7_75t_L g5514 ( 
.A(n_5324),
.Y(n_5514)
);

OAI221xp5_ASAP7_75t_L g5515 ( 
.A1(n_5447),
.A2(n_5343),
.B1(n_5361),
.B2(n_5304),
.C(n_5329),
.Y(n_5515)
);

INVx2_ASAP7_75t_L g5516 ( 
.A(n_5435),
.Y(n_5516)
);

AND4x1_ASAP7_75t_L g5517 ( 
.A(n_5503),
.B(n_5346),
.C(n_5372),
.D(n_5371),
.Y(n_5517)
);

HB1xp67_ASAP7_75t_L g5518 ( 
.A(n_5447),
.Y(n_5518)
);

OAI22xp5_ASAP7_75t_SL g5519 ( 
.A1(n_5507),
.A2(n_5328),
.B1(n_5287),
.B2(n_5368),
.Y(n_5519)
);

OAI22xp5_ASAP7_75t_L g5520 ( 
.A1(n_5414),
.A2(n_5290),
.B1(n_5306),
.B2(n_5281),
.Y(n_5520)
);

AOI221xp5_ASAP7_75t_L g5521 ( 
.A1(n_5511),
.A2(n_5349),
.B1(n_5377),
.B2(n_5397),
.C(n_5378),
.Y(n_5521)
);

OAI33xp33_ASAP7_75t_L g5522 ( 
.A1(n_5482),
.A2(n_5376),
.A3(n_5275),
.B1(n_5400),
.B2(n_5296),
.B3(n_5344),
.Y(n_5522)
);

OAI222xp33_ASAP7_75t_L g5523 ( 
.A1(n_5428),
.A2(n_5356),
.B1(n_5335),
.B2(n_5374),
.C1(n_5348),
.C2(n_5322),
.Y(n_5523)
);

BUFx12f_ASAP7_75t_L g5524 ( 
.A(n_5421),
.Y(n_5524)
);

AOI221xp5_ASAP7_75t_L g5525 ( 
.A1(n_5482),
.A2(n_5379),
.B1(n_5381),
.B2(n_5297),
.C(n_5318),
.Y(n_5525)
);

INVx2_ASAP7_75t_L g5526 ( 
.A(n_5435),
.Y(n_5526)
);

INVxp67_ASAP7_75t_L g5527 ( 
.A(n_5430),
.Y(n_5527)
);

OAI22xp5_ASAP7_75t_L g5528 ( 
.A1(n_5428),
.A2(n_5341),
.B1(n_5394),
.B2(n_5392),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_5497),
.B(n_5495),
.Y(n_5529)
);

OAI22xp33_ASAP7_75t_L g5530 ( 
.A1(n_5508),
.A2(n_5504),
.B1(n_5506),
.B2(n_5496),
.Y(n_5530)
);

NAND4xp25_ASAP7_75t_L g5531 ( 
.A(n_5503),
.B(n_5507),
.C(n_5505),
.D(n_5493),
.Y(n_5531)
);

AND2x4_ASAP7_75t_SL g5532 ( 
.A(n_5467),
.B(n_5383),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_5408),
.Y(n_5533)
);

AOI21xp33_ASAP7_75t_SL g5534 ( 
.A1(n_5421),
.A2(n_5389),
.B(n_5388),
.Y(n_5534)
);

OAI221xp5_ASAP7_75t_L g5535 ( 
.A1(n_5505),
.A2(n_384),
.B1(n_381),
.B2(n_382),
.C(n_387),
.Y(n_5535)
);

INVx2_ASAP7_75t_L g5536 ( 
.A(n_5429),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5415),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_5416),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_5433),
.Y(n_5539)
);

AND2x2_ASAP7_75t_L g5540 ( 
.A(n_5425),
.B(n_381),
.Y(n_5540)
);

OAI22xp33_ASAP7_75t_L g5541 ( 
.A1(n_5508),
.A2(n_389),
.B1(n_384),
.B2(n_388),
.Y(n_5541)
);

OA21x2_ASAP7_75t_L g5542 ( 
.A1(n_5424),
.A2(n_388),
.B(n_390),
.Y(n_5542)
);

AOI22xp33_ASAP7_75t_L g5543 ( 
.A1(n_5499),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_5543)
);

NOR2xp33_ASAP7_75t_L g5544 ( 
.A(n_5437),
.B(n_392),
.Y(n_5544)
);

AOI22xp33_ASAP7_75t_L g5545 ( 
.A1(n_5500),
.A2(n_397),
.B1(n_394),
.B2(n_396),
.Y(n_5545)
);

INVx2_ASAP7_75t_L g5546 ( 
.A(n_5429),
.Y(n_5546)
);

OAI31xp33_ASAP7_75t_SL g5547 ( 
.A1(n_5450),
.A2(n_5493),
.A3(n_5510),
.B(n_5441),
.Y(n_5547)
);

OAI22xp5_ASAP7_75t_L g5548 ( 
.A1(n_5412),
.A2(n_397),
.B1(n_394),
.B2(n_396),
.Y(n_5548)
);

AOI22xp33_ASAP7_75t_L g5549 ( 
.A1(n_5514),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_5549)
);

AND2x2_ASAP7_75t_L g5550 ( 
.A(n_5420),
.B(n_398),
.Y(n_5550)
);

NAND2x1p5_ASAP7_75t_L g5551 ( 
.A(n_5453),
.B(n_400),
.Y(n_5551)
);

OAI211xp5_ASAP7_75t_SL g5552 ( 
.A1(n_5459),
.A2(n_404),
.B(n_402),
.C(n_403),
.Y(n_5552)
);

AOI22xp5_ASAP7_75t_L g5553 ( 
.A1(n_5498),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_5553)
);

AOI22xp5_ASAP7_75t_L g5554 ( 
.A1(n_5498),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_5554)
);

INVx1_ASAP7_75t_L g5555 ( 
.A(n_5442),
.Y(n_5555)
);

AOI22xp33_ASAP7_75t_L g5556 ( 
.A1(n_5514),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_5556)
);

INVx2_ASAP7_75t_L g5557 ( 
.A(n_5453),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_5449),
.Y(n_5558)
);

NAND3xp33_ASAP7_75t_L g5559 ( 
.A(n_5412),
.B(n_5483),
.C(n_5459),
.Y(n_5559)
);

AOI22xp33_ASAP7_75t_L g5560 ( 
.A1(n_5513),
.A2(n_412),
.B1(n_409),
.B2(n_410),
.Y(n_5560)
);

AND2x4_ASAP7_75t_L g5561 ( 
.A(n_5409),
.B(n_409),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_5474),
.Y(n_5562)
);

AOI33xp33_ASAP7_75t_L g5563 ( 
.A1(n_5501),
.A2(n_412),
.A3(n_413),
.B1(n_414),
.B2(n_416),
.B3(n_417),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5477),
.Y(n_5564)
);

AOI221xp5_ASAP7_75t_L g5565 ( 
.A1(n_5441),
.A2(n_5501),
.B1(n_5513),
.B2(n_5509),
.C(n_5483),
.Y(n_5565)
);

AOI22xp33_ASAP7_75t_L g5566 ( 
.A1(n_5512),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_5566)
);

NAND4xp25_ASAP7_75t_L g5567 ( 
.A(n_5443),
.B(n_420),
.C(n_418),
.D(n_419),
.Y(n_5567)
);

NAND4xp25_ASAP7_75t_L g5568 ( 
.A(n_5450),
.B(n_422),
.C(n_420),
.D(n_421),
.Y(n_5568)
);

OAI22xp5_ASAP7_75t_L g5569 ( 
.A1(n_5409),
.A2(n_5401),
.B1(n_5487),
.B2(n_5431),
.Y(n_5569)
);

AND2x2_ASAP7_75t_L g5570 ( 
.A(n_5407),
.B(n_421),
.Y(n_5570)
);

NOR3xp33_ASAP7_75t_L g5571 ( 
.A(n_5437),
.B(n_422),
.C(n_423),
.Y(n_5571)
);

AOI22xp33_ASAP7_75t_L g5572 ( 
.A1(n_5402),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_5572)
);

BUFx3_ASAP7_75t_L g5573 ( 
.A(n_5467),
.Y(n_5573)
);

NAND3xp33_ASAP7_75t_L g5574 ( 
.A(n_5502),
.B(n_424),
.C(n_428),
.Y(n_5574)
);

HB1xp67_ASAP7_75t_L g5575 ( 
.A(n_5436),
.Y(n_5575)
);

AND2x2_ASAP7_75t_L g5576 ( 
.A(n_5410),
.B(n_429),
.Y(n_5576)
);

NAND2xp5_ASAP7_75t_L g5577 ( 
.A(n_5494),
.B(n_431),
.Y(n_5577)
);

NAND2xp5_ASAP7_75t_L g5578 ( 
.A(n_5494),
.B(n_5489),
.Y(n_5578)
);

NAND3xp33_ASAP7_75t_L g5579 ( 
.A(n_5424),
.B(n_432),
.C(n_433),
.Y(n_5579)
);

INVx2_ASAP7_75t_L g5580 ( 
.A(n_5481),
.Y(n_5580)
);

NAND2x1p5_ASAP7_75t_L g5581 ( 
.A(n_5403),
.B(n_432),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_5472),
.Y(n_5582)
);

OR2x2_ASAP7_75t_L g5583 ( 
.A(n_5492),
.B(n_433),
.Y(n_5583)
);

INVx2_ASAP7_75t_L g5584 ( 
.A(n_5445),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_5436),
.Y(n_5585)
);

OAI21xp5_ASAP7_75t_L g5586 ( 
.A1(n_5423),
.A2(n_434),
.B(n_435),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5454),
.Y(n_5587)
);

AOI221xp5_ASAP7_75t_L g5588 ( 
.A1(n_5492),
.A2(n_434),
.B1(n_436),
.B2(n_440),
.C(n_441),
.Y(n_5588)
);

AND2x2_ASAP7_75t_L g5589 ( 
.A(n_5427),
.B(n_441),
.Y(n_5589)
);

AND2x2_ASAP7_75t_L g5590 ( 
.A(n_5468),
.B(n_442),
.Y(n_5590)
);

INVx2_ASAP7_75t_L g5591 ( 
.A(n_5582),
.Y(n_5591)
);

AND2x2_ASAP7_75t_L g5592 ( 
.A(n_5516),
.B(n_5403),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5575),
.Y(n_5593)
);

AND2x2_ASAP7_75t_L g5594 ( 
.A(n_5526),
.B(n_5431),
.Y(n_5594)
);

INVx2_ASAP7_75t_L g5595 ( 
.A(n_5561),
.Y(n_5595)
);

OR2x2_ASAP7_75t_L g5596 ( 
.A(n_5518),
.B(n_5454),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_5585),
.Y(n_5597)
);

AND2x2_ASAP7_75t_L g5598 ( 
.A(n_5527),
.B(n_5418),
.Y(n_5598)
);

NAND2xp5_ASAP7_75t_L g5599 ( 
.A(n_5541),
.B(n_5489),
.Y(n_5599)
);

AND2x2_ASAP7_75t_L g5600 ( 
.A(n_5557),
.B(n_5580),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_5542),
.Y(n_5601)
);

INVx2_ASAP7_75t_L g5602 ( 
.A(n_5561),
.Y(n_5602)
);

INVx2_ASAP7_75t_L g5603 ( 
.A(n_5542),
.Y(n_5603)
);

AND2x4_ASAP7_75t_L g5604 ( 
.A(n_5536),
.B(n_5405),
.Y(n_5604)
);

AND2x2_ASAP7_75t_L g5605 ( 
.A(n_5546),
.B(n_5405),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5587),
.Y(n_5606)
);

NOR2xp33_ASAP7_75t_L g5607 ( 
.A(n_5573),
.B(n_5461),
.Y(n_5607)
);

INVx2_ASAP7_75t_L g5608 ( 
.A(n_5581),
.Y(n_5608)
);

AND2x2_ASAP7_75t_L g5609 ( 
.A(n_5584),
.B(n_5479),
.Y(n_5609)
);

AOI22xp33_ASAP7_75t_L g5610 ( 
.A1(n_5531),
.A2(n_5502),
.B1(n_5484),
.B2(n_5491),
.Y(n_5610)
);

NAND2xp5_ASAP7_75t_L g5611 ( 
.A(n_5565),
.B(n_5547),
.Y(n_5611)
);

AND2x2_ASAP7_75t_L g5612 ( 
.A(n_5529),
.B(n_5445),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_5578),
.Y(n_5613)
);

NAND2xp5_ASAP7_75t_L g5614 ( 
.A(n_5589),
.B(n_5401),
.Y(n_5614)
);

OR2x2_ASAP7_75t_L g5615 ( 
.A(n_5559),
.B(n_5564),
.Y(n_5615)
);

INVx3_ASAP7_75t_L g5616 ( 
.A(n_5524),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5533),
.Y(n_5617)
);

INVx1_ASAP7_75t_L g5618 ( 
.A(n_5537),
.Y(n_5618)
);

NAND2xp5_ASAP7_75t_L g5619 ( 
.A(n_5550),
.B(n_5456),
.Y(n_5619)
);

INVx2_ASAP7_75t_L g5620 ( 
.A(n_5551),
.Y(n_5620)
);

AND2x4_ASAP7_75t_L g5621 ( 
.A(n_5574),
.B(n_5456),
.Y(n_5621)
);

AND2x2_ASAP7_75t_L g5622 ( 
.A(n_5569),
.B(n_5411),
.Y(n_5622)
);

AND2x2_ASAP7_75t_L g5623 ( 
.A(n_5570),
.B(n_5411),
.Y(n_5623)
);

NOR2xp33_ASAP7_75t_L g5624 ( 
.A(n_5522),
.B(n_5462),
.Y(n_5624)
);

INVx1_ASAP7_75t_L g5625 ( 
.A(n_5538),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5539),
.Y(n_5626)
);

AND2x2_ASAP7_75t_L g5627 ( 
.A(n_5576),
.B(n_5455),
.Y(n_5627)
);

NAND2xp5_ASAP7_75t_L g5628 ( 
.A(n_5530),
.B(n_5423),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5583),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_L g5630 ( 
.A(n_5525),
.B(n_5480),
.Y(n_5630)
);

INVx2_ASAP7_75t_L g5631 ( 
.A(n_5540),
.Y(n_5631)
);

AND2x2_ASAP7_75t_L g5632 ( 
.A(n_5555),
.B(n_5460),
.Y(n_5632)
);

AND2x2_ASAP7_75t_L g5633 ( 
.A(n_5558),
.B(n_5463),
.Y(n_5633)
);

INVx1_ASAP7_75t_L g5634 ( 
.A(n_5562),
.Y(n_5634)
);

AND2x4_ASAP7_75t_SL g5635 ( 
.A(n_5571),
.B(n_5413),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5579),
.Y(n_5636)
);

INVxp67_ASAP7_75t_SL g5637 ( 
.A(n_5579),
.Y(n_5637)
);

AND2x2_ASAP7_75t_L g5638 ( 
.A(n_5590),
.B(n_5464),
.Y(n_5638)
);

INVx2_ASAP7_75t_L g5639 ( 
.A(n_5577),
.Y(n_5639)
);

INVx1_ASAP7_75t_L g5640 ( 
.A(n_5596),
.Y(n_5640)
);

AND2x2_ASAP7_75t_L g5641 ( 
.A(n_5592),
.B(n_5470),
.Y(n_5641)
);

INVx2_ASAP7_75t_L g5642 ( 
.A(n_5596),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_5593),
.Y(n_5643)
);

AO22x1_ASAP7_75t_L g5644 ( 
.A1(n_5637),
.A2(n_5586),
.B1(n_5544),
.B2(n_5548),
.Y(n_5644)
);

INVx2_ASAP7_75t_L g5645 ( 
.A(n_5608),
.Y(n_5645)
);

INVx1_ASAP7_75t_L g5646 ( 
.A(n_5593),
.Y(n_5646)
);

AOI211xp5_ASAP7_75t_L g5647 ( 
.A1(n_5611),
.A2(n_5515),
.B(n_5535),
.C(n_5568),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_5606),
.Y(n_5648)
);

AND2x2_ASAP7_75t_L g5649 ( 
.A(n_5592),
.B(n_5476),
.Y(n_5649)
);

BUFx12f_ASAP7_75t_L g5650 ( 
.A(n_5621),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_5606),
.Y(n_5651)
);

NAND3xp33_ASAP7_75t_L g5652 ( 
.A(n_5610),
.B(n_5517),
.C(n_5588),
.Y(n_5652)
);

INVx2_ASAP7_75t_L g5653 ( 
.A(n_5608),
.Y(n_5653)
);

INVx2_ASAP7_75t_L g5654 ( 
.A(n_5620),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_5620),
.Y(n_5655)
);

AND2x2_ASAP7_75t_L g5656 ( 
.A(n_5616),
.B(n_5466),
.Y(n_5656)
);

AND2x2_ASAP7_75t_L g5657 ( 
.A(n_5616),
.B(n_5466),
.Y(n_5657)
);

OR2x2_ASAP7_75t_L g5658 ( 
.A(n_5636),
.B(n_5426),
.Y(n_5658)
);

INVx2_ASAP7_75t_L g5659 ( 
.A(n_5595),
.Y(n_5659)
);

AND2x2_ASAP7_75t_L g5660 ( 
.A(n_5616),
.B(n_5440),
.Y(n_5660)
);

AOI33xp33_ASAP7_75t_L g5661 ( 
.A1(n_5636),
.A2(n_5545),
.A3(n_5556),
.B1(n_5549),
.B2(n_5543),
.B3(n_5572),
.Y(n_5661)
);

AND2x4_ASAP7_75t_L g5662 ( 
.A(n_5604),
.B(n_5422),
.Y(n_5662)
);

OAI211xp5_ASAP7_75t_L g5663 ( 
.A1(n_5628),
.A2(n_5534),
.B(n_5567),
.C(n_5521),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5618),
.Y(n_5664)
);

INVx2_ASAP7_75t_L g5665 ( 
.A(n_5595),
.Y(n_5665)
);

OR2x2_ASAP7_75t_L g5666 ( 
.A(n_5603),
.B(n_5426),
.Y(n_5666)
);

AOI22xp33_ASAP7_75t_L g5667 ( 
.A1(n_5624),
.A2(n_5519),
.B1(n_5520),
.B2(n_5528),
.Y(n_5667)
);

AND2x2_ASAP7_75t_L g5668 ( 
.A(n_5623),
.B(n_5444),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_5618),
.Y(n_5669)
);

AND2x2_ASAP7_75t_L g5670 ( 
.A(n_5623),
.B(n_5438),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_5626),
.Y(n_5671)
);

NAND4xp25_ASAP7_75t_SL g5672 ( 
.A(n_5630),
.B(n_5534),
.C(n_5563),
.D(n_5554),
.Y(n_5672)
);

AND2x2_ASAP7_75t_L g5673 ( 
.A(n_5656),
.B(n_5605),
.Y(n_5673)
);

AND2x2_ASAP7_75t_L g5674 ( 
.A(n_5656),
.B(n_5605),
.Y(n_5674)
);

INVx1_ASAP7_75t_SL g5675 ( 
.A(n_5650),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5642),
.Y(n_5676)
);

HB1xp67_ASAP7_75t_L g5677 ( 
.A(n_5650),
.Y(n_5677)
);

AND2x2_ASAP7_75t_L g5678 ( 
.A(n_5657),
.B(n_5627),
.Y(n_5678)
);

OR2x2_ASAP7_75t_L g5679 ( 
.A(n_5645),
.B(n_5602),
.Y(n_5679)
);

AND2x4_ASAP7_75t_L g5680 ( 
.A(n_5657),
.B(n_5602),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_L g5681 ( 
.A(n_5652),
.B(n_5601),
.Y(n_5681)
);

INVx2_ASAP7_75t_L g5682 ( 
.A(n_5662),
.Y(n_5682)
);

BUFx2_ASAP7_75t_L g5683 ( 
.A(n_5662),
.Y(n_5683)
);

OAI21xp33_ASAP7_75t_L g5684 ( 
.A1(n_5667),
.A2(n_5663),
.B(n_5672),
.Y(n_5684)
);

INVx2_ASAP7_75t_L g5685 ( 
.A(n_5662),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_5642),
.Y(n_5686)
);

INVx1_ASAP7_75t_L g5687 ( 
.A(n_5659),
.Y(n_5687)
);

AND2x2_ASAP7_75t_L g5688 ( 
.A(n_5641),
.B(n_5627),
.Y(n_5688)
);

OR2x2_ASAP7_75t_L g5689 ( 
.A(n_5645),
.B(n_5599),
.Y(n_5689)
);

OR2x6_ASAP7_75t_L g5690 ( 
.A(n_5644),
.B(n_5631),
.Y(n_5690)
);

NAND2xp5_ASAP7_75t_L g5691 ( 
.A(n_5647),
.B(n_5640),
.Y(n_5691)
);

AND2x2_ASAP7_75t_L g5692 ( 
.A(n_5641),
.B(n_5598),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5659),
.Y(n_5693)
);

BUFx3_ASAP7_75t_L g5694 ( 
.A(n_5665),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_L g5695 ( 
.A(n_5665),
.B(n_5601),
.Y(n_5695)
);

INVx2_ASAP7_75t_L g5696 ( 
.A(n_5683),
.Y(n_5696)
);

AND2x2_ASAP7_75t_L g5697 ( 
.A(n_5692),
.B(n_5649),
.Y(n_5697)
);

NAND3xp33_ASAP7_75t_L g5698 ( 
.A(n_5690),
.B(n_5603),
.C(n_5517),
.Y(n_5698)
);

INVx1_ASAP7_75t_SL g5699 ( 
.A(n_5690),
.Y(n_5699)
);

AND2x2_ASAP7_75t_L g5700 ( 
.A(n_5678),
.B(n_5649),
.Y(n_5700)
);

NOR2xp33_ASAP7_75t_L g5701 ( 
.A(n_5675),
.B(n_5660),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5694),
.Y(n_5702)
);

NAND2xp5_ASAP7_75t_L g5703 ( 
.A(n_5688),
.B(n_5631),
.Y(n_5703)
);

INVx1_ASAP7_75t_L g5704 ( 
.A(n_5694),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_5679),
.Y(n_5705)
);

NAND2xp5_ASAP7_75t_L g5706 ( 
.A(n_5684),
.B(n_5653),
.Y(n_5706)
);

INVxp67_ASAP7_75t_L g5707 ( 
.A(n_5690),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5682),
.Y(n_5708)
);

INVx2_ASAP7_75t_SL g5709 ( 
.A(n_5680),
.Y(n_5709)
);

NAND2xp5_ASAP7_75t_L g5710 ( 
.A(n_5681),
.B(n_5653),
.Y(n_5710)
);

AND2x2_ASAP7_75t_L g5711 ( 
.A(n_5673),
.B(n_5660),
.Y(n_5711)
);

AND2x2_ASAP7_75t_L g5712 ( 
.A(n_5674),
.B(n_5668),
.Y(n_5712)
);

AND2x2_ASAP7_75t_L g5713 ( 
.A(n_5680),
.B(n_5668),
.Y(n_5713)
);

INVx2_ASAP7_75t_L g5714 ( 
.A(n_5682),
.Y(n_5714)
);

AOI22xp5_ASAP7_75t_L g5715 ( 
.A1(n_5681),
.A2(n_5519),
.B1(n_5622),
.B2(n_5635),
.Y(n_5715)
);

NOR2xp33_ASAP7_75t_L g5716 ( 
.A(n_5677),
.B(n_5607),
.Y(n_5716)
);

NAND2xp5_ASAP7_75t_L g5717 ( 
.A(n_5676),
.B(n_5654),
.Y(n_5717)
);

NOR3xp33_ASAP7_75t_L g5718 ( 
.A(n_5677),
.B(n_5691),
.C(n_5689),
.Y(n_5718)
);

AND2x2_ASAP7_75t_L g5719 ( 
.A(n_5711),
.B(n_5670),
.Y(n_5719)
);

NAND2x1_ASAP7_75t_L g5720 ( 
.A(n_5713),
.B(n_5604),
.Y(n_5720)
);

OR2x2_ASAP7_75t_L g5721 ( 
.A(n_5709),
.B(n_5691),
.Y(n_5721)
);

O2A1O1Ixp33_ASAP7_75t_L g5722 ( 
.A1(n_5698),
.A2(n_5695),
.B(n_5686),
.C(n_5615),
.Y(n_5722)
);

OR2x2_ASAP7_75t_L g5723 ( 
.A(n_5696),
.B(n_5703),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5714),
.Y(n_5724)
);

NOR2xp33_ASAP7_75t_L g5725 ( 
.A(n_5716),
.B(n_5701),
.Y(n_5725)
);

NAND4xp25_ASAP7_75t_SL g5726 ( 
.A(n_5715),
.B(n_5661),
.C(n_5622),
.D(n_5615),
.Y(n_5726)
);

OR2x2_ASAP7_75t_L g5727 ( 
.A(n_5699),
.B(n_5654),
.Y(n_5727)
);

INVx1_ASAP7_75t_L g5728 ( 
.A(n_5708),
.Y(n_5728)
);

AND2x2_ASAP7_75t_L g5729 ( 
.A(n_5700),
.B(n_5670),
.Y(n_5729)
);

NAND2xp5_ASAP7_75t_L g5730 ( 
.A(n_5712),
.B(n_5685),
.Y(n_5730)
);

INVx1_ASAP7_75t_SL g5731 ( 
.A(n_5699),
.Y(n_5731)
);

OR2x2_ASAP7_75t_L g5732 ( 
.A(n_5710),
.B(n_5655),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_5702),
.Y(n_5733)
);

NOR2xp33_ASAP7_75t_L g5734 ( 
.A(n_5697),
.B(n_5629),
.Y(n_5734)
);

NOR2xp33_ASAP7_75t_L g5735 ( 
.A(n_5707),
.B(n_5706),
.Y(n_5735)
);

BUFx2_ASAP7_75t_L g5736 ( 
.A(n_5729),
.Y(n_5736)
);

AND2x2_ASAP7_75t_L g5737 ( 
.A(n_5719),
.B(n_5718),
.Y(n_5737)
);

AND2x2_ASAP7_75t_L g5738 ( 
.A(n_5731),
.B(n_5704),
.Y(n_5738)
);

AND2x2_ASAP7_75t_L g5739 ( 
.A(n_5735),
.B(n_5591),
.Y(n_5739)
);

INVxp67_ASAP7_75t_SL g5740 ( 
.A(n_5720),
.Y(n_5740)
);

NAND2xp5_ASAP7_75t_L g5741 ( 
.A(n_5734),
.B(n_5685),
.Y(n_5741)
);

AOI221xp5_ASAP7_75t_L g5742 ( 
.A1(n_5726),
.A2(n_5710),
.B1(n_5706),
.B2(n_5646),
.C(n_5643),
.Y(n_5742)
);

INVxp67_ASAP7_75t_L g5743 ( 
.A(n_5725),
.Y(n_5743)
);

INVx1_ASAP7_75t_SL g5744 ( 
.A(n_5721),
.Y(n_5744)
);

AND2x2_ASAP7_75t_L g5745 ( 
.A(n_5730),
.B(n_5591),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5727),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5732),
.Y(n_5747)
);

INVx2_ASAP7_75t_L g5748 ( 
.A(n_5723),
.Y(n_5748)
);

NAND2xp5_ASAP7_75t_L g5749 ( 
.A(n_5740),
.B(n_5705),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_5736),
.Y(n_5750)
);

OR2x2_ASAP7_75t_L g5751 ( 
.A(n_5744),
.B(n_5655),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5738),
.Y(n_5752)
);

AND2x2_ASAP7_75t_L g5753 ( 
.A(n_5737),
.B(n_5733),
.Y(n_5753)
);

OAI22xp5_ASAP7_75t_L g5754 ( 
.A1(n_5744),
.A2(n_5635),
.B1(n_5621),
.B2(n_5604),
.Y(n_5754)
);

NAND2xp5_ASAP7_75t_L g5755 ( 
.A(n_5746),
.B(n_5724),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_5741),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5741),
.Y(n_5757)
);

OAI21xp5_ASAP7_75t_L g5758 ( 
.A1(n_5742),
.A2(n_5722),
.B(n_5717),
.Y(n_5758)
);

INVx2_ASAP7_75t_L g5759 ( 
.A(n_5739),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5745),
.Y(n_5760)
);

INVx2_ASAP7_75t_L g5761 ( 
.A(n_5748),
.Y(n_5761)
);

INVx1_ASAP7_75t_SL g5762 ( 
.A(n_5747),
.Y(n_5762)
);

AND2x2_ASAP7_75t_L g5763 ( 
.A(n_5743),
.B(n_5598),
.Y(n_5763)
);

OAI31xp33_ASAP7_75t_L g5764 ( 
.A1(n_5744),
.A2(n_5695),
.A3(n_5717),
.B(n_5693),
.Y(n_5764)
);

AOI221xp5_ASAP7_75t_L g5765 ( 
.A1(n_5758),
.A2(n_5648),
.B1(n_5651),
.B2(n_5728),
.C(n_5687),
.Y(n_5765)
);

AND2x2_ASAP7_75t_L g5766 ( 
.A(n_5763),
.B(n_5600),
.Y(n_5766)
);

AOI22xp5_ASAP7_75t_L g5767 ( 
.A1(n_5754),
.A2(n_5600),
.B1(n_5612),
.B2(n_5594),
.Y(n_5767)
);

NOR2xp33_ASAP7_75t_L g5768 ( 
.A(n_5762),
.B(n_5629),
.Y(n_5768)
);

INVx1_ASAP7_75t_L g5769 ( 
.A(n_5751),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5749),
.Y(n_5770)
);

INVx1_ASAP7_75t_L g5771 ( 
.A(n_5750),
.Y(n_5771)
);

NAND2xp5_ASAP7_75t_L g5772 ( 
.A(n_5762),
.B(n_5621),
.Y(n_5772)
);

AO22x2_ASAP7_75t_L g5773 ( 
.A1(n_5752),
.A2(n_5669),
.B1(n_5671),
.B2(n_5664),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5753),
.Y(n_5774)
);

AND2x2_ASAP7_75t_L g5775 ( 
.A(n_5759),
.B(n_5761),
.Y(n_5775)
);

OAI21xp33_ASAP7_75t_L g5776 ( 
.A1(n_5755),
.A2(n_5658),
.B(n_5612),
.Y(n_5776)
);

INVx1_ASAP7_75t_L g5777 ( 
.A(n_5772),
.Y(n_5777)
);

A2O1A1Ixp33_ASAP7_75t_L g5778 ( 
.A1(n_5768),
.A2(n_5764),
.B(n_5757),
.C(n_5756),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_5766),
.Y(n_5779)
);

INVx1_ASAP7_75t_L g5780 ( 
.A(n_5773),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_5773),
.Y(n_5781)
);

OAI21xp5_ASAP7_75t_L g5782 ( 
.A1(n_5767),
.A2(n_5760),
.B(n_5764),
.Y(n_5782)
);

INVx1_ASAP7_75t_SL g5783 ( 
.A(n_5775),
.Y(n_5783)
);

NAND2xp5_ASAP7_75t_L g5784 ( 
.A(n_5776),
.B(n_5639),
.Y(n_5784)
);

OAI21xp33_ASAP7_75t_L g5785 ( 
.A1(n_5774),
.A2(n_5771),
.B(n_5770),
.Y(n_5785)
);

OAI221xp5_ASAP7_75t_L g5786 ( 
.A1(n_5765),
.A2(n_5658),
.B1(n_5597),
.B2(n_5613),
.C(n_5639),
.Y(n_5786)
);

AND2x2_ASAP7_75t_L g5787 ( 
.A(n_5769),
.B(n_5594),
.Y(n_5787)
);

OR2x2_ASAP7_75t_L g5788 ( 
.A(n_5783),
.B(n_5617),
.Y(n_5788)
);

NAND2xp5_ASAP7_75t_L g5789 ( 
.A(n_5787),
.B(n_5619),
.Y(n_5789)
);

INVx2_ASAP7_75t_L g5790 ( 
.A(n_5780),
.Y(n_5790)
);

AND2x2_ASAP7_75t_L g5791 ( 
.A(n_5779),
.B(n_5782),
.Y(n_5791)
);

AOI21xp33_ASAP7_75t_L g5792 ( 
.A1(n_5785),
.A2(n_5666),
.B(n_5634),
.Y(n_5792)
);

OAI21xp5_ASAP7_75t_L g5793 ( 
.A1(n_5778),
.A2(n_5666),
.B(n_5634),
.Y(n_5793)
);

XOR2x2_ASAP7_75t_L g5794 ( 
.A(n_5784),
.B(n_5553),
.Y(n_5794)
);

AOI21xp5_ASAP7_75t_L g5795 ( 
.A1(n_5781),
.A2(n_5777),
.B(n_5786),
.Y(n_5795)
);

INVxp67_ASAP7_75t_L g5796 ( 
.A(n_5787),
.Y(n_5796)
);

NAND2xp33_ASAP7_75t_L g5797 ( 
.A(n_5787),
.B(n_5626),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5787),
.Y(n_5798)
);

INVxp67_ASAP7_75t_L g5799 ( 
.A(n_5787),
.Y(n_5799)
);

NAND3xp33_ASAP7_75t_L g5800 ( 
.A(n_5778),
.B(n_5554),
.C(n_5553),
.Y(n_5800)
);

NOR2xp33_ASAP7_75t_L g5801 ( 
.A(n_5783),
.B(n_5625),
.Y(n_5801)
);

CKINVDCx16_ASAP7_75t_R g5802 ( 
.A(n_5782),
.Y(n_5802)
);

AOI22xp5_ASAP7_75t_L g5803 ( 
.A1(n_5783),
.A2(n_5609),
.B1(n_5633),
.B2(n_5632),
.Y(n_5803)
);

NAND3xp33_ASAP7_75t_L g5804 ( 
.A(n_5778),
.B(n_5661),
.C(n_5560),
.Y(n_5804)
);

INVx1_ASAP7_75t_L g5805 ( 
.A(n_5787),
.Y(n_5805)
);

INVx1_ASAP7_75t_SL g5806 ( 
.A(n_5787),
.Y(n_5806)
);

NOR3xp33_ASAP7_75t_L g5807 ( 
.A(n_5802),
.B(n_5552),
.C(n_5614),
.Y(n_5807)
);

NOR4xp25_ASAP7_75t_L g5808 ( 
.A(n_5806),
.B(n_5609),
.C(n_5633),
.D(n_5632),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5803),
.Y(n_5809)
);

AOI211xp5_ASAP7_75t_L g5810 ( 
.A1(n_5792),
.A2(n_5523),
.B(n_5638),
.C(n_5422),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5789),
.Y(n_5811)
);

NOR3xp33_ASAP7_75t_SL g5812 ( 
.A(n_5795),
.B(n_443),
.C(n_444),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_5791),
.Y(n_5813)
);

HB1xp67_ASAP7_75t_L g5814 ( 
.A(n_5793),
.Y(n_5814)
);

AOI21xp33_ASAP7_75t_SL g5815 ( 
.A1(n_5788),
.A2(n_5638),
.B(n_443),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5797),
.Y(n_5816)
);

AOI22xp5_ASAP7_75t_L g5817 ( 
.A1(n_5800),
.A2(n_5566),
.B1(n_5532),
.B2(n_5419),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5794),
.Y(n_5818)
);

OAI22xp5_ASAP7_75t_L g5819 ( 
.A1(n_5804),
.A2(n_5446),
.B1(n_5448),
.B2(n_5404),
.Y(n_5819)
);

NAND2xp5_ASAP7_75t_L g5820 ( 
.A(n_5798),
.B(n_5432),
.Y(n_5820)
);

AO22x2_ASAP7_75t_L g5821 ( 
.A1(n_5805),
.A2(n_5451),
.B1(n_5439),
.B2(n_5432),
.Y(n_5821)
);

NOR2x1_ASAP7_75t_L g5822 ( 
.A(n_5790),
.B(n_5439),
.Y(n_5822)
);

NOR2xp33_ASAP7_75t_L g5823 ( 
.A(n_5796),
.B(n_5490),
.Y(n_5823)
);

NOR2x1_ASAP7_75t_SL g5824 ( 
.A(n_5799),
.B(n_5465),
.Y(n_5824)
);

NOR3xp33_ASAP7_75t_L g5825 ( 
.A(n_5801),
.B(n_5485),
.C(n_5458),
.Y(n_5825)
);

NAND4xp75_ASAP7_75t_L g5826 ( 
.A(n_5795),
.B(n_5502),
.C(n_446),
.D(n_444),
.Y(n_5826)
);

NAND4xp75_ASAP7_75t_L g5827 ( 
.A(n_5795),
.B(n_447),
.C(n_445),
.D(n_446),
.Y(n_5827)
);

AOI21xp5_ASAP7_75t_L g5828 ( 
.A1(n_5789),
.A2(n_5458),
.B(n_5465),
.Y(n_5828)
);

NAND2xp5_ASAP7_75t_L g5829 ( 
.A(n_5803),
.B(n_5469),
.Y(n_5829)
);

NOR3xp33_ASAP7_75t_L g5830 ( 
.A(n_5802),
.B(n_5457),
.C(n_5452),
.Y(n_5830)
);

NOR2xp33_ASAP7_75t_SL g5831 ( 
.A(n_5806),
.B(n_5473),
.Y(n_5831)
);

AOI211xp5_ASAP7_75t_L g5832 ( 
.A1(n_5792),
.A2(n_5457),
.B(n_5452),
.C(n_5471),
.Y(n_5832)
);

OAI221xp5_ASAP7_75t_SL g5833 ( 
.A1(n_5810),
.A2(n_5475),
.B1(n_5471),
.B2(n_5434),
.C(n_5478),
.Y(n_5833)
);

XOR2xp5_ASAP7_75t_L g5834 ( 
.A(n_5827),
.B(n_445),
.Y(n_5834)
);

XNOR2xp5_ASAP7_75t_L g5835 ( 
.A(n_5813),
.B(n_448),
.Y(n_5835)
);

OAI22xp33_ASAP7_75t_L g5836 ( 
.A1(n_5831),
.A2(n_5475),
.B1(n_5417),
.B2(n_5488),
.Y(n_5836)
);

AOI221xp5_ASAP7_75t_L g5837 ( 
.A1(n_5815),
.A2(n_5488),
.B1(n_5486),
.B2(n_5406),
.C(n_453),
.Y(n_5837)
);

AOI21xp5_ASAP7_75t_L g5838 ( 
.A1(n_5814),
.A2(n_448),
.B(n_449),
.Y(n_5838)
);

AOI22xp33_ASAP7_75t_L g5839 ( 
.A1(n_5807),
.A2(n_5825),
.B1(n_5830),
.B2(n_5809),
.Y(n_5839)
);

NAND3xp33_ASAP7_75t_L g5840 ( 
.A(n_5812),
.B(n_452),
.C(n_453),
.Y(n_5840)
);

AOI321xp33_ASAP7_75t_L g5841 ( 
.A1(n_5808),
.A2(n_454),
.A3(n_455),
.B1(n_456),
.B2(n_457),
.C(n_458),
.Y(n_5841)
);

NOR2xp33_ASAP7_75t_L g5842 ( 
.A(n_5820),
.B(n_5823),
.Y(n_5842)
);

O2A1O1Ixp33_ASAP7_75t_SL g5843 ( 
.A1(n_5816),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_5843)
);

XOR2x2_ASAP7_75t_L g5844 ( 
.A(n_5818),
.B(n_459),
.Y(n_5844)
);

AOI22xp5_ASAP7_75t_L g5845 ( 
.A1(n_5811),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.Y(n_5845)
);

XNOR2x1_ASAP7_75t_L g5846 ( 
.A(n_5822),
.B(n_460),
.Y(n_5846)
);

AOI21xp5_ASAP7_75t_L g5847 ( 
.A1(n_5824),
.A2(n_461),
.B(n_462),
.Y(n_5847)
);

AOI21xp5_ASAP7_75t_L g5848 ( 
.A1(n_5829),
.A2(n_463),
.B(n_464),
.Y(n_5848)
);

NOR2xp33_ASAP7_75t_SL g5849 ( 
.A(n_5826),
.B(n_464),
.Y(n_5849)
);

AOI211xp5_ASAP7_75t_L g5850 ( 
.A1(n_5819),
.A2(n_468),
.B(n_466),
.C(n_467),
.Y(n_5850)
);

OR2x2_ASAP7_75t_L g5851 ( 
.A(n_5817),
.B(n_466),
.Y(n_5851)
);

AOI211xp5_ASAP7_75t_SL g5852 ( 
.A1(n_5828),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_5852)
);

AOI22xp33_ASAP7_75t_L g5853 ( 
.A1(n_5821),
.A2(n_473),
.B1(n_470),
.B2(n_471),
.Y(n_5853)
);

INVx1_ASAP7_75t_L g5854 ( 
.A(n_5821),
.Y(n_5854)
);

A2O1A1Ixp33_ASAP7_75t_L g5855 ( 
.A1(n_5832),
.A2(n_471),
.B(n_474),
.C(n_475),
.Y(n_5855)
);

NAND3xp33_ASAP7_75t_L g5856 ( 
.A(n_5812),
.B(n_474),
.C(n_478),
.Y(n_5856)
);

OAI21xp33_ASAP7_75t_L g5857 ( 
.A1(n_5808),
.A2(n_478),
.B(n_479),
.Y(n_5857)
);

NOR3xp33_ASAP7_75t_L g5858 ( 
.A(n_5813),
.B(n_479),
.C(n_480),
.Y(n_5858)
);

XNOR2x1_ASAP7_75t_L g5859 ( 
.A(n_5827),
.B(n_482),
.Y(n_5859)
);

NAND5xp2_ASAP7_75t_L g5860 ( 
.A(n_5839),
.B(n_483),
.C(n_484),
.D(n_486),
.E(n_487),
.Y(n_5860)
);

INVx2_ASAP7_75t_SL g5861 ( 
.A(n_5846),
.Y(n_5861)
);

NOR3xp33_ASAP7_75t_L g5862 ( 
.A(n_5842),
.B(n_483),
.C(n_484),
.Y(n_5862)
);

NOR3x1_ASAP7_75t_L g5863 ( 
.A(n_5840),
.B(n_486),
.C(n_487),
.Y(n_5863)
);

AND5x1_ASAP7_75t_L g5864 ( 
.A(n_5849),
.B(n_488),
.C(n_489),
.D(n_490),
.E(n_492),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5835),
.Y(n_5865)
);

NOR2x1_ASAP7_75t_L g5866 ( 
.A(n_5854),
.B(n_490),
.Y(n_5866)
);

NAND4xp75_ASAP7_75t_L g5867 ( 
.A(n_5848),
.B(n_493),
.C(n_494),
.D(n_495),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5834),
.Y(n_5868)
);

NOR2xp33_ASAP7_75t_SL g5869 ( 
.A(n_5857),
.B(n_493),
.Y(n_5869)
);

INVx1_ASAP7_75t_L g5870 ( 
.A(n_5841),
.Y(n_5870)
);

NOR3xp33_ASAP7_75t_L g5871 ( 
.A(n_5856),
.B(n_496),
.C(n_497),
.Y(n_5871)
);

NOR3xp33_ASAP7_75t_L g5872 ( 
.A(n_5838),
.B(n_496),
.C(n_498),
.Y(n_5872)
);

AND2x4_ASAP7_75t_L g5873 ( 
.A(n_5847),
.B(n_498),
.Y(n_5873)
);

NAND2xp33_ASAP7_75t_SL g5874 ( 
.A(n_5859),
.B(n_499),
.Y(n_5874)
);

NOR3xp33_ASAP7_75t_L g5875 ( 
.A(n_5851),
.B(n_499),
.C(n_500),
.Y(n_5875)
);

NAND3xp33_ASAP7_75t_SL g5876 ( 
.A(n_5852),
.B(n_500),
.C(n_502),
.Y(n_5876)
);

NAND2xp5_ASAP7_75t_L g5877 ( 
.A(n_5858),
.B(n_502),
.Y(n_5877)
);

NOR2x1_ASAP7_75t_L g5878 ( 
.A(n_5855),
.B(n_503),
.Y(n_5878)
);

AND2x2_ASAP7_75t_L g5879 ( 
.A(n_5837),
.B(n_503),
.Y(n_5879)
);

NAND4xp25_ASAP7_75t_L g5880 ( 
.A(n_5850),
.B(n_504),
.C(n_505),
.D(n_506),
.Y(n_5880)
);

INVx3_ASAP7_75t_L g5881 ( 
.A(n_5844),
.Y(n_5881)
);

NOR2x1p5_ASAP7_75t_L g5882 ( 
.A(n_5843),
.B(n_504),
.Y(n_5882)
);

CKINVDCx20_ASAP7_75t_R g5883 ( 
.A(n_5845),
.Y(n_5883)
);

NAND2xp5_ASAP7_75t_L g5884 ( 
.A(n_5873),
.B(n_5853),
.Y(n_5884)
);

NOR2x1_ASAP7_75t_L g5885 ( 
.A(n_5866),
.B(n_5836),
.Y(n_5885)
);

NOR2x1p5_ASAP7_75t_L g5886 ( 
.A(n_5867),
.B(n_5833),
.Y(n_5886)
);

AOI221xp5_ASAP7_75t_L g5887 ( 
.A1(n_5874),
.A2(n_506),
.B1(n_507),
.B2(n_508),
.C(n_509),
.Y(n_5887)
);

O2A1O1Ixp33_ASAP7_75t_L g5888 ( 
.A1(n_5876),
.A2(n_507),
.B(n_508),
.C(n_511),
.Y(n_5888)
);

AO22x2_ASAP7_75t_L g5889 ( 
.A1(n_5861),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_5889)
);

AOI221xp5_ASAP7_75t_L g5890 ( 
.A1(n_5870),
.A2(n_512),
.B1(n_515),
.B2(n_516),
.C(n_517),
.Y(n_5890)
);

OAI21xp5_ASAP7_75t_SL g5891 ( 
.A1(n_5880),
.A2(n_5871),
.B(n_5879),
.Y(n_5891)
);

NOR2xp67_ASAP7_75t_SL g5892 ( 
.A(n_5881),
.B(n_515),
.Y(n_5892)
);

INVx1_ASAP7_75t_L g5893 ( 
.A(n_5882),
.Y(n_5893)
);

XNOR2xp5_ASAP7_75t_L g5894 ( 
.A(n_5865),
.B(n_516),
.Y(n_5894)
);

OAI311xp33_ASAP7_75t_L g5895 ( 
.A1(n_5868),
.A2(n_518),
.A3(n_519),
.B1(n_520),
.C1(n_521),
.Y(n_5895)
);

AO22x2_ASAP7_75t_L g5896 ( 
.A1(n_5873),
.A2(n_518),
.B1(n_519),
.B2(n_520),
.Y(n_5896)
);

NAND4xp25_ASAP7_75t_L g5897 ( 
.A(n_5863),
.B(n_521),
.C(n_522),
.D(n_523),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5877),
.Y(n_5898)
);

NAND3xp33_ASAP7_75t_L g5899 ( 
.A(n_5875),
.B(n_522),
.C(n_524),
.Y(n_5899)
);

OAI22xp5_ASAP7_75t_L g5900 ( 
.A1(n_5883),
.A2(n_524),
.B1(n_525),
.B2(n_526),
.Y(n_5900)
);

NOR4xp25_ASAP7_75t_L g5901 ( 
.A(n_5869),
.B(n_525),
.C(n_527),
.D(n_528),
.Y(n_5901)
);

NOR3xp33_ASAP7_75t_SL g5902 ( 
.A(n_5891),
.B(n_5860),
.C(n_5878),
.Y(n_5902)
);

AND4x1_ASAP7_75t_L g5903 ( 
.A(n_5892),
.B(n_5872),
.C(n_5862),
.D(n_5864),
.Y(n_5903)
);

NAND2xp5_ASAP7_75t_SL g5904 ( 
.A(n_5901),
.B(n_528),
.Y(n_5904)
);

NOR3xp33_ASAP7_75t_L g5905 ( 
.A(n_5893),
.B(n_530),
.C(n_531),
.Y(n_5905)
);

OAI22xp5_ASAP7_75t_L g5906 ( 
.A1(n_5899),
.A2(n_531),
.B1(n_532),
.B2(n_534),
.Y(n_5906)
);

INVx2_ASAP7_75t_L g5907 ( 
.A(n_5889),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_5896),
.Y(n_5908)
);

NOR2xp33_ASAP7_75t_L g5909 ( 
.A(n_5897),
.B(n_532),
.Y(n_5909)
);

NOR3xp33_ASAP7_75t_L g5910 ( 
.A(n_5884),
.B(n_534),
.C(n_535),
.Y(n_5910)
);

NAND3xp33_ASAP7_75t_L g5911 ( 
.A(n_5887),
.B(n_536),
.C(n_537),
.Y(n_5911)
);

OAI22xp5_ASAP7_75t_L g5912 ( 
.A1(n_5885),
.A2(n_536),
.B1(n_538),
.B2(n_539),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5894),
.Y(n_5913)
);

NAND2xp5_ASAP7_75t_SL g5914 ( 
.A(n_5888),
.B(n_539),
.Y(n_5914)
);

NOR2xp33_ASAP7_75t_L g5915 ( 
.A(n_5898),
.B(n_5900),
.Y(n_5915)
);

XNOR2x1_ASAP7_75t_L g5916 ( 
.A(n_5886),
.B(n_540),
.Y(n_5916)
);

NAND5xp2_ASAP7_75t_L g5917 ( 
.A(n_5890),
.B(n_540),
.C(n_541),
.D(n_542),
.E(n_543),
.Y(n_5917)
);

AOI21xp33_ASAP7_75t_L g5918 ( 
.A1(n_5916),
.A2(n_5889),
.B(n_5895),
.Y(n_5918)
);

NAND2xp5_ASAP7_75t_L g5919 ( 
.A(n_5905),
.B(n_5910),
.Y(n_5919)
);

OR3x1_ASAP7_75t_L g5920 ( 
.A(n_5917),
.B(n_5909),
.C(n_5908),
.Y(n_5920)
);

NOR3xp33_ASAP7_75t_L g5921 ( 
.A(n_5915),
.B(n_5913),
.C(n_5914),
.Y(n_5921)
);

NAND2x1_ASAP7_75t_L g5922 ( 
.A(n_5907),
.B(n_541),
.Y(n_5922)
);

A2O1A1Ixp33_ASAP7_75t_L g5923 ( 
.A1(n_5911),
.A2(n_542),
.B(n_544),
.C(n_545),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5904),
.Y(n_5924)
);

NAND4xp25_ASAP7_75t_L g5925 ( 
.A(n_5906),
.B(n_5912),
.C(n_5903),
.D(n_5902),
.Y(n_5925)
);

OAI21xp5_ASAP7_75t_L g5926 ( 
.A1(n_5909),
.A2(n_544),
.B(n_545),
.Y(n_5926)
);

AOI22xp5_ASAP7_75t_L g5927 ( 
.A1(n_5909),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.Y(n_5927)
);

NOR3xp33_ASAP7_75t_L g5928 ( 
.A(n_5915),
.B(n_551),
.C(n_552),
.Y(n_5928)
);

AOI22xp33_ASAP7_75t_L g5929 ( 
.A1(n_5909),
.A2(n_552),
.B1(n_554),
.B2(n_556),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5916),
.Y(n_5930)
);

NAND3xp33_ASAP7_75t_SL g5931 ( 
.A(n_5908),
.B(n_556),
.C(n_557),
.Y(n_5931)
);

NAND3xp33_ASAP7_75t_SL g5932 ( 
.A(n_5908),
.B(n_557),
.C(n_558),
.Y(n_5932)
);

AO22x2_ASAP7_75t_L g5933 ( 
.A1(n_5916),
.A2(n_558),
.B1(n_559),
.B2(n_561),
.Y(n_5933)
);

NOR3xp33_ASAP7_75t_L g5934 ( 
.A(n_5915),
.B(n_561),
.C(n_562),
.Y(n_5934)
);

OAI22xp5_ASAP7_75t_SL g5935 ( 
.A1(n_5922),
.A2(n_563),
.B1(n_564),
.B2(n_566),
.Y(n_5935)
);

NAND2xp5_ASAP7_75t_L g5936 ( 
.A(n_5928),
.B(n_563),
.Y(n_5936)
);

OAI21x1_ASAP7_75t_L g5937 ( 
.A1(n_5926),
.A2(n_566),
.B(n_568),
.Y(n_5937)
);

INVx1_ASAP7_75t_L g5938 ( 
.A(n_5933),
.Y(n_5938)
);

INVx2_ASAP7_75t_L g5939 ( 
.A(n_5933),
.Y(n_5939)
);

AND2x2_ASAP7_75t_SL g5940 ( 
.A(n_5921),
.B(n_570),
.Y(n_5940)
);

AND2x4_ASAP7_75t_L g5941 ( 
.A(n_5924),
.B(n_570),
.Y(n_5941)
);

OAI22xp5_ASAP7_75t_SL g5942 ( 
.A1(n_5920),
.A2(n_572),
.B1(n_573),
.B2(n_574),
.Y(n_5942)
);

NAND2xp5_ASAP7_75t_L g5943 ( 
.A(n_5934),
.B(n_573),
.Y(n_5943)
);

HB1xp67_ASAP7_75t_L g5944 ( 
.A(n_5931),
.Y(n_5944)
);

INVx1_ASAP7_75t_L g5945 ( 
.A(n_5932),
.Y(n_5945)
);

AOI221xp5_ASAP7_75t_L g5946 ( 
.A1(n_5918),
.A2(n_574),
.B1(n_575),
.B2(n_576),
.C(n_577),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_5923),
.Y(n_5947)
);

NAND2x1_ASAP7_75t_L g5948 ( 
.A(n_5938),
.B(n_5927),
.Y(n_5948)
);

OR4x2_ASAP7_75t_L g5949 ( 
.A(n_5940),
.B(n_5925),
.C(n_5919),
.D(n_5930),
.Y(n_5949)
);

XNOR2xp5_ASAP7_75t_L g5950 ( 
.A(n_5942),
.B(n_5929),
.Y(n_5950)
);

O2A1O1Ixp33_ASAP7_75t_L g5951 ( 
.A1(n_5939),
.A2(n_579),
.B(n_580),
.C(n_581),
.Y(n_5951)
);

OAI22x1_ASAP7_75t_L g5952 ( 
.A1(n_5945),
.A2(n_580),
.B1(n_582),
.B2(n_583),
.Y(n_5952)
);

INVx1_ASAP7_75t_L g5953 ( 
.A(n_5937),
.Y(n_5953)
);

XOR2xp5_ASAP7_75t_L g5954 ( 
.A(n_5944),
.B(n_584),
.Y(n_5954)
);

OAI22xp5_ASAP7_75t_SL g5955 ( 
.A1(n_5949),
.A2(n_5935),
.B1(n_5947),
.B2(n_5943),
.Y(n_5955)
);

AOI21xp5_ASAP7_75t_L g5956 ( 
.A1(n_5948),
.A2(n_5936),
.B(n_5946),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5954),
.Y(n_5957)
);

XNOR2x1_ASAP7_75t_L g5958 ( 
.A(n_5950),
.B(n_5941),
.Y(n_5958)
);

INVx1_ASAP7_75t_L g5959 ( 
.A(n_5953),
.Y(n_5959)
);

AND4x1_ASAP7_75t_L g5960 ( 
.A(n_5951),
.B(n_584),
.C(n_586),
.D(n_588),
.Y(n_5960)
);

NAND2xp5_ASAP7_75t_L g5961 ( 
.A(n_5952),
.B(n_586),
.Y(n_5961)
);

AND2x4_ASAP7_75t_L g5962 ( 
.A(n_5957),
.B(n_588),
.Y(n_5962)
);

HB1xp67_ASAP7_75t_L g5963 ( 
.A(n_5960),
.Y(n_5963)
);

AND2x2_ASAP7_75t_SL g5964 ( 
.A(n_5961),
.B(n_589),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5955),
.Y(n_5965)
);

AOI21xp5_ASAP7_75t_L g5966 ( 
.A1(n_5956),
.A2(n_590),
.B(n_591),
.Y(n_5966)
);

INVx3_ASAP7_75t_L g5967 ( 
.A(n_5958),
.Y(n_5967)
);

CKINVDCx20_ASAP7_75t_R g5968 ( 
.A(n_5967),
.Y(n_5968)
);

AOI22x1_ASAP7_75t_L g5969 ( 
.A1(n_5965),
.A2(n_5959),
.B1(n_593),
.B2(n_594),
.Y(n_5969)
);

CKINVDCx20_ASAP7_75t_R g5970 ( 
.A(n_5963),
.Y(n_5970)
);

CKINVDCx20_ASAP7_75t_R g5971 ( 
.A(n_5966),
.Y(n_5971)
);

AO22x2_ASAP7_75t_L g5972 ( 
.A1(n_5964),
.A2(n_592),
.B1(n_595),
.B2(n_596),
.Y(n_5972)
);

OAI22x1_ASAP7_75t_L g5973 ( 
.A1(n_5969),
.A2(n_5962),
.B1(n_5968),
.B2(n_5970),
.Y(n_5973)
);

NAND2xp5_ASAP7_75t_L g5974 ( 
.A(n_5972),
.B(n_597),
.Y(n_5974)
);

INVx1_ASAP7_75t_L g5975 ( 
.A(n_5971),
.Y(n_5975)
);

XOR2xp5_ASAP7_75t_L g5976 ( 
.A(n_5968),
.B(n_597),
.Y(n_5976)
);

OAI21xp5_ASAP7_75t_L g5977 ( 
.A1(n_5974),
.A2(n_598),
.B(n_599),
.Y(n_5977)
);

NOR4xp75_ASAP7_75t_L g5978 ( 
.A(n_5973),
.B(n_600),
.C(n_602),
.D(n_603),
.Y(n_5978)
);

INVx2_ASAP7_75t_L g5979 ( 
.A(n_5976),
.Y(n_5979)
);

AO21x2_ASAP7_75t_L g5980 ( 
.A1(n_5975),
.A2(n_603),
.B(n_604),
.Y(n_5980)
);

AO21x1_ASAP7_75t_L g5981 ( 
.A1(n_5975),
.A2(n_605),
.B(n_606),
.Y(n_5981)
);

AOI222xp33_ASAP7_75t_L g5982 ( 
.A1(n_5979),
.A2(n_606),
.B1(n_607),
.B2(n_608),
.C1(n_611),
.C2(n_612),
.Y(n_5982)
);

OR2x2_ASAP7_75t_L g5983 ( 
.A(n_5977),
.B(n_607),
.Y(n_5983)
);

OAI22xp5_ASAP7_75t_L g5984 ( 
.A1(n_5978),
.A2(n_608),
.B1(n_613),
.B2(n_615),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5980),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5981),
.Y(n_5986)
);

INVxp67_ASAP7_75t_L g5987 ( 
.A(n_5979),
.Y(n_5987)
);

HB1xp67_ASAP7_75t_L g5988 ( 
.A(n_5978),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5980),
.Y(n_5989)
);

AO21x2_ASAP7_75t_L g5990 ( 
.A1(n_5985),
.A2(n_617),
.B(n_619),
.Y(n_5990)
);

OAI21xp5_ASAP7_75t_L g5991 ( 
.A1(n_5987),
.A2(n_619),
.B(n_621),
.Y(n_5991)
);

OA21x2_ASAP7_75t_L g5992 ( 
.A1(n_5989),
.A2(n_621),
.B(n_622),
.Y(n_5992)
);

OAI22xp5_ASAP7_75t_L g5993 ( 
.A1(n_5983),
.A2(n_623),
.B1(n_624),
.B2(n_625),
.Y(n_5993)
);

OAI21xp5_ASAP7_75t_SL g5994 ( 
.A1(n_5988),
.A2(n_623),
.B(n_624),
.Y(n_5994)
);

NAND2xp5_ASAP7_75t_L g5995 ( 
.A(n_5984),
.B(n_626),
.Y(n_5995)
);

AOI21xp5_ASAP7_75t_L g5996 ( 
.A1(n_5986),
.A2(n_627),
.B(n_628),
.Y(n_5996)
);

AOI21xp33_ASAP7_75t_L g5997 ( 
.A1(n_5982),
.A2(n_629),
.B(n_630),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5995),
.Y(n_5998)
);

AO21x2_ASAP7_75t_L g5999 ( 
.A1(n_5997),
.A2(n_631),
.B(n_663),
.Y(n_5999)
);

OAI22xp33_ASAP7_75t_L g6000 ( 
.A1(n_5994),
.A2(n_668),
.B1(n_670),
.B2(n_671),
.Y(n_6000)
);

OAI22xp33_ASAP7_75t_L g6001 ( 
.A1(n_5993),
.A2(n_672),
.B1(n_674),
.B2(n_678),
.Y(n_6001)
);

OAI211xp5_ASAP7_75t_SL g6002 ( 
.A1(n_5996),
.A2(n_679),
.B(n_680),
.C(n_682),
.Y(n_6002)
);

BUFx3_ASAP7_75t_L g6003 ( 
.A(n_5992),
.Y(n_6003)
);

OR2x6_ASAP7_75t_L g6004 ( 
.A(n_6003),
.B(n_5991),
.Y(n_6004)
);

OR2x6_ASAP7_75t_L g6005 ( 
.A(n_5998),
.B(n_5990),
.Y(n_6005)
);

AOI21xp5_ASAP7_75t_L g6006 ( 
.A1(n_6004),
.A2(n_5999),
.B(n_6001),
.Y(n_6006)
);

AOI211xp5_ASAP7_75t_L g6007 ( 
.A1(n_6006),
.A2(n_6002),
.B(n_6000),
.C(n_6005),
.Y(n_6007)
);


endmodule