module real_jpeg_7826_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_1),
.A2(n_53),
.B1(n_61),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_1),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_121),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_1),
.A2(n_38),
.B1(n_41),
.B2(n_121),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_121),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_40),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_4),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_4),
.A2(n_55),
.B(n_59),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_4),
.A2(n_53),
.B1(n_61),
.B2(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_4),
.B(n_65),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_38),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_4),
.B(n_38),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_4),
.A2(n_82),
.B1(n_83),
.B2(n_201),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_53),
.B1(n_61),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_5),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_102),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_102),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_5),
.A2(n_38),
.B1(n_41),
.B2(n_102),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_SL g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_38),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_48),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_12),
.A2(n_29),
.B1(n_58),
.B2(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_12),
.A2(n_29),
.B1(n_38),
.B2(n_41),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_13),
.A2(n_35),
.B1(n_53),
.B2(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_13),
.A2(n_35),
.B1(n_58),
.B2(n_59),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_13),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_15),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_15),
.A2(n_27),
.B1(n_30),
.B2(n_62),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_15),
.A2(n_38),
.B1(n_41),
.B2(n_62),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_106),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_90),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_78),
.B2(n_79),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_24),
.B(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_25),
.A2(n_83),
.B(n_128),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_32),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_30),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_27),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_30),
.B(n_46),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_30),
.B(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_31),
.A2(n_32),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_32),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_33),
.A2(n_82),
.B(n_185),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_34),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_37),
.A2(n_45),
.B(n_96),
.Y(n_95)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_43),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_41),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_38),
.B(n_69),
.Y(n_229)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_41),
.A2(n_74),
.B1(n_224),
.B2(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_47),
.B(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_42),
.A2(n_45),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_42),
.A2(n_45),
.B1(n_191),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_42),
.A2(n_45),
.B1(n_214),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_42),
.A2(n_222),
.B(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_44),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_45),
.B(n_125),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_45),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_66),
.B2(n_77),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_60),
.B(n_63),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_57),
.B1(n_60),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_52),
.A2(n_57),
.B1(n_101),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_52),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B(n_56),
.C(n_57),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_53),
.A2(n_54),
.B(n_125),
.C(n_126),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_55),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_68),
.B(n_69),
.C(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_69),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g224 ( 
.A(n_59),
.B(n_125),
.CON(n_224),
.SN(n_224)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_65),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B(n_72),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_76),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_67),
.A2(n_115),
.B1(n_116),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_67),
.A2(n_115),
.B1(n_145),
.B2(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_67),
.B(n_125),
.Y(n_212)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_104),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_68),
.A2(n_73),
.B1(n_169),
.B2(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_73),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_73),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_89),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_82),
.A2(n_83),
.B1(n_93),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_82),
.A2(n_83),
.B1(n_183),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_82),
.A2(n_84),
.B(n_94),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_83),
.B(n_125),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_87),
.A2(n_98),
.B(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.C(n_103),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_92),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_111),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_110),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_112),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_122),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B(n_117),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_174),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_155),
.B(n_173),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_175),
.C(n_256),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_152),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_152),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.C(n_141),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_150),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_144),
.B1(n_150),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_151),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_156),
.B(n_158),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_159),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_162),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.C(n_171),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_166),
.A2(n_167),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_170),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_250),
.B(n_255),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_233),
.B(n_249),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_217),
.B(n_232),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_208),
.B(n_216),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_197),
.B(n_207),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_186),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_196),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_196),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_190),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_202),
.B(n_206),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_199),
.B(n_200),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_210),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_211),
.B(n_218),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.CI(n_215),
.CON(n_211),
.SN(n_211)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_227),
.B2(n_231),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_221),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_223),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_226),
.C(n_231),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_227),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_230),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_234),
.B(n_235),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_241),
.B2(n_242),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_244),
.C(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_243),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);


endmodule