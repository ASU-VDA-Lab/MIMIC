module real_jpeg_5156_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_2),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_2),
.Y(n_134)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_5),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_5),
.A2(n_33),
.B1(n_188),
.B2(n_191),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_64),
.B1(n_94),
.B2(n_97),
.Y(n_93)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_7),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_8),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_8),
.B(n_122),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_8),
.A2(n_119),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_8),
.B(n_165),
.C(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_8),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_8),
.B(n_92),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_9),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_10),
.A2(n_40),
.B1(n_80),
.B2(n_83),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_10),
.A2(n_40),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_150),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_148),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_86),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_86),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_52),
.C(n_60),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_15),
.A2(n_16),
.B1(n_52),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_28),
.B(n_36),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_20),
.B1(n_24),
.B2(n_26),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_21),
.Y(n_135)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_25),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_28),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_89)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_44)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_31),
.Y(n_156)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_32),
.Y(n_146)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_32),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_37),
.B(n_92),
.Y(n_159)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_39),
.A2(n_121),
.A3(n_139),
.B1(n_142),
.B2(n_144),
.Y(n_138)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_42),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_52),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_60),
.B(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_69),
.B(n_76),
.Y(n_60)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_61),
.Y(n_200)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_69),
.A2(n_76),
.B(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_79),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_70),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_75),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_129),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_98),
.B2(n_99),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_90),
.A2(n_154),
.B(n_159),
.Y(n_153)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_114),
.B(n_123),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_105),
.Y(n_110)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_119),
.B(n_120),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_138),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_136),
.B(n_137),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_187),
.B(n_193),
.Y(n_186)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_171),
.B(n_205),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_168),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_168),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_160),
.B1(n_161),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_197),
.B(n_204),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_185),
.B(n_196),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_184),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_181),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_195),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_195),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_202),
.Y(n_204)
);


endmodule