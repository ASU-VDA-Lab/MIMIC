module fake_jpeg_1141_n_12 (n_3, n_2, n_1, n_0, n_4, n_12);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_12;

wire n_11;
wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx1_ASAP7_75t_L g5 ( 
.A(n_2),
.Y(n_5)
);

AOI22xp5_ASAP7_75t_L g6 ( 
.A1(n_1),
.A2(n_3),
.B1(n_0),
.B2(n_4),
.Y(n_6)
);

CKINVDCx16_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_7),
.Y(n_9)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

AOI322xp5_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_6),
.A3(n_8),
.B1(n_10),
.B2(n_5),
.C1(n_9),
.C2(n_0),
.Y(n_12)
);


endmodule