module fake_netlist_5_835_n_1717 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1717);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1717;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_SL g158 ( 
.A(n_150),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_28),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_42),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_129),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_93),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_43),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_61),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_64),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_98),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_101),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_34),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_55),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_123),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_20),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_8),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_69),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_108),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_119),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_131),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_15),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_79),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_88),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_9),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_34),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_74),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_51),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_40),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_112),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_16),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_103),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_122),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_11),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_32),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_16),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_0),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_156),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_6),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_54),
.Y(n_211)
);

HB1xp67_ASAP7_75t_SL g212 ( 
.A(n_49),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_102),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_8),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_146),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_11),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_151),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_121),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_115),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_75),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_136),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_113),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_86),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_22),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_152),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_107),
.Y(n_228)
);

INVxp33_ASAP7_75t_R g229 ( 
.A(n_27),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_33),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_58),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_59),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_46),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_138),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_25),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_39),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_41),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_111),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_117),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_80),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_97),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_82),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_70),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_27),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_84),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_85),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_31),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_23),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_65),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_44),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_96),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_52),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_35),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_7),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_25),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_47),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_130),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_77),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_45),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_144),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_143),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_100),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_155),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_21),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_21),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_153),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_44),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_140),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_30),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_147),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_31),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_81),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_116),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_29),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_60),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_53),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_1),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_124),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_30),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_50),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_142),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_48),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_106),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_141),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_66),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_18),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_118),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_35),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_1),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_83),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_15),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_2),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_41),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_76),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_104),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_48),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_26),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_148),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_22),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_6),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_109),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_110),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_42),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_134),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_26),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_46),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_90),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_5),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_43),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_259),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_230),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_230),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_263),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_192),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_206),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_230),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_230),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_223),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_181),
.B(n_0),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_245),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_230),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_166),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_186),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_230),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_188),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_190),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_191),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_2),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_313),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_307),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_161),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_243),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_197),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_200),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_249),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_193),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_295),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_204),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_184),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_194),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_257),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_208),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_160),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_160),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_181),
.B(n_3),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_212),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_210),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_163),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_215),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_205),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_238),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_187),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_217),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_163),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_294),
.B(n_3),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_241),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_226),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_189),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_241),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_262),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_262),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_201),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_202),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_168),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_170),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_198),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_209),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_185),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_213),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_233),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_214),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_195),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_R g387 ( 
.A(n_216),
.B(n_89),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_169),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_235),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_169),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_321),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_328),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_315),
.B(n_306),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_306),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_322),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_322),
.B(n_205),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_350),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_325),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_329),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_329),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_329),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_316),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_183),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_366),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_372),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_339),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_327),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_376),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_341),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_183),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_316),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_331),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_199),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_R g425 ( 
.A(n_377),
.B(n_218),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_317),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_373),
.B(n_199),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g429 ( 
.A(n_318),
.B(n_282),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_315),
.B(n_234),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_320),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_340),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_362),
.B(n_270),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_270),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_323),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_381),
.Y(n_436)
);

NAND2x1_ASAP7_75t_L g437 ( 
.A(n_326),
.B(n_166),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_383),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_319),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_385),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_343),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_330),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_324),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_330),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_388),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_332),
.Y(n_446)
);

OA21x2_ASAP7_75t_L g447 ( 
.A1(n_379),
.A2(n_203),
.B(n_196),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_388),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_390),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_365),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_342),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_347),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_351),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_386),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_332),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_352),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_333),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_333),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_346),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_397),
.B(n_319),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_422),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_449),
.Y(n_466)
);

INVx6_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_422),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_412),
.B(n_166),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_412),
.B(n_166),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_423),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_412),
.B(n_359),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_456),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_428),
.B(n_166),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_427),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_436),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_421),
.A2(n_338),
.B1(n_369),
.B2(n_304),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_437),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_435),
.B(n_334),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_400),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_435),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_456),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_400),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_453),
.Y(n_492)
);

OAI22xp33_ASAP7_75t_L g493 ( 
.A1(n_404),
.A2(n_250),
.B1(n_284),
.B2(n_260),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_413),
.B(n_334),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_451),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_428),
.B(n_368),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_456),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_428),
.B(n_303),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_428),
.B(n_303),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_449),
.B(n_370),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_429),
.B(n_303),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_402),
.B(n_344),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_437),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_L g505 ( 
.A(n_414),
.B(n_303),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_399),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_454),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_429),
.B(n_303),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_425),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_430),
.B(n_344),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_404),
.B(n_345),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_442),
.B(n_345),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_456),
.B(n_349),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_444),
.B(n_349),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_454),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_SL g518 ( 
.A(n_439),
.B(n_251),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_396),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_456),
.Y(n_520)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_447),
.B(n_296),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_411),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_SL g523 ( 
.A1(n_424),
.A2(n_375),
.B(n_304),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_455),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_411),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_406),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

OAI21xp33_ASAP7_75t_L g529 ( 
.A1(n_462),
.A2(n_361),
.B(n_353),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_413),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_413),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_426),
.B(n_353),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_426),
.B(n_361),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_456),
.B(n_363),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_398),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_411),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_398),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_431),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_426),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_426),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_431),
.B(n_363),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_431),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_440),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_439),
.B(n_364),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_443),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_446),
.B(n_367),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_411),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_401),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_458),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_SL g553 ( 
.A(n_457),
.B(n_271),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_393),
.B(n_395),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_459),
.B(n_367),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_458),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_460),
.B(n_371),
.Y(n_557)
);

CKINVDCx11_ASAP7_75t_R g558 ( 
.A(n_391),
.Y(n_558)
);

NOR2x1p5_ASAP7_75t_L g559 ( 
.A(n_415),
.B(n_371),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_433),
.B(n_384),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_393),
.B(n_384),
.Y(n_561)
);

OAI21xp33_ASAP7_75t_SL g562 ( 
.A1(n_395),
.A2(n_296),
.B(n_211),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_458),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_434),
.A2(n_255),
.B1(n_277),
.B2(n_247),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_411),
.Y(n_566)
);

BUFx8_ASAP7_75t_SL g567 ( 
.A(n_407),
.Y(n_567)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_441),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_434),
.B(n_355),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_434),
.B(n_207),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_418),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_458),
.B(n_389),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_403),
.B(n_389),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_405),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_452),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_434),
.B(n_222),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_447),
.A2(n_356),
.B1(n_231),
.B2(n_228),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_403),
.B(n_158),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_447),
.A2(n_232),
.B1(n_289),
.B2(n_300),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_447),
.A2(n_348),
.B1(n_246),
.B2(n_314),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_417),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_452),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_417),
.B(n_176),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_L g584 ( 
.A(n_416),
.B(n_285),
.C(n_236),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_452),
.B(n_290),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_445),
.B(n_205),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_445),
.A2(n_234),
.B1(n_266),
.B2(n_272),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_405),
.Y(n_588)
);

INVxp33_ASAP7_75t_L g589 ( 
.A(n_448),
.Y(n_589)
);

AND2x4_ASAP7_75t_SL g590 ( 
.A(n_432),
.B(n_234),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_405),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_420),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_452),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_420),
.B(n_311),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_408),
.B(n_219),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_452),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_448),
.B(n_162),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_408),
.B(n_220),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_452),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_448),
.B(n_450),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_408),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_409),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_450),
.B(n_221),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_461),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_450),
.B(n_162),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_409),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_409),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_410),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_419),
.B(n_311),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_438),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_410),
.A2(n_237),
.B1(n_312),
.B2(n_182),
.Y(n_611)
);

BUFx10_ASAP7_75t_L g612 ( 
.A(n_410),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_428),
.B(n_266),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_507),
.B(n_224),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_495),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_507),
.B(n_521),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_521),
.B(n_225),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_560),
.A2(n_227),
.B1(n_239),
.B2(n_240),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_490),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_502),
.B(n_164),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_589),
.B(n_242),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_465),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_589),
.B(n_244),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_508),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_463),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_465),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_464),
.B(n_248),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_468),
.B(n_253),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_586),
.B(n_311),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_470),
.B(n_261),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_472),
.B(n_475),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_500),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_517),
.Y(n_634)
);

INVxp33_ASAP7_75t_L g635 ( 
.A(n_567),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_480),
.B(n_264),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_483),
.A2(n_265),
.B(n_267),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_488),
.B(n_274),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_524),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_573),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_572),
.B(n_473),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_551),
.B(n_291),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_565),
.A2(n_577),
.B1(n_579),
.B2(n_483),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_545),
.B(n_159),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_525),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_467),
.B(n_276),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_485),
.B(n_159),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_565),
.A2(n_504),
.B1(n_570),
.B2(n_613),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_487),
.B(n_164),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_528),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_467),
.B(n_279),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_504),
.B(n_287),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_467),
.B(n_288),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_474),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_494),
.B(n_532),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_533),
.B(n_165),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_529),
.B(n_165),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_581),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_610),
.B(n_229),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_541),
.B(n_167),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_600),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_474),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_482),
.B(n_269),
.C(n_252),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_512),
.A2(n_167),
.B(n_312),
.C(n_174),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_503),
.B(n_171),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_503),
.B(n_496),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_551),
.B(n_254),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_561),
.B(n_580),
.C(n_587),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_SL g669 ( 
.A1(n_568),
.A2(n_310),
.B1(n_308),
.B2(n_305),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_594),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_612),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_515),
.A2(n_171),
.B1(n_172),
.B2(n_309),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_611),
.B(n_273),
.C(n_256),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_496),
.B(n_172),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_592),
.Y(n_675)
);

NAND3xp33_ASAP7_75t_L g676 ( 
.A(n_584),
.B(n_275),
.C(n_258),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_565),
.A2(n_293),
.B1(n_310),
.B2(n_175),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_500),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_609),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_518),
.Y(n_680)
);

NAND2x1_ASAP7_75t_L g681 ( 
.A(n_600),
.B(n_56),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_500),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_549),
.B(n_268),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_496),
.B(n_173),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_487),
.B(n_173),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_466),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_513),
.B(n_280),
.C(n_278),
.Y(n_687)
);

AND2x6_ASAP7_75t_SL g688 ( 
.A(n_514),
.B(n_179),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_530),
.B(n_174),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_531),
.B(n_182),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_487),
.B(n_237),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_600),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_539),
.B(n_292),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_516),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_604),
.B(n_559),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_555),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_540),
.B(n_292),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_597),
.B(n_309),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_605),
.B(n_177),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_608),
.B(n_466),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_600),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_569),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_558),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_608),
.B(n_299),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_484),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_477),
.B(n_299),
.Y(n_706)
);

AND2x6_ASAP7_75t_SL g707 ( 
.A(n_557),
.B(n_308),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_612),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_553),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_570),
.A2(n_175),
.B1(n_305),
.B2(n_302),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_515),
.B(n_177),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_570),
.A2(n_178),
.B1(n_302),
.B2(n_298),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_477),
.A2(n_180),
.B1(n_283),
.B2(n_281),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_571),
.B(n_298),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_554),
.B(n_606),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_613),
.B(n_387),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_534),
.A2(n_180),
.B1(n_272),
.B2(n_266),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_534),
.A2(n_513),
.B1(n_613),
.B2(n_569),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_527),
.Y(n_719)
);

AO221x1_ASAP7_75t_L g720 ( 
.A1(n_493),
.A2(n_272),
.B1(n_293),
.B2(n_179),
.C(n_178),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_606),
.B(n_132),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_569),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_606),
.B(n_126),
.Y(n_723)
);

NAND2x1p5_ASAP7_75t_L g724 ( 
.A(n_499),
.B(n_120),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_595),
.B(n_99),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_598),
.B(n_95),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_578),
.B(n_94),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_603),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_613),
.A2(n_87),
.B1(n_73),
.B2(n_67),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_575),
.B(n_62),
.Y(n_730)
);

INVx8_ASAP7_75t_L g731 ( 
.A(n_613),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_603),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_575),
.B(n_57),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_518),
.B(n_4),
.Y(n_734)
);

BUFx12f_ASAP7_75t_L g735 ( 
.A(n_558),
.Y(n_735)
);

NOR2x1p5_ASAP7_75t_L g736 ( 
.A(n_527),
.B(n_4),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_570),
.A2(n_478),
.B1(n_498),
.B2(n_505),
.Y(n_737)
);

NAND2x1_ASAP7_75t_L g738 ( 
.A(n_536),
.B(n_5),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_583),
.B(n_53),
.Y(n_739)
);

BUFx5_ASAP7_75t_L g740 ( 
.A(n_570),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_576),
.B(n_7),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_582),
.B(n_10),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_582),
.B(n_10),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_484),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_486),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_553),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_510),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_593),
.B(n_12),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_510),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_590),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_SL g751 ( 
.A(n_469),
.B(n_12),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_511),
.B(n_52),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_568),
.B(n_13),
.C(n_14),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_590),
.B(n_13),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_481),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_486),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_570),
.A2(n_14),
.B1(n_17),
.B2(n_18),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_566),
.B(n_19),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_519),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_491),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_593),
.B(n_19),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_576),
.B(n_20),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_519),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_535),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_546),
.B(n_23),
.Y(n_765)
);

AND2x6_ASAP7_75t_SL g766 ( 
.A(n_544),
.B(n_24),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_538),
.B(n_28),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_523),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_538),
.B(n_36),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_505),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_535),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_542),
.B(n_547),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_543),
.B(n_37),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_543),
.B(n_50),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_562),
.B(n_38),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_547),
.B(n_49),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_501),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_491),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_588),
.B(n_591),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_499),
.A2(n_509),
.B1(n_501),
.B2(n_471),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_588),
.B(n_39),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_596),
.B(n_40),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_469),
.B(n_471),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_719),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_641),
.B(n_506),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_655),
.B(n_506),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_661),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_715),
.A2(n_520),
.B(n_497),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_640),
.B(n_591),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_783),
.A2(n_616),
.B(n_617),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_660),
.B(n_591),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_667),
.B(n_537),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_757),
.A2(n_509),
.B1(n_498),
.B2(n_478),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_779),
.A2(n_520),
.B(n_497),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_616),
.A2(n_552),
.B1(n_564),
.B2(n_556),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_772),
.A2(n_666),
.B(n_627),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_660),
.B(n_588),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_741),
.A2(n_537),
.B(n_602),
.C(n_607),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_711),
.B(n_585),
.C(n_548),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_714),
.B(n_585),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_728),
.B(n_591),
.Y(n_801)
);

AOI33xp33_ASAP7_75t_L g802 ( 
.A1(n_677),
.A2(n_45),
.A3(n_47),
.B1(n_607),
.B2(n_563),
.B3(n_599),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_741),
.A2(n_596),
.B(n_574),
.C(n_601),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_771),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_783),
.A2(n_476),
.B(n_497),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_661),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_633),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_742),
.A2(n_601),
.B(n_574),
.C(n_478),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_732),
.B(n_588),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_SL g810 ( 
.A(n_680),
.B(n_526),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_747),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_749),
.Y(n_812)
);

AOI21x1_ASAP7_75t_L g813 ( 
.A1(n_617),
.A2(n_612),
.B(n_476),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_759),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_630),
.B(n_683),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_731),
.A2(n_489),
.B(n_550),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_694),
.B(n_489),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_735),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_718),
.A2(n_601),
.B1(n_574),
.B2(n_550),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_646),
.A2(n_536),
.B(n_479),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_651),
.A2(n_479),
.B(n_522),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_757),
.A2(n_478),
.B1(n_498),
.B2(n_479),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_661),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_633),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_711),
.B(n_479),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_661),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_762),
.A2(n_522),
.B(n_526),
.C(n_478),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_653),
.A2(n_522),
.B(n_526),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_742),
.A2(n_478),
.B(n_498),
.C(n_522),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_700),
.A2(n_526),
.B(n_498),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_671),
.A2(n_498),
.B(n_708),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_682),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_696),
.B(n_626),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_763),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_755),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_668),
.B(n_709),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_743),
.A2(n_782),
.B(n_748),
.C(n_761),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_780),
.A2(n_716),
.B(n_652),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_652),
.A2(n_632),
.B(n_723),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_701),
.B(n_681),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_643),
.A2(n_777),
.B1(n_648),
.B2(n_746),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_721),
.A2(n_727),
.B(n_764),
.Y(n_842)
);

NOR2xp67_ASAP7_75t_L g843 ( 
.A(n_615),
.B(n_679),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_670),
.A2(n_678),
.B1(n_722),
.B2(n_702),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_762),
.A2(n_775),
.B(n_657),
.C(n_734),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_622),
.A2(n_624),
.B(n_643),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_619),
.B(n_621),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_682),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_625),
.B(n_634),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_725),
.A2(n_726),
.B(n_665),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_L g851 ( 
.A(n_687),
.B(n_676),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_647),
.B(n_691),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_737),
.A2(n_629),
.B(n_631),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_743),
.A2(n_782),
.B(n_748),
.C(n_761),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_639),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_645),
.B(n_650),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_623),
.A2(n_745),
.B(n_778),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_739),
.A2(n_664),
.B(n_693),
.C(n_689),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_737),
.A2(n_628),
.B(n_656),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_658),
.B(n_675),
.Y(n_860)
);

OAI321xp33_ASAP7_75t_L g861 ( 
.A1(n_768),
.A2(n_677),
.A3(n_717),
.B1(n_657),
.B2(n_775),
.C(n_770),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_710),
.A2(n_712),
.B(n_691),
.C(n_751),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_L g863 ( 
.A(n_750),
.B(n_672),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_654),
.A2(n_744),
.B(n_756),
.Y(n_864)
);

BUFx12f_ASAP7_75t_L g865 ( 
.A(n_695),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_758),
.A2(n_781),
.B(n_730),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_701),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_673),
.B(n_663),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_698),
.B(n_699),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_648),
.B(n_740),
.Y(n_870)
);

NAND2x1_ASAP7_75t_L g871 ( 
.A(n_662),
.B(n_705),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_710),
.A2(n_712),
.B(n_692),
.C(n_729),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_636),
.A2(n_638),
.B(n_706),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_740),
.B(n_686),
.Y(n_874)
);

O2A1O1Ixp5_ASAP7_75t_L g875 ( 
.A1(n_767),
.A2(n_776),
.B(n_774),
.C(n_773),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_686),
.B(n_614),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_695),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_690),
.A2(n_684),
.B(n_674),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_704),
.A2(n_760),
.B(n_637),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_642),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_614),
.A2(n_733),
.B(n_730),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_769),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_754),
.A2(n_753),
.B(n_738),
.C(n_733),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_689),
.A2(n_697),
.B(n_693),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_697),
.B(n_618),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_620),
.B(n_765),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_703),
.Y(n_887)
);

BUFx2_ASAP7_75t_L g888 ( 
.A(n_659),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_644),
.B(n_649),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_685),
.B(n_713),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_736),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_724),
.A2(n_740),
.B(n_752),
.Y(n_892)
);

NAND2x1p5_ASAP7_75t_L g893 ( 
.A(n_740),
.B(n_695),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_659),
.B(n_720),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_740),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_L g896 ( 
.A(n_659),
.B(n_635),
.C(n_669),
.Y(n_896)
);

AO21x1_ASAP7_75t_L g897 ( 
.A1(n_740),
.A2(n_688),
.B(n_707),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_766),
.A2(n_641),
.B(n_783),
.Y(n_898)
);

OR2x6_ASAP7_75t_L g899 ( 
.A(n_659),
.B(n_695),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_741),
.A2(n_762),
.B(n_711),
.C(n_775),
.Y(n_900)
);

AO21x1_ASAP7_75t_L g901 ( 
.A1(n_641),
.A2(n_711),
.B(n_616),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_633),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_641),
.B(n_655),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_641),
.B(n_655),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_661),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_641),
.A2(n_783),
.B(n_616),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_771),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_661),
.B(n_718),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_661),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_741),
.A2(n_762),
.B(n_711),
.C(n_775),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_757),
.A2(n_521),
.B1(n_762),
.B2(n_741),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_661),
.B(n_718),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_655),
.A2(n_616),
.B1(n_732),
.B2(n_728),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_640),
.B(n_694),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_661),
.B(n_718),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_714),
.B(n_365),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_771),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_626),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_616),
.A2(n_782),
.B(n_742),
.C(n_748),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_641),
.B(n_655),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_641),
.A2(n_783),
.B(n_616),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_641),
.B(n_655),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_640),
.B(n_397),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_640),
.B(n_694),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_661),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_641),
.B(n_655),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_626),
.Y(n_938)
);

OAI321xp33_ASAP7_75t_L g939 ( 
.A1(n_768),
.A2(n_493),
.A3(n_668),
.B1(n_757),
.B2(n_677),
.C(n_717),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_771),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_661),
.B(n_718),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_640),
.B(n_694),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_641),
.B(n_655),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_641),
.B(n_655),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_661),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_661),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_641),
.B(n_655),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_633),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_616),
.A2(n_641),
.B1(n_718),
.B2(n_643),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_741),
.A2(n_762),
.B(n_711),
.C(n_775),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_741),
.A2(n_762),
.B(n_711),
.C(n_775),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_641),
.B(n_655),
.Y(n_955)
);

AO21x1_ASAP7_75t_L g956 ( 
.A1(n_641),
.A2(n_711),
.B(n_616),
.Y(n_956)
);

AO21x1_ASAP7_75t_L g957 ( 
.A1(n_641),
.A2(n_711),
.B(n_616),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_771),
.Y(n_958)
);

NAND3xp33_ASAP7_75t_L g959 ( 
.A(n_711),
.B(n_640),
.C(n_657),
.Y(n_959)
);

AO21x1_ASAP7_75t_L g960 ( 
.A1(n_641),
.A2(n_711),
.B(n_616),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_633),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_771),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_641),
.B(n_655),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_641),
.A2(n_655),
.B(n_783),
.C(n_473),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_715),
.A2(n_641),
.B(n_779),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_641),
.B(n_655),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_640),
.B(n_397),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_823),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_SL g971 ( 
.A(n_784),
.B(n_835),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_823),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_906),
.A2(n_917),
.B(n_916),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_900),
.A2(n_953),
.B(n_954),
.C(n_911),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_855),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_903),
.B(n_904),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_918),
.A2(n_924),
.B(n_920),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_887),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_807),
.Y(n_979)
);

NAND3xp33_ASAP7_75t_L g980 ( 
.A(n_852),
.B(n_959),
.C(n_911),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_928),
.B(n_930),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_811),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_807),
.Y(n_983)
);

AOI211x1_ASAP7_75t_L g984 ( 
.A1(n_898),
.A2(n_841),
.B(n_936),
.C(n_968),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_931),
.B(n_969),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_925),
.A2(n_934),
.B(n_927),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_945),
.B(n_946),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_935),
.A2(n_943),
.B(n_937),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_832),
.Y(n_990)
);

AOI21xp33_ASAP7_75t_L g991 ( 
.A1(n_852),
.A2(n_939),
.B(n_861),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_921),
.B(n_880),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_944),
.A2(n_962),
.B(n_952),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_949),
.B(n_955),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_964),
.B(n_869),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_966),
.A2(n_967),
.B(n_951),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_824),
.B(n_848),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_965),
.A2(n_846),
.B(n_907),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_821),
.A2(n_828),
.B(n_820),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_812),
.Y(n_1000)
);

AOI21x1_ASAP7_75t_L g1001 ( 
.A1(n_813),
.A2(n_825),
.B(n_797),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_965),
.A2(n_929),
.B(n_790),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_838),
.A2(n_941),
.B(n_919),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_912),
.A2(n_836),
.B1(n_901),
.B2(n_960),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_926),
.A2(n_859),
.B(n_853),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_902),
.B(n_950),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_909),
.A2(n_941),
.B(n_913),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_815),
.B(n_915),
.Y(n_1008)
);

AOI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_885),
.A2(n_845),
.B(n_858),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_915),
.B(n_932),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_932),
.B(n_942),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_942),
.B(n_833),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_792),
.B(n_914),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_817),
.B(n_876),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_879),
.A2(n_842),
.B(n_788),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_833),
.B(n_889),
.Y(n_1016)
);

AOI221x1_ASAP7_75t_L g1017 ( 
.A1(n_862),
.A2(n_839),
.B1(n_827),
.B2(n_872),
.C(n_881),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_817),
.B(n_786),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_909),
.A2(n_913),
.B(n_919),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_805),
.A2(n_791),
.B(n_870),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_816),
.A2(n_819),
.B(n_831),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_889),
.B(n_832),
.Y(n_1022)
);

AO31x2_ASAP7_75t_L g1023 ( 
.A1(n_956),
.A2(n_957),
.A3(n_803),
.B(n_798),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_857),
.A2(n_830),
.B(n_808),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_870),
.A2(n_785),
.B(n_878),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_843),
.B(n_961),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_873),
.A2(n_837),
.B(n_854),
.Y(n_1027)
);

NAND2x1p5_ASAP7_75t_L g1028 ( 
.A(n_826),
.B(n_933),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_814),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_850),
.A2(n_822),
.B(n_827),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_875),
.A2(n_829),
.B(n_840),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_826),
.B(n_933),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_884),
.A2(n_872),
.B(n_868),
.C(n_883),
.Y(n_1033)
);

AO21x1_ASAP7_75t_L g1034 ( 
.A1(n_810),
.A2(n_874),
.B(n_886),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_847),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_875),
.A2(n_840),
.B(n_795),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_818),
.Y(n_1037)
);

OA22x2_ASAP7_75t_L g1038 ( 
.A1(n_891),
.A2(n_894),
.B1(n_899),
.B2(n_890),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_822),
.A2(n_866),
.B(n_809),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_801),
.A2(n_803),
.B(n_874),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_834),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_883),
.A2(n_892),
.B(n_851),
.C(n_800),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_923),
.B(n_938),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_798),
.A2(n_882),
.A3(n_849),
.B(n_856),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_789),
.A2(n_793),
.B(n_799),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_860),
.B(n_963),
.Y(n_1046)
);

AO31x2_ASAP7_75t_L g1047 ( 
.A1(n_897),
.A2(n_867),
.A3(n_802),
.B(n_940),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_958),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_793),
.A2(n_871),
.B(n_922),
.Y(n_1049)
);

AOI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_804),
.A2(n_908),
.B(n_844),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_787),
.B(n_948),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_863),
.A2(n_947),
.B(n_806),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_806),
.A2(n_905),
.B1(n_910),
.B2(n_823),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_802),
.A2(n_893),
.B(n_896),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_823),
.A2(n_910),
.B(n_877),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_910),
.A2(n_877),
.B1(n_899),
.B2(n_888),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_899),
.B(n_865),
.Y(n_1057)
);

OAI22x1_ASAP7_75t_L g1058 ( 
.A1(n_852),
.A2(n_959),
.B1(n_680),
.B2(n_513),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_784),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_906),
.A2(n_917),
.B(n_916),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_903),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_811),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_906),
.A2(n_917),
.B(n_916),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_903),
.B(n_904),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_823),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_824),
.B(n_848),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_895),
.B(n_823),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_903),
.B(n_904),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_903),
.B(n_904),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_824),
.B(n_848),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_784),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_903),
.B(n_904),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_921),
.B(n_495),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_855),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_965),
.A2(n_846),
.B(n_900),
.Y(n_1075)
);

OAI22x1_ASAP7_75t_L g1076 ( 
.A1(n_852),
.A2(n_959),
.B1(n_680),
.B2(n_513),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_921),
.B(n_495),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_835),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_903),
.B(n_904),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_823),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_824),
.B(n_848),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_903),
.B(n_904),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_903),
.B(n_904),
.Y(n_1087)
);

INVx4_ASAP7_75t_L g1088 ( 
.A(n_823),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_965),
.A2(n_846),
.B(n_900),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_965),
.A2(n_846),
.B(n_900),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_931),
.B(n_969),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_835),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_790),
.A2(n_803),
.B(n_798),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_903),
.B(n_904),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_903),
.B(n_904),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_900),
.A2(n_953),
.B(n_954),
.C(n_911),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_823),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_835),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_912),
.A2(n_904),
.B1(n_928),
.B2(n_903),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_807),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_903),
.B(n_904),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_811),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_855),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_900),
.A2(n_953),
.B(n_954),
.C(n_911),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_823),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_864),
.A2(n_796),
.B(n_794),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_975),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1010),
.B(n_1008),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1074),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_1092),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_985),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_1057),
.B(n_1038),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_978),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1106),
.Y(n_1118)
);

BUFx12f_ASAP7_75t_L g1119 ( 
.A(n_1037),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_982),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1082),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1011),
.B(n_1012),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_976),
.B(n_987),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_994),
.B(n_1064),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_1073),
.B(n_1077),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1078),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1100),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1082),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_1059),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_997),
.B(n_1006),
.Y(n_1130)
);

O2A1O1Ixp5_ASAP7_75t_L g1131 ( 
.A1(n_991),
.A2(n_1009),
.B(n_1089),
.C(n_1090),
.Y(n_1131)
);

INVx3_ASAP7_75t_SL g1132 ( 
.A(n_992),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1091),
.B(n_1016),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_1017),
.A2(n_1097),
.A3(n_1107),
.B(n_974),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1068),
.A2(n_1072),
.B1(n_1096),
.B2(n_1069),
.Y(n_1135)
);

OAI21xp33_ASAP7_75t_L g1136 ( 
.A1(n_1011),
.A2(n_995),
.B(n_1012),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1100),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1080),
.A2(n_1086),
.B1(n_1104),
.B2(n_1094),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1071),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_979),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1087),
.B(n_1035),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1061),
.B(n_1102),
.Y(n_1142)
);

OA21x2_ASAP7_75t_L g1143 ( 
.A1(n_1075),
.A2(n_998),
.B(n_1005),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1000),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1145)
);

O2A1O1Ixp5_ASAP7_75t_SL g1146 ( 
.A1(n_1002),
.A2(n_1054),
.B(n_981),
.C(n_1050),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1061),
.B(n_981),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1082),
.Y(n_1148)
);

OR2x2_ASAP7_75t_L g1149 ( 
.A(n_1046),
.B(n_979),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_984),
.B(n_980),
.Y(n_1150)
);

INVx6_ASAP7_75t_L g1151 ( 
.A(n_1043),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_997),
.B(n_1006),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1014),
.B(n_1018),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1004),
.A2(n_1033),
.B1(n_1013),
.B2(n_1038),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_990),
.Y(n_1155)
);

INVx4_ASAP7_75t_SL g1156 ( 
.A(n_1067),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1029),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1004),
.B(n_1042),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1041),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_990),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1103),
.A2(n_1056),
.B(n_983),
.C(n_1027),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1030),
.A2(n_1020),
.B1(n_996),
.B2(n_1027),
.Y(n_1162)
);

O2A1O1Ixp5_ASAP7_75t_SL g1163 ( 
.A1(n_1053),
.A2(n_970),
.B(n_1065),
.C(n_1103),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1098),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1007),
.B(n_1019),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1066),
.B(n_1070),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1062),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1066),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1070),
.B(n_1084),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1084),
.B(n_1105),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1048),
.Y(n_1171)
);

AOI222xp33_ASAP7_75t_L g1172 ( 
.A1(n_1058),
.A2(n_1076),
.B1(n_971),
.B2(n_1051),
.C1(n_1067),
.C2(n_970),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1034),
.B(n_1052),
.Y(n_1173)
);

CKINVDCx8_ASAP7_75t_R g1174 ( 
.A(n_1098),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_977),
.A2(n_1063),
.B(n_986),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1109),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1047),
.B(n_1065),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1047),
.Y(n_1178)
);

OR2x2_ASAP7_75t_SL g1179 ( 
.A(n_1109),
.B(n_1093),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1047),
.B(n_1044),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_L g1181 ( 
.A(n_1052),
.B(n_972),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1025),
.B(n_1020),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1047),
.B(n_972),
.Y(n_1183)
);

NAND2x1_ASAP7_75t_L g1184 ( 
.A(n_1067),
.B(n_1088),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1028),
.B(n_1032),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1109),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1109),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1088),
.B(n_1028),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1055),
.B(n_1025),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_988),
.A2(n_1060),
.B(n_993),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1045),
.B(n_1003),
.Y(n_1191)
);

NAND2x1_ASAP7_75t_L g1192 ( 
.A(n_1067),
.B(n_1049),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1032),
.B(n_1023),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_1023),
.B(n_1045),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1003),
.B(n_1039),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1093),
.Y(n_1196)
);

NAND2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1036),
.B(n_1031),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1023),
.B(n_1049),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1024),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1040),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1021),
.B(n_1040),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_999),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1039),
.B(n_1030),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1060),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1001),
.B(n_1015),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_989),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1079),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1081),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1083),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1085),
.A2(n_1095),
.B(n_1099),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1101),
.B(n_1108),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1110),
.B(n_826),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1010),
.B(n_1008),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_976),
.B(n_987),
.Y(n_1214)
);

CKINVDCx11_ASAP7_75t_R g1215 ( 
.A(n_978),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1082),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1011),
.B(n_694),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_973),
.A2(n_986),
.B(n_977),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1010),
.B(n_1008),
.Y(n_1219)
);

NAND2x1p5_ASAP7_75t_L g1220 ( 
.A(n_972),
.B(n_826),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_976),
.B(n_987),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_SL g1222 ( 
.A1(n_1075),
.A2(n_852),
.B(n_512),
.C(n_516),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_976),
.B(n_987),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_975),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_991),
.A2(n_954),
.B(n_900),
.C(n_953),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1010),
.B(n_1008),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_997),
.B(n_1006),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_991),
.A2(n_954),
.B(n_900),
.C(n_953),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_997),
.B(n_1006),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_1059),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1082),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_975),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_976),
.B(n_987),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_976),
.B(n_987),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_976),
.B(n_987),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_975),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_SL g1237 ( 
.A(n_1059),
.B(n_511),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1010),
.B(n_1008),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_975),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1138),
.B(n_1123),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1178),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1118),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1122),
.A2(n_1217),
.B1(n_1136),
.B2(n_1125),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1179),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1123),
.B(n_1124),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1132),
.A2(n_1133),
.B1(n_1135),
.B2(n_1154),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1135),
.A2(n_1154),
.B1(n_1115),
.B2(n_1116),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1236),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1112),
.B(n_1213),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1239),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1115),
.A2(n_1116),
.B1(n_1219),
.B2(n_1226),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1215),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1165),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1114),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1124),
.B(n_1214),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1214),
.B(n_1221),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1111),
.Y(n_1257)
);

INVx6_ASAP7_75t_L g1258 ( 
.A(n_1156),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1121),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1155),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1230),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1113),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1156),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1160),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1224),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1232),
.Y(n_1266)
);

BUFx12f_ASAP7_75t_L g1267 ( 
.A(n_1129),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1157),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1130),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1158),
.A2(n_1145),
.B1(n_1221),
.B2(n_1223),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_1139),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1223),
.B(n_1233),
.Y(n_1272)
);

CKINVDCx8_ASAP7_75t_R g1273 ( 
.A(n_1130),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1210),
.A2(n_1211),
.B(n_1175),
.Y(n_1274)
);

NAND3xp33_ASAP7_75t_L g1275 ( 
.A(n_1222),
.B(n_1225),
.C(n_1228),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1196),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1159),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1120),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_SL g1279 ( 
.A1(n_1158),
.A2(n_1233),
.B1(n_1235),
.B2(n_1234),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1144),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1234),
.A2(n_1235),
.B1(n_1141),
.B2(n_1116),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1167),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1238),
.A2(n_1172),
.B1(n_1150),
.B2(n_1153),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1149),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1156),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1147),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1153),
.B(n_1152),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1119),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1147),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1146),
.A2(n_1131),
.B(n_1142),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1172),
.A2(n_1150),
.B1(n_1151),
.B2(n_1168),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1177),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1161),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1192),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1184),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1151),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1185),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1170),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1140),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1204),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1200),
.Y(n_1301)
);

AOI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1211),
.A2(n_1218),
.B(n_1190),
.Y(n_1302)
);

AO21x1_ASAP7_75t_SL g1303 ( 
.A1(n_1142),
.A2(n_1203),
.B(n_1195),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1140),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1186),
.Y(n_1305)
);

BUFx8_ASAP7_75t_L g1306 ( 
.A(n_1127),
.Y(n_1306)
);

BUFx4f_ASAP7_75t_SL g1307 ( 
.A(n_1117),
.Y(n_1307)
);

INVx6_ASAP7_75t_L g1308 ( 
.A(n_1166),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1114),
.Y(n_1309)
);

CKINVDCx11_ASAP7_75t_R g1310 ( 
.A(n_1174),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1183),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1137),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1169),
.B(n_1229),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1134),
.B(n_1198),
.Y(n_1314)
);

BUFx2_ASAP7_75t_R g1315 ( 
.A(n_1191),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1134),
.B(n_1180),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1182),
.A2(n_1162),
.B(n_1203),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1227),
.A2(n_1229),
.B1(n_1171),
.B2(n_1126),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1121),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1227),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1197),
.A2(n_1207),
.B(n_1212),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1143),
.A2(n_1237),
.B1(n_1193),
.B2(n_1201),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1143),
.A2(n_1173),
.B1(n_1199),
.B2(n_1194),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1134),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1199),
.A2(n_1195),
.B1(n_1189),
.B2(n_1185),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1185),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1176),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1205),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1188),
.A2(n_1181),
.B1(n_1176),
.B2(n_1231),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1128),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1206),
.A2(n_1209),
.B(n_1163),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1164),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1212),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1202),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1231),
.A2(n_1220),
.B(n_1208),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1148),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1208),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1187),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1220),
.B(n_1187),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1187),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1275),
.A2(n_1216),
.B(n_1243),
.Y(n_1341)
);

AO21x2_ASAP7_75t_L g1342 ( 
.A1(n_1290),
.A2(n_1274),
.B(n_1302),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1314),
.B(n_1316),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1314),
.B(n_1316),
.Y(n_1344)
);

BUFx4f_ASAP7_75t_L g1345 ( 
.A(n_1258),
.Y(n_1345)
);

INVxp33_ASAP7_75t_L g1346 ( 
.A(n_1249),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1324),
.Y(n_1347)
);

INVx3_ASAP7_75t_SL g1348 ( 
.A(n_1258),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1245),
.B(n_1256),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1260),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1253),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1260),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1252),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1326),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1264),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1245),
.B(n_1256),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1311),
.B(n_1292),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1328),
.B(n_1276),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1264),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1326),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1303),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1303),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1293),
.A2(n_1279),
.B(n_1255),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1309),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1241),
.B(n_1323),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1327),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1317),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1244),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1240),
.B(n_1272),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1241),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1244),
.Y(n_1371)
);

AO31x2_ASAP7_75t_L g1372 ( 
.A1(n_1334),
.A2(n_1301),
.A3(n_1337),
.B(n_1300),
.Y(n_1372)
);

CKINVDCx10_ASAP7_75t_R g1373 ( 
.A(n_1252),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1286),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1289),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1301),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1240),
.B(n_1300),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1262),
.B(n_1265),
.Y(n_1378)
);

INVxp33_ASAP7_75t_L g1379 ( 
.A(n_1313),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1287),
.B(n_1307),
.Y(n_1380)
);

CKINVDCx6p67_ASAP7_75t_R g1381 ( 
.A(n_1310),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1310),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1320),
.B(n_1254),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1266),
.B(n_1322),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1246),
.A2(n_1270),
.B(n_1283),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1337),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1321),
.A2(n_1294),
.B(n_1335),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1331),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1333),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1247),
.B(n_1284),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1257),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1331),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1325),
.A2(n_1251),
.B(n_1305),
.Y(n_1393)
);

OAI22x1_ASAP7_75t_L g1394 ( 
.A1(n_1329),
.A2(n_1304),
.B1(n_1299),
.B2(n_1297),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1331),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1281),
.A2(n_1277),
.B(n_1268),
.Y(n_1396)
);

AO21x2_ASAP7_75t_L g1397 ( 
.A1(n_1242),
.A2(n_1248),
.B(n_1250),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1330),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1330),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1278),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1280),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1298),
.B(n_1282),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1387),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1347),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1361),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1392),
.A2(n_1291),
.B(n_1332),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1365),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1343),
.B(n_1338),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1343),
.B(n_1338),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1369),
.B(n_1312),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1344),
.B(n_1340),
.Y(n_1411)
);

INVxp67_ASAP7_75t_L g1412 ( 
.A(n_1398),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1344),
.B(n_1340),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1392),
.B(n_1318),
.Y(n_1414)
);

INVxp67_ASAP7_75t_R g1415 ( 
.A(n_1387),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1395),
.B(n_1336),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1399),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1351),
.B(n_1295),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1370),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1370),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1385),
.A2(n_1308),
.B1(n_1269),
.B2(n_1306),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1345),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1350),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1372),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1372),
.Y(n_1425)
);

AND2x4_ASAP7_75t_SL g1426 ( 
.A(n_1361),
.B(n_1285),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1395),
.B(n_1388),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1362),
.B(n_1263),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1342),
.B(n_1259),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1342),
.B(n_1259),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1342),
.B(n_1259),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1388),
.B(n_1259),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1388),
.B(n_1259),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1363),
.A2(n_1315),
.B(n_1339),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1367),
.B(n_1319),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1365),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1434),
.A2(n_1341),
.B(n_1379),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1434),
.B(n_1390),
.C(n_1364),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1407),
.B(n_1384),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1410),
.B(n_1352),
.Y(n_1440)
);

OAI221xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1421),
.A2(n_1390),
.B1(n_1410),
.B2(n_1436),
.C(n_1407),
.Y(n_1441)
);

OAI221xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1421),
.A2(n_1377),
.B1(n_1371),
.B2(n_1368),
.C(n_1381),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1423),
.B(n_1355),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1422),
.A2(n_1273),
.B1(n_1345),
.B2(n_1346),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1422),
.B(n_1362),
.Y(n_1445)
);

AOI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1423),
.A2(n_1394),
.B1(n_1359),
.B2(n_1366),
.C(n_1383),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1407),
.B(n_1384),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1436),
.B(n_1362),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1412),
.B(n_1349),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1436),
.B(n_1362),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1422),
.B(n_1394),
.Y(n_1451)
);

OAI221xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1414),
.A2(n_1368),
.B1(n_1371),
.B2(n_1381),
.C(n_1380),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1426),
.A2(n_1356),
.B(n_1373),
.Y(n_1453)
);

OAI21xp33_ASAP7_75t_L g1454 ( 
.A1(n_1414),
.A2(n_1402),
.B(n_1357),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1417),
.B(n_1374),
.Y(n_1455)
);

OAI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1414),
.A2(n_1273),
.B1(n_1360),
.B2(n_1269),
.C(n_1308),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1408),
.B(n_1357),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1411),
.B(n_1375),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1422),
.A2(n_1393),
.B1(n_1354),
.B2(n_1382),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1422),
.B(n_1345),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1426),
.A2(n_1373),
.B(n_1429),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1413),
.B(n_1376),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1408),
.B(n_1391),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1429),
.B(n_1393),
.C(n_1360),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1408),
.B(n_1391),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1409),
.B(n_1432),
.Y(n_1466)
);

NAND3xp33_ASAP7_75t_L g1467 ( 
.A(n_1406),
.B(n_1401),
.C(n_1400),
.Y(n_1467)
);

NAND3xp33_ASAP7_75t_L g1468 ( 
.A(n_1406),
.B(n_1401),
.C(n_1400),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1409),
.B(n_1396),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1409),
.B(n_1396),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1419),
.B(n_1396),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1432),
.B(n_1358),
.Y(n_1472)
);

NAND4xp25_ASAP7_75t_L g1473 ( 
.A(n_1418),
.B(n_1402),
.C(n_1354),
.D(n_1378),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1406),
.B(n_1306),
.C(n_1393),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1426),
.A2(n_1382),
.B(n_1353),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1419),
.B(n_1397),
.Y(n_1476)
);

NAND3xp33_ASAP7_75t_L g1477 ( 
.A(n_1406),
.B(n_1306),
.C(n_1393),
.Y(n_1477)
);

NAND4xp25_ASAP7_75t_L g1478 ( 
.A(n_1418),
.B(n_1354),
.C(n_1378),
.D(n_1389),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1406),
.B(n_1386),
.C(n_1389),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1420),
.B(n_1397),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1440),
.B(n_1435),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1466),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1449),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1469),
.B(n_1416),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1476),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1448),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1443),
.B(n_1439),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1470),
.B(n_1416),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1448),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1480),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1439),
.B(n_1416),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1447),
.B(n_1430),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1438),
.A2(n_1428),
.B1(n_1348),
.B2(n_1345),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1471),
.Y(n_1494)
);

NOR2xp67_ASAP7_75t_L g1495 ( 
.A(n_1464),
.B(n_1403),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1463),
.B(n_1427),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1450),
.B(n_1405),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1465),
.B(n_1427),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1455),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1462),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1458),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1450),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1457),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1472),
.B(n_1430),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1460),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1457),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1479),
.B(n_1424),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1473),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1454),
.B(n_1431),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1454),
.B(n_1433),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1478),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1479),
.B(n_1425),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1467),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1503),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1494),
.B(n_1446),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1482),
.B(n_1415),
.Y(n_1516)
);

OAI21xp33_ASAP7_75t_L g1517 ( 
.A1(n_1513),
.A2(n_1438),
.B(n_1437),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1503),
.Y(n_1518)
);

NAND4xp75_ASAP7_75t_L g1519 ( 
.A(n_1495),
.B(n_1451),
.C(n_1445),
.D(n_1475),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1493),
.B(n_1459),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1482),
.B(n_1509),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1482),
.B(n_1415),
.Y(n_1522)
);

NAND2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1495),
.B(n_1405),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1482),
.B(n_1415),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1511),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1513),
.B(n_1467),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1508),
.A2(n_1444),
.B1(n_1474),
.B2(n_1477),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1507),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1483),
.A2(n_1477),
.B1(n_1474),
.B2(n_1468),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1509),
.B(n_1425),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1490),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_L g1532 ( 
.A(n_1490),
.B(n_1468),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1505),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1506),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1506),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1491),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1491),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1499),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1507),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1496),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1499),
.B(n_1404),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1512),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1498),
.Y(n_1544)
);

NOR2xp67_ASAP7_75t_L g1545 ( 
.A(n_1512),
.B(n_1461),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1523),
.B(n_1486),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1517),
.A2(n_1456),
.B1(n_1510),
.B2(n_1502),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1519),
.A2(n_1452),
.B1(n_1442),
.B2(n_1441),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1523),
.B(n_1486),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1523),
.B(n_1489),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1514),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1517),
.B(n_1525),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1521),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1526),
.B(n_1484),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1526),
.B(n_1488),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1525),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1528),
.B(n_1488),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1528),
.B(n_1539),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1514),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1528),
.B(n_1485),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1523),
.B(n_1489),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1545),
.B(n_1489),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1539),
.B(n_1485),
.Y(n_1565)
);

AOI32xp33_ASAP7_75t_L g1566 ( 
.A1(n_1529),
.A2(n_1510),
.A3(n_1502),
.B1(n_1497),
.B2(n_1492),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1545),
.B(n_1502),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1518),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1521),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1536),
.B(n_1504),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1515),
.B(n_1500),
.Y(n_1571)
);

NAND2x1p5_ASAP7_75t_L g1572 ( 
.A(n_1532),
.B(n_1405),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1520),
.A2(n_1453),
.B(n_1501),
.C(n_1487),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1518),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1538),
.B(n_1497),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1533),
.B(n_1288),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1519),
.A2(n_1497),
.B1(n_1481),
.B2(n_1500),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1533),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1538),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1534),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1538),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1532),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1536),
.B(n_1504),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1534),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1535),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1533),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1586),
.B(n_1288),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1557),
.B(n_1515),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1552),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1578),
.B(n_1537),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1552),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1582),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1548),
.B(n_1543),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1564),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1568),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1553),
.B(n_1537),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1559),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1571),
.B(n_1547),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1559),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1572),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1568),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1564),
.B(n_1540),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1567),
.B(n_1540),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1567),
.B(n_1541),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1582),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1575),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_L g1607 ( 
.A(n_1573),
.B(n_1543),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1572),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1549),
.A2(n_1527),
.B1(n_1529),
.B2(n_1544),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1580),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1580),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1548),
.B(n_1555),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1577),
.A2(n_1544),
.B1(n_1541),
.B2(n_1530),
.Y(n_1613)
);

INVxp67_ASAP7_75t_SL g1614 ( 
.A(n_1572),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1579),
.B(n_1542),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1585),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1579),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1555),
.B(n_1542),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1560),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1551),
.B(n_1530),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1574),
.Y(n_1622)
);

AOI21xp33_ASAP7_75t_L g1623 ( 
.A1(n_1607),
.A2(n_1581),
.B(n_1566),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1607),
.A2(n_1576),
.B(n_1581),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1606),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1612),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1609),
.B(n_1570),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1587),
.B(n_1267),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1570),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1589),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1594),
.B(n_1575),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1606),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1594),
.B(n_1583),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1602),
.B(n_1575),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1612),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1589),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1591),
.Y(n_1637)
);

NOR3xp33_ASAP7_75t_L g1638 ( 
.A(n_1588),
.B(n_1563),
.C(n_1554),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1613),
.A2(n_1562),
.B(n_1551),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1618),
.B(n_1583),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1591),
.Y(n_1641)
);

OAI211xp5_ASAP7_75t_L g1642 ( 
.A1(n_1614),
.A2(n_1550),
.B(n_1546),
.C(n_1554),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1595),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1608),
.A2(n_1562),
.B1(n_1550),
.B2(n_1546),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1590),
.Y(n_1645)
);

NOR2x1p5_ASAP7_75t_L g1646 ( 
.A(n_1596),
.B(n_1267),
.Y(n_1646)
);

AOI21xp33_ASAP7_75t_SL g1647 ( 
.A1(n_1593),
.A2(n_1556),
.B(n_1558),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1626),
.B(n_1602),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1635),
.B(n_1597),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1635),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1625),
.B(n_1603),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1641),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1631),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1625),
.B(n_1603),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1631),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1641),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1630),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1623),
.A2(n_1605),
.B1(n_1592),
.B2(n_1620),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1632),
.B(n_1627),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1632),
.B(n_1604),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1636),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1637),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1624),
.B(n_1604),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1645),
.B(n_1605),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1643),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1634),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1629),
.B(n_1621),
.Y(n_1667)
);

AOI222xp33_ASAP7_75t_L g1668 ( 
.A1(n_1658),
.A2(n_1639),
.B1(n_1642),
.B2(n_1633),
.C1(n_1640),
.C2(n_1646),
.Y(n_1668)
);

NAND4xp25_ASAP7_75t_L g1669 ( 
.A(n_1658),
.B(n_1644),
.C(n_1638),
.D(n_1628),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1663),
.A2(n_1647),
.B1(n_1634),
.B2(n_1599),
.C(n_1597),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1659),
.A2(n_1608),
.B(n_1628),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1664),
.A2(n_1599),
.B(n_1597),
.Y(n_1672)
);

AOI21xp33_ASAP7_75t_L g1673 ( 
.A1(n_1653),
.A2(n_1599),
.B(n_1593),
.Y(n_1673)
);

AOI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1655),
.A2(n_1600),
.B(n_1622),
.C(n_1620),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1666),
.B(n_1621),
.Y(n_1675)
);

OAI222xp33_ASAP7_75t_L g1676 ( 
.A1(n_1648),
.A2(n_1600),
.B1(n_1619),
.B2(n_1615),
.C1(n_1556),
.C2(n_1563),
.Y(n_1676)
);

OAI21xp33_ASAP7_75t_L g1677 ( 
.A1(n_1666),
.A2(n_1619),
.B(n_1622),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1668),
.B(n_1651),
.Y(n_1678)
);

AOI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1669),
.A2(n_1660),
.B(n_1649),
.C(n_1654),
.Y(n_1679)
);

NOR2xp67_ASAP7_75t_L g1680 ( 
.A(n_1672),
.B(n_1649),
.Y(n_1680)
);

NOR2x1_ASAP7_75t_L g1681 ( 
.A(n_1671),
.B(n_1650),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1675),
.B(n_1650),
.Y(n_1682)
);

NOR3x1_ASAP7_75t_L g1683 ( 
.A(n_1674),
.B(n_1667),
.C(n_1661),
.Y(n_1683)
);

NOR2x1_ASAP7_75t_L g1684 ( 
.A(n_1676),
.B(n_1652),
.Y(n_1684)
);

NOR3x1_ASAP7_75t_L g1685 ( 
.A(n_1670),
.B(n_1662),
.C(n_1657),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1677),
.Y(n_1686)
);

AOI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1678),
.A2(n_1673),
.B1(n_1665),
.B2(n_1656),
.C(n_1617),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1680),
.B(n_1595),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_L g1689 ( 
.A(n_1681),
.B(n_1601),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1684),
.A2(n_1600),
.B1(n_1616),
.B2(n_1611),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1682),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1689),
.B(n_1685),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1688),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1691),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1690),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1687),
.A2(n_1686),
.B1(n_1679),
.B2(n_1683),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1689),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1692),
.B(n_1601),
.Y(n_1698)
);

OAI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1696),
.A2(n_1617),
.B1(n_1616),
.B2(n_1611),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1697),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1692),
.B(n_1610),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1693),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1702),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1698),
.Y(n_1704)
);

AND2x2_ASAP7_75t_SL g1705 ( 
.A(n_1700),
.B(n_1696),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1703),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1705),
.B1(n_1695),
.B2(n_1699),
.Y(n_1707)
);

AOI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1705),
.B(n_1693),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1707),
.A2(n_1694),
.B1(n_1704),
.B2(n_1701),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1708),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1709),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1610),
.B1(n_1569),
.B2(n_1271),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1710),
.A2(n_1261),
.B(n_1569),
.Y(n_1713)
);

AOI22x1_ASAP7_75t_L g1714 ( 
.A1(n_1713),
.A2(n_1296),
.B1(n_1271),
.B2(n_1261),
.Y(n_1714)
);

AOI322xp5_ASAP7_75t_L g1715 ( 
.A1(n_1714),
.A2(n_1712),
.A3(n_1584),
.B1(n_1531),
.B2(n_1524),
.C1(n_1522),
.C2(n_1516),
.Y(n_1715)
);

AOI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1584),
.B1(n_1531),
.B2(n_1565),
.C(n_1561),
.Y(n_1716)
);

AOI211xp5_ASAP7_75t_L g1717 ( 
.A1(n_1716),
.A2(n_1271),
.B(n_1565),
.C(n_1561),
.Y(n_1717)
);


endmodule