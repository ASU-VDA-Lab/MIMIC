module fake_jpeg_1966_n_232 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_232);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_1),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_81),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_0),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_54),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_2),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_70),
.B1(n_56),
.B2(n_65),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_97),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_55),
.B1(n_68),
.B2(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_55),
.B1(n_68),
.B2(n_72),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_59),
.B(n_71),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_71),
.B(n_61),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_65),
.B1(n_64),
.B2(n_62),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_114),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_77),
.B1(n_73),
.B2(n_76),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_115),
.B1(n_57),
.B2(n_7),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_63),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_113),
.Y(n_122)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_61),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_64),
.B1(n_82),
.B2(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_2),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_3),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_4),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_94),
.C(n_79),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_125),
.C(n_137),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_98),
.B1(n_79),
.B2(n_80),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_25),
.B1(n_51),
.B2(n_47),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_75),
.C(n_74),
.Y(n_125)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_126),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_57),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_26),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_75),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_74),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_138),
.B(n_9),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_100),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_149),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_112),
.B1(n_111),
.B2(n_105),
.Y(n_145)
);

OAI22x1_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_146),
.A2(n_157),
.B(n_15),
.Y(n_176)
);

AO22x1_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_99),
.B1(n_27),
.B2(n_28),
.Y(n_147)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_155),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_24),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_12),
.C(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_11),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_130),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_159),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_12),
.B(n_13),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_139),
.B(n_138),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_170),
.B(n_176),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_153),
.A2(n_120),
.B1(n_126),
.B2(n_119),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_175),
.B1(n_158),
.B2(n_18),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_162),
.A2(n_125),
.B1(n_29),
.B2(n_31),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_181),
.B(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_162),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_34),
.B(n_45),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_141),
.B(n_156),
.C(n_143),
.D(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_32),
.C(n_44),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_147),
.B1(n_151),
.B2(n_161),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_191),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_158),
.B(n_19),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_190),
.A2(n_196),
.B(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_194),
.B(n_195),
.Y(n_200)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_20),
.B(n_21),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_198),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_165),
.C(n_166),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_207),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_179),
.B(n_178),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_174),
.C(n_173),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_182),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.C(n_193),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_183),
.C(n_175),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.Y(n_220)
);

NAND4xp25_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_216),
.C(n_218),
.D(n_200),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_203),
.A2(n_194),
.B1(n_197),
.B2(n_186),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_171),
.Y(n_222)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

AO221x1_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_186),
.B1(n_195),
.B2(n_205),
.C(n_206),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_222),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_213),
.B(n_216),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_214),
.C(n_212),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_223),
.B(n_224),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_220),
.Y(n_227)
);

OAI321xp33_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_225),
.A3(n_40),
.B1(n_41),
.B2(n_42),
.C(n_43),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_52),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_22),
.Y(n_232)
);


endmodule