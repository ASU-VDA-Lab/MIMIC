module fake_jpeg_10662_n_273 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_62),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_60),
.B1(n_25),
.B2(n_24),
.Y(n_96)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_34),
.B(n_25),
.Y(n_92)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NAND2x1_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_33),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_33),
.B(n_25),
.C(n_24),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_26),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_18),
.B1(n_29),
.B2(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_21),
.B1(n_33),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_61),
.B1(n_63),
.B2(n_23),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_26),
.C(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_66),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_18),
.B1(n_32),
.B2(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_17),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_18),
.B1(n_31),
.B2(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_24),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_100),
.C(n_46),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_40),
.B1(n_33),
.B2(n_25),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_46),
.B1(n_65),
.B2(n_3),
.Y(n_107)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_71),
.B(n_94),
.Y(n_119)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_73),
.A2(n_76),
.B1(n_86),
.B2(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_34),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_34),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_77),
.Y(n_109)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

CKINVDCx6p67_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_81),
.B(n_88),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_85),
.A2(n_97),
.B1(n_101),
.B2(n_16),
.Y(n_120)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_34),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_6),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_0),
.C(n_2),
.Y(n_113)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_128)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_68),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_58),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_46),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_107),
.A2(n_87),
.B1(n_73),
.B2(n_101),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_120),
.B1(n_128),
.B2(n_76),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_102),
.Y(n_139)
);

XOR2x1_ASAP7_75t_SL g153 ( 
.A(n_113),
.B(n_79),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_94),
.B1(n_91),
.B2(n_80),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_82),
.B(n_71),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_6),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_69),
.B(n_7),
.C(n_8),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_97),
.C(n_9),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_129),
.B(n_118),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_104),
.B1(n_115),
.B2(n_109),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_99),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_140),
.C(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_132),
.B(n_133),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_127),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_147),
.B(n_155),
.Y(n_166)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_106),
.B(n_88),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_139),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_72),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_156),
.B1(n_158),
.B2(n_142),
.Y(n_172)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_111),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_100),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_157),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_79),
.C(n_70),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NOR2xp67_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_89),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_126),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_181),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_178),
.B(n_179),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_125),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_136),
.C(n_138),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_104),
.B1(n_106),
.B2(n_103),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_168),
.A2(n_170),
.B1(n_173),
.B2(n_176),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_105),
.B1(n_109),
.B2(n_116),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_116),
.B1(n_98),
.B2(n_128),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_117),
.B(n_79),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_117),
.B(n_124),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_124),
.B(n_121),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_133),
.A2(n_95),
.B1(n_78),
.B2(n_75),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_156),
.B1(n_158),
.B2(n_121),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_135),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_197),
.C(n_199),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_135),
.Y(n_191)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_163),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_195),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_151),
.Y(n_196)
);

AOI21x1_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_198),
.B(n_205),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_150),
.C(n_149),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_168),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_171),
.B1(n_175),
.B2(n_183),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_159),
.B(n_147),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_148),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_167),
.C(n_160),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_210),
.C(n_214),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_174),
.C(n_179),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_181),
.C(n_165),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_186),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_174),
.C(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_173),
.C(n_165),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_219),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_165),
.C(n_171),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_176),
.B1(n_86),
.B2(n_84),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_186),
.B(n_195),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_217),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_192),
.B(n_191),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_224),
.A2(n_236),
.B1(n_222),
.B2(n_187),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_230),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_232),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_185),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_196),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_206),
.C(n_210),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_242),
.C(n_243),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_8),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_206),
.C(n_214),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_209),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_246),
.C(n_231),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_221),
.C(n_212),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_185),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_196),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_246),
.A2(n_236),
.B(n_226),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_234),
.B(n_227),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_9),
.B(n_10),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_253),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_254),
.C(n_248),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_230),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_201),
.C(n_198),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_245),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_255),
.C(n_89),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_250),
.A2(n_240),
.B1(n_237),
.B2(n_245),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_260),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_258),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_84),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_264),
.A2(n_259),
.B1(n_260),
.B2(n_256),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_268),
.A3(n_265),
.B1(n_262),
.B2(n_13),
.C1(n_14),
.C2(n_16),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_257),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_10),
.C2(n_15),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_269),
.B1(n_12),
.B2(n_13),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_11),
.Y(n_273)
);


endmodule