module fake_jpeg_29902_n_371 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_371);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_371;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_4),
.B(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_45),
.B(n_50),
.Y(n_116)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_46),
.Y(n_102)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_21),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_53),
.Y(n_103)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_9),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_59),
.B(n_17),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_74),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_24),
.B(n_9),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_26),
.B(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_71),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_26),
.B(n_10),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_20),
.C(n_19),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_79),
.B(n_17),
.C(n_16),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_87),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_42),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_93),
.A2(n_98),
.B1(n_36),
.B2(n_35),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_47),
.A2(n_38),
.B1(n_40),
.B2(n_37),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_117),
.B1(n_121),
.B2(n_123),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_28),
.B1(n_30),
.B2(n_37),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_37),
.B1(n_33),
.B2(n_40),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_113),
.B1(n_119),
.B2(n_0),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_43),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_43),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_108),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_50),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_38),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_112),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_37),
.B1(n_40),
.B2(n_18),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_44),
.B1(n_32),
.B2(n_29),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_66),
.A2(n_44),
.B1(n_32),
.B2(n_29),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_35),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_45),
.A2(n_44),
.B1(n_29),
.B2(n_27),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_35),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_122),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_45),
.A2(n_44),
.B1(n_27),
.B2(n_22),
.Y(n_123)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_126),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_18),
.B(n_27),
.C(n_22),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_22),
.B1(n_18),
.B2(n_36),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_0),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_137),
.Y(n_171)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_96),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_36),
.B1(n_35),
.B2(n_12),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_142),
.B1(n_144),
.B2(n_150),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_147),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_36),
.B1(n_12),
.B2(n_13),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_36),
.B1(n_17),
.B2(n_16),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_81),
.B(n_0),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_133),
.Y(n_172)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_151),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_162),
.B1(n_129),
.B2(n_87),
.Y(n_178)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_155),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_101),
.A2(n_15),
.B(n_1),
.C(n_2),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_86),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_112),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_156),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_116),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_159),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_163),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_113),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_97),
.B1(n_85),
.B2(n_88),
.Y(n_187)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_8),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_174),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_119),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_79),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_87),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_178),
.A2(n_193),
.B1(n_197),
.B2(n_126),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_88),
.B1(n_97),
.B2(n_114),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_182),
.A2(n_187),
.B1(n_191),
.B2(n_159),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_89),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_189),
.C(n_198),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_89),
.C(n_106),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_114),
.B1(n_85),
.B2(n_82),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_194),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_99),
.B1(n_82),
.B2(n_90),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_162),
.A2(n_99),
.B1(n_106),
.B2(n_78),
.Y(n_193)
);

AO22x2_ASAP7_75t_L g194 ( 
.A1(n_127),
.A2(n_103),
.B1(n_84),
.B2(n_80),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_136),
.A2(n_84),
.B1(n_90),
.B2(n_80),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_202),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_143),
.A2(n_80),
.B1(n_103),
.B2(n_108),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_103),
.C(n_80),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_7),
.C(n_8),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_173),
.C(n_174),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_137),
.B(n_158),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_208),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_177),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_211),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_135),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_214),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_124),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_215),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_128),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_217),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_147),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_131),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_220),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_139),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_155),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_221),
.B(n_236),
.Y(n_258)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_194),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_SL g262 ( 
.A(n_224),
.B(n_231),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_134),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_225),
.B(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_229),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_168),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_171),
.B(n_148),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_168),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_194),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_165),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_192),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_156),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_234),
.B(n_235),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_243),
.B(n_257),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_178),
.C(n_196),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_259),
.C(n_209),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_242),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_196),
.B(n_175),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_SL g244 ( 
.A1(n_214),
.A2(n_154),
.A3(n_167),
.B1(n_197),
.B2(n_193),
.C1(n_199),
.C2(n_194),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_244),
.B(n_163),
.CI(n_153),
.CON(n_282),
.SN(n_282)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_192),
.B(n_200),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_250),
.B(n_179),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_192),
.B(n_195),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_260),
.B(n_218),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_167),
.B1(n_187),
.B2(n_190),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_160),
.B1(n_180),
.B2(n_151),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_206),
.A2(n_169),
.B(n_185),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_209),
.B(n_184),
.C(n_185),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_179),
.B(n_169),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_236),
.A2(n_138),
.B(n_146),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_225),
.B(n_227),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_221),
.A2(n_179),
.B1(n_160),
.B2(n_159),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_254),
.B1(n_261),
.B2(n_257),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_205),
.A3(n_219),
.B1(n_212),
.B2(n_204),
.C1(n_207),
.C2(n_220),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_266),
.A2(n_274),
.B(n_265),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_268),
.C(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_210),
.C(n_204),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_242),
.B(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g272 ( 
.A1(n_241),
.A2(n_205),
.A3(n_213),
.B1(n_212),
.B2(n_218),
.C1(n_217),
.C2(n_231),
.Y(n_272)
);

NOR3xp33_ASAP7_75t_SL g307 ( 
.A(n_272),
.B(n_287),
.C(n_262),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_273),
.B(n_276),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_252),
.B(n_232),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_289),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_232),
.B1(n_203),
.B2(n_228),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_226),
.C(n_215),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_280),
.A2(n_245),
.B1(n_250),
.B2(n_246),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_222),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_249),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_8),
.Y(n_283)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_237),
.A2(n_248),
.B(n_245),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_285),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_240),
.C(n_253),
.Y(n_286)
);

OAI321xp33_ASAP7_75t_L g287 ( 
.A1(n_245),
.A2(n_238),
.A3(n_263),
.B1(n_262),
.B2(n_258),
.C(n_248),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_265),
.C(n_241),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_268),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_249),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_279),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_291),
.B(n_292),
.Y(n_325)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_279),
.A2(n_245),
.B1(n_250),
.B2(n_244),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_303),
.B(n_273),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_309),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_280),
.A2(n_250),
.B1(n_256),
.B2(n_248),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_282),
.Y(n_315)
);

AOI321xp33_ASAP7_75t_L g308 ( 
.A1(n_269),
.A2(n_255),
.A3(n_260),
.B1(n_246),
.B2(n_251),
.C(n_247),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_308),
.A2(n_281),
.B(n_283),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_286),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_275),
.C(n_289),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_311),
.B(n_317),
.C(n_318),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_294),
.B(n_288),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_315),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_278),
.B(n_270),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_319),
.B(n_297),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_271),
.C(n_282),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_277),
.C(n_284),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_301),
.A2(n_278),
.B(n_270),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_321),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_277),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_297),
.A2(n_274),
.B1(n_287),
.B2(n_276),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_322),
.A2(n_303),
.B1(n_295),
.B2(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_305),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_323),
.Y(n_328)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_323),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_302),
.C(n_298),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_331),
.B(n_334),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_332),
.A2(n_335),
.B1(n_308),
.B2(n_266),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_299),
.C(n_290),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_322),
.A2(n_320),
.B1(n_316),
.B2(n_324),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_316),
.A2(n_299),
.B1(n_307),
.B2(n_306),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_326),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_293),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_337),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_325),
.B(n_313),
.Y(n_340)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_340),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_318),
.B(n_317),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_343),
.B(n_345),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_330),
.A2(n_319),
.B(n_314),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_334),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_333),
.A2(n_311),
.B(n_285),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_346),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_332),
.Y(n_353)
);

NOR2x1_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_321),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_339),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_327),
.C(n_331),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_352),
.A2(n_356),
.B(n_353),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_353),
.A2(n_357),
.B1(n_349),
.B2(n_348),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_345),
.B(n_327),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_356),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_335),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_359),
.B(n_361),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_351),
.A2(n_354),
.B1(n_358),
.B2(n_329),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_364),
.C(n_337),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_358),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_362),
.B(n_352),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_366),
.C(n_328),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g370 ( 
.A1(n_368),
.A2(n_369),
.B(n_357),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_367),
.B(n_363),
.C(n_329),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_339),
.Y(n_371)
);


endmodule