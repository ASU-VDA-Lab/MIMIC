module fake_aes_12658_n_20 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_20);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_7;
BUFx6f_ASAP7_75t_L g7 ( .A(n_2), .Y(n_7) );
INVx3_ASAP7_75t_L g8 ( .A(n_1), .Y(n_8) );
OA21x2_ASAP7_75t_L g9 ( .A1(n_3), .A2(n_5), .B(n_6), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_8), .B(n_0), .Y(n_10) );
BUFx3_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
OAI21x1_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_9), .B(n_4), .Y(n_12) );
INVx1_ASAP7_75t_SL g13 ( .A(n_12), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_14), .B(n_11), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
XNOR2xp5_ASAP7_75t_L g19 ( .A(n_18), .B(n_7), .Y(n_19) );
INVx2_ASAP7_75t_SL g20 ( .A(n_19), .Y(n_20) );
endmodule