module fake_jpeg_32176_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_2),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx6f_ASAP7_75t_SL g71 ( 
.A(n_26),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_84),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_59),
.B1(n_62),
.B2(n_75),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_91),
.B1(n_99),
.B2(n_57),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_59),
.B1(n_75),
.B2(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_73),
.Y(n_93)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_63),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_70),
.B1(n_53),
.B2(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_52),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_52),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_71),
.B1(n_54),
.B2(n_70),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_112),
.B1(n_7),
.B2(n_8),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_53),
.B1(n_74),
.B2(n_55),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_117),
.B1(n_29),
.B2(n_50),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_64),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_114),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_56),
.B1(n_64),
.B2(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_76),
.B1(n_2),
.B2(n_3),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_21),
.B1(n_49),
.B2(n_48),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_22),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_134),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_3),
.B(n_4),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_10),
.B(n_11),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_4),
.C(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_136),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_6),
.B(n_7),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_24),
.C(n_41),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_122),
.C(n_139),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_8),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_10),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_40),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_149),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_28),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_125),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_155),
.A2(n_156),
.B(n_133),
.Y(n_163)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_30),
.A3(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_158),
.B(n_19),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_161),
.B1(n_119),
.B2(n_141),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_162),
.A2(n_165),
.B1(n_166),
.B2(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_167),
.C(n_158),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_135),
.B(n_121),
.Y(n_165)
);

NAND4xp25_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_127),
.C(n_120),
.D(n_128),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_154),
.C(n_146),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_174),
.C(n_168),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_142),
.C(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_147),
.B1(n_173),
.B2(n_152),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_147),
.B1(n_159),
.B2(n_161),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_170),
.B(n_151),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_177),
.B1(n_164),
.B2(n_165),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_145),
.B(n_150),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_166),
.B(n_136),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_31),
.C(n_32),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_185),
.B(n_39),
.Y(n_186)
);


endmodule