module fake_jpeg_23472_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_23),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_64),
.Y(n_97)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_51),
.Y(n_77)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_55),
.Y(n_81)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_35),
.B1(n_16),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_67),
.B1(n_35),
.B2(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_35),
.B1(n_16),
.B2(n_28),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_75),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_92),
.B1(n_96),
.B2(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_94),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_74),
.A2(n_89),
.B1(n_95),
.B2(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_79),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_37),
.B1(n_39),
.B2(n_18),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_78),
.A2(n_93),
.B1(n_91),
.B2(n_70),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_21),
.Y(n_82)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_84),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_66),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_30),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_44),
.B1(n_42),
.B2(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_22),
.Y(n_125)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_12),
.C(n_15),
.Y(n_135)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_36),
.B1(n_29),
.B2(n_20),
.Y(n_126)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_43),
.C(n_38),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_107),
.C(n_29),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_64),
.B(n_39),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_45),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_112),
.A2(n_113),
.B(n_134),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_72),
.A2(n_22),
.B(n_37),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_128),
.C(n_77),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_129),
.B1(n_136),
.B2(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_22),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_44),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_42),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_33),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_88),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_0),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_9),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_95),
.A2(n_20),
.B1(n_32),
.B2(n_31),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_84),
.A2(n_33),
.B1(n_34),
.B2(n_32),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_80),
.B1(n_108),
.B2(n_100),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_151),
.C(n_150),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_141),
.B1(n_159),
.B2(n_127),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_130),
.B1(n_131),
.B2(n_110),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_142),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_81),
.B(n_17),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_148),
.B(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_157),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_149),
.B1(n_153),
.B2(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_117),
.B(n_73),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_84),
.B1(n_69),
.B2(n_80),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_102),
.B(n_108),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_84),
.C(n_103),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_98),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_152),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_83),
.B1(n_87),
.B2(n_79),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_32),
.B1(n_27),
.B2(n_34),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_17),
.B(n_27),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_158),
.B(n_168),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_31),
.B1(n_27),
.B2(n_17),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_31),
.B(n_88),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_161),
.A2(n_170),
.B1(n_15),
.B2(n_9),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_33),
.B(n_1),
.Y(n_162)
);

NOR2x1_ASAP7_75t_R g191 ( 
.A(n_162),
.B(n_1),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_0),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_1),
.Y(n_173)
);

AO22x1_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_33),
.B1(n_90),
.B2(n_88),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_165),
.A2(n_138),
.B1(n_121),
.B2(n_137),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_120),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_169),
.Y(n_174)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_1),
.B(n_2),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_191),
.B(n_200),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_189),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_169),
.A2(n_124),
.B1(n_109),
.B2(n_121),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_175),
.A2(n_195),
.B1(n_141),
.B2(n_142),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_179),
.C(n_182),
.Y(n_224)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_177),
.B(n_181),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_119),
.C(n_116),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_119),
.C(n_116),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_147),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_194),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_123),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_127),
.B1(n_123),
.B2(n_4),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_143),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_9),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_162),
.B(n_166),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_144),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_159),
.B1(n_140),
.B2(n_155),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_3),
.C(n_4),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_11),
.C(n_13),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_170),
.B1(n_149),
.B2(n_145),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_204),
.A2(n_220),
.B1(n_226),
.B2(n_173),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_206),
.A2(n_230),
.B1(n_209),
.B2(n_205),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_207),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_151),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_179),
.Y(n_233)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_211),
.B(n_216),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_212),
.Y(n_250)
);

NAND2x1_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_143),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_219),
.B(n_229),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_178),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_225),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_197),
.A2(n_146),
.B(n_157),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_192),
.A2(n_156),
.B1(n_164),
.B2(n_167),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_222),
.Y(n_252)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_164),
.B1(n_154),
.B2(n_8),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_164),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_203),
.C(n_180),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g231 ( 
.A(n_198),
.Y(n_231)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_245),
.C(n_256),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_235),
.B(n_222),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_180),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_239),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_171),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_199),
.A3(n_188),
.B1(n_172),
.B2(n_186),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_204),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_210),
.A2(n_197),
.B(n_185),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_241),
.A2(n_213),
.B(n_227),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_171),
.B1(n_177),
.B2(n_202),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_242),
.A2(n_247),
.B1(n_226),
.B2(n_217),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_195),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_191),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_249),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_187),
.B1(n_173),
.B2(n_8),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_232),
.B1(n_214),
.B2(n_229),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_205),
.B(n_10),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_209),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_218),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_10),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_250),
.Y(n_257)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_273),
.C(n_245),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_276),
.B1(n_244),
.B2(n_204),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_269),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_254),
.A2(n_214),
.B1(n_216),
.B2(n_212),
.Y(n_267)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_220),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_221),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_270),
.B(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_234),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_246),
.B(n_243),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_230),
.C(n_223),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_237),
.A2(n_211),
.B1(n_204),
.B2(n_207),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_275),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_242),
.B(n_223),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_238),
.B1(n_234),
.B2(n_248),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_283),
.B1(n_291),
.B2(n_11),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_281),
.C(n_285),
.Y(n_302)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_258),
.B(n_259),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_235),
.C(n_236),
.Y(n_281)
);

XOR2x1_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_240),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_263),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_256),
.B1(n_247),
.B2(n_249),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_228),
.C(n_7),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_294),
.B(n_298),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_303),
.CI(n_285),
.CON(n_311),
.SN(n_311)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_297),
.B(n_300),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_290),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_291),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_277),
.B(n_268),
.CI(n_262),
.CON(n_299),
.SN(n_299)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_301),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_292),
.A2(n_257),
.B(n_262),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_283),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_11),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_278),
.C(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_307),
.C(n_14),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_300),
.C(n_304),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_289),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_306),
.B(n_308),
.Y(n_317)
);

NOR2x1_ASAP7_75t_R g315 ( 
.A(n_311),
.B(n_299),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_284),
.B(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_293),
.B1(n_280),
.B2(n_299),
.Y(n_314)
);

NAND2x1p5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_319),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g321 ( 
.A(n_319),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_321),
.A2(n_320),
.B(n_315),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_316),
.B(n_311),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_318),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_317),
.B(n_322),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_305),
.C(n_307),
.Y(n_328)
);


endmodule