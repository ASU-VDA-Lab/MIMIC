module fake_jpeg_3369_n_530 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_530);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_46),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_1),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_49),
.B(n_24),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_50),
.Y(n_139)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_52),
.Y(n_143)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_53),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_95),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx2_ASAP7_75t_R g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_24),
.Y(n_100)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_96),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_100),
.B(n_125),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_46),
.A2(n_21),
.B1(n_33),
.B2(n_37),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_113),
.A2(n_74),
.B1(n_69),
.B2(n_19),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_47),
.A2(n_24),
.B1(n_32),
.B2(n_15),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_114),
.A2(n_128),
.B1(n_136),
.B2(n_155),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_40),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_116),
.B(n_117),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_55),
.B(n_40),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_71),
.B(n_43),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_88),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_55),
.B(n_43),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_123),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_24),
.B1(n_15),
.B2(n_27),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_67),
.A2(n_24),
.B1(n_15),
.B2(n_27),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_70),
.B(n_42),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_142),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_70),
.B(n_94),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_94),
.A2(n_42),
.B1(n_39),
.B2(n_23),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_77),
.A2(n_39),
.B1(n_44),
.B2(n_18),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_157),
.A2(n_75),
.B1(n_44),
.B2(n_17),
.Y(n_202)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_167),
.Y(n_208)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_97),
.B(n_72),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_162),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_79),
.B1(n_91),
.B2(n_85),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_163),
.A2(n_164),
.B1(n_177),
.B2(n_183),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_59),
.B1(n_66),
.B2(n_52),
.Y(n_164)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_102),
.B(n_72),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_166),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_115),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_107),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_169),
.B(n_180),
.Y(n_235)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_103),
.B(n_33),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_110),
.B(n_37),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_84),
.B1(n_83),
.B2(n_81),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_179),
.A2(n_143),
.B1(n_17),
.B2(n_133),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_107),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_186),
.Y(n_223)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_96),
.B1(n_18),
.B2(n_19),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_135),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_156),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_192),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_21),
.B1(n_37),
.B2(n_76),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_196),
.B1(n_17),
.B2(n_119),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_111),
.B(n_37),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_101),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_195),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_99),
.A2(n_44),
.B1(n_19),
.B2(n_18),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_197),
.Y(n_236)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_200),
.A2(n_138),
.B1(n_137),
.B2(n_119),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_202),
.A2(n_75),
.B1(n_137),
.B2(n_118),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_180),
.B1(n_169),
.B2(n_190),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_209),
.A2(n_203),
.B1(n_101),
.B2(n_197),
.Y(n_259)
);

AO22x2_ASAP7_75t_L g211 ( 
.A1(n_164),
.A2(n_128),
.B1(n_136),
.B2(n_114),
.Y(n_211)
);

AO21x2_ASAP7_75t_L g243 ( 
.A1(n_211),
.A2(n_221),
.B(n_231),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_127),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_226),
.C(n_166),
.Y(n_240)
);

BUFx8_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_162),
.B(n_106),
.C(n_151),
.Y(n_226)
);

AOI32xp33_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_149),
.A3(n_130),
.B1(n_138),
.B2(n_112),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_166),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_162),
.A2(n_133),
.B1(n_126),
.B2(n_141),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_195),
.B1(n_158),
.B2(n_172),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_167),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_241),
.B(n_264),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_171),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_265),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_209),
.A2(n_179),
.B1(n_204),
.B2(n_174),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_253),
.B1(n_257),
.B2(n_258),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_204),
.C(n_160),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_246),
.B(n_250),
.C(n_267),
.Y(n_298)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_248),
.Y(n_293)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_204),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_256),
.B(n_269),
.Y(n_290)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_228),
.B(n_203),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_266),
.B(n_207),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_160),
.B(n_191),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_192),
.B1(n_203),
.B2(n_193),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_218),
.A2(n_203),
.B1(n_184),
.B2(n_168),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_262),
.B1(n_231),
.B2(n_205),
.Y(n_280)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_261),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_219),
.A2(n_131),
.B1(n_141),
.B2(n_126),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_229),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_268),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_234),
.B(n_189),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_234),
.B(n_194),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_232),
.A2(n_170),
.B(n_178),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_228),
.C(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_SL g269 ( 
.A(n_237),
.B(n_178),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_241),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_271),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_264),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_276),
.C(n_284),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_246),
.C(n_240),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_213),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_279),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_278),
.A2(n_281),
.B(n_288),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_244),
.B(n_213),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_243),
.B1(n_258),
.B2(n_262),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_211),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_227),
.C(n_223),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_250),
.B(n_236),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_254),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_243),
.A2(n_211),
.B1(n_221),
.B2(n_223),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_294),
.B1(n_243),
.B2(n_257),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_223),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_263),
.Y(n_291)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_291),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_255),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_220),
.C(n_199),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_211),
.B1(n_223),
.B2(n_214),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_252),
.B(n_236),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_297),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_253),
.Y(n_299)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_299),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_272),
.B(n_245),
.Y(n_300)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_295),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_301),
.B(n_312),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_302),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_280),
.B1(n_288),
.B2(n_292),
.Y(n_336)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_243),
.B1(n_255),
.B2(n_242),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_275),
.A2(n_243),
.B1(n_211),
.B2(n_247),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_291),
.A2(n_247),
.B1(n_205),
.B2(n_249),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_275),
.A2(n_211),
.B1(n_247),
.B2(n_260),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_311),
.A2(n_314),
.B1(n_324),
.B2(n_328),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_295),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_313),
.B(n_319),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_247),
.B1(n_268),
.B2(n_248),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_SL g315 ( 
.A(n_272),
.B(n_233),
.C(n_205),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_176),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_270),
.A2(n_261),
.B1(n_230),
.B2(n_224),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_318),
.A2(n_330),
.B(n_288),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_271),
.B(n_230),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_279),
.B(n_214),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_322),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_277),
.B(n_214),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_292),
.B(n_298),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_285),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_278),
.A2(n_206),
.B1(n_165),
.B2(n_200),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_296),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_173),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_217),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_331),
.C(n_298),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_283),
.A2(n_224),
.B1(n_198),
.B2(n_181),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_220),
.B1(n_215),
.B2(n_210),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_293),
.B1(n_215),
.B2(n_210),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_186),
.B(n_238),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_316),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_336),
.A2(n_341),
.B1(n_350),
.B2(n_351),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_276),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_338),
.B(n_342),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_344),
.C(n_357),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_309),
.A2(n_289),
.B1(n_286),
.B2(n_282),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_340),
.A2(n_305),
.B1(n_358),
.B2(n_313),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_304),
.A2(n_274),
.B1(n_289),
.B2(n_284),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_323),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_284),
.C(n_285),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_273),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_124),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_318),
.Y(n_346)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_346),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_348),
.B(n_326),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_308),
.A2(n_282),
.B1(n_293),
.B2(n_283),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_317),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_352),
.B(n_361),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_302),
.A2(n_182),
.B1(n_175),
.B2(n_161),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_353),
.A2(n_354),
.B1(n_360),
.B2(n_303),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_SL g355 ( 
.A(n_312),
.B(n_176),
.Y(n_355)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_314),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_149),
.C(n_120),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_140),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_359),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_301),
.A2(n_139),
.B1(n_188),
.B2(n_144),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_317),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_300),
.A2(n_187),
.B(n_139),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_176),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_320),
.Y(n_364)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

NAND4xp25_ASAP7_75t_SL g395 ( 
.A(n_366),
.B(n_356),
.C(n_335),
.D(n_355),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_369),
.A2(n_379),
.B1(n_392),
.B2(n_346),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_326),
.C(n_319),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_372),
.C(n_376),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_371),
.B(n_378),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_321),
.C(n_311),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_374),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_341),
.B(n_306),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_384),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_322),
.C(n_325),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_345),
.B(n_306),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_334),
.A2(n_332),
.B1(n_324),
.B2(n_316),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_329),
.C(n_332),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_393),
.C(n_359),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_108),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_336),
.A2(n_315),
.B1(n_303),
.B2(n_131),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_382),
.A2(n_362),
.B1(n_359),
.B2(n_368),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_333),
.B(n_315),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_340),
.B(n_140),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_387),
.Y(n_408)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_388),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_333),
.B(n_303),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_389),
.B(n_391),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_349),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_337),
.A2(n_98),
.B1(n_132),
.B2(n_80),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_86),
.C(n_48),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_353),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_395),
.B(n_1),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_410),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_357),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_404),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_401),
.A2(n_382),
.B1(n_379),
.B2(n_368),
.Y(n_428)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_347),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_403),
.Y(n_430)
);

XNOR2x2_ASAP7_75t_SL g404 ( 
.A(n_388),
.B(n_347),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_363),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_412),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_411),
.A2(n_419),
.B1(n_390),
.B2(n_392),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_350),
.C(n_356),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_364),
.C(n_343),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_4),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_360),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_386),
.Y(n_435)
);

AO221x1_ASAP7_75t_L g415 ( 
.A1(n_369),
.A2(n_343),
.B1(n_124),
.B2(n_108),
.C(n_21),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_415),
.B(n_4),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_416),
.B(n_380),
.Y(n_423)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_367),
.A2(n_30),
.B1(n_2),
.B2(n_4),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_377),
.B(n_371),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_378),
.Y(n_434)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_421),
.Y(n_437)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_423),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_407),
.A2(n_383),
.B(n_366),
.Y(n_425)
);

CKINVDCx14_ASAP7_75t_R g455 ( 
.A(n_425),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_393),
.C(n_394),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_436),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_428),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_429),
.A2(n_433),
.B1(n_409),
.B2(n_5),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_399),
.A2(n_381),
.B(n_386),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_431),
.A2(n_4),
.B(n_5),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_418),
.A2(n_411),
.B1(n_400),
.B2(n_404),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_434),
.B(n_441),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_435),
.B(n_442),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_25),
.C(n_4),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_438),
.A2(n_6),
.B(n_7),
.Y(n_465)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_419),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_440),
.Y(n_457)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_396),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_413),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g460 ( 
.A(n_443),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_30),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_6),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_30),
.B1(n_5),
.B2(n_6),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_445),
.A2(n_408),
.B1(n_397),
.B2(n_395),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_430),
.Y(n_447)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_447),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_431),
.A2(n_412),
.B(n_416),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_448),
.A2(n_428),
.B(n_426),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_410),
.C(n_414),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_451),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_420),
.C(n_409),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_463),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_454),
.A2(n_436),
.B1(n_9),
.B2(n_10),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_SL g471 ( 
.A(n_456),
.B(n_437),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_446),
.B(n_5),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_458),
.B(n_8),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_461),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_438),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_25),
.C(n_7),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_465),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_433),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_470),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_473),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_427),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_SL g474 ( 
.A(n_449),
.B(n_427),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_474),
.A2(n_466),
.B(n_452),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_432),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_475),
.B(n_476),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_444),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_462),
.B(n_435),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_478),
.A2(n_482),
.B1(n_465),
.B2(n_461),
.Y(n_491)
);

OAI21xp33_ASAP7_75t_SL g484 ( 
.A1(n_479),
.A2(n_480),
.B(n_481),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_454),
.A2(n_429),
.B(n_434),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_448),
.A2(n_423),
.B(n_445),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_453),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_488),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_472),
.A2(n_450),
.B1(n_451),
.B2(n_466),
.Y(n_486)
);

XOR2x2_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_492),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_479),
.A2(n_453),
.B(n_450),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_497),
.B(n_483),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_460),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_25),
.C(n_9),
.Y(n_508)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_491),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_473),
.B(n_464),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_458),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_498),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_456),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_496),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_471),
.A2(n_459),
.B(n_30),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_30),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_508),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_495),
.A2(n_489),
.B(n_486),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_500),
.A2(n_503),
.B(n_8),
.Y(n_514)
);

OAI321xp33_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_492),
.A3(n_484),
.B1(n_496),
.B2(n_468),
.C(n_482),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_484),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g518 ( 
.A(n_506),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_25),
.C(n_9),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_509),
.B(n_510),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_489),
.A2(n_25),
.B1(n_9),
.B2(n_10),
.Y(n_510)
);

NOR3xp33_ASAP7_75t_L g511 ( 
.A(n_504),
.B(n_8),
.C(n_9),
.Y(n_511)
);

O2A1O1Ixp33_ASAP7_75t_SL g523 ( 
.A1(n_511),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_501),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_512),
.A2(n_514),
.B(n_516),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_11),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_515),
.A2(n_518),
.B(n_513),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_13),
.C(n_11),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_505),
.B(n_507),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_520),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_521),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_517),
.A2(n_505),
.B(n_12),
.Y(n_522)
);

NOR3xp33_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_523),
.C(n_11),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_524),
.B(n_519),
.C(n_12),
.Y(n_528)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_525),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_528),
.B(n_526),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_529),
.A2(n_11),
.B(n_13),
.Y(n_530)
);


endmodule