module fake_netlist_5_1887_n_1609 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1609);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1609;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_109),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_30),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_37),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_11),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_60),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_41),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_55),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_105),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_32),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_33),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_48),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_8),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_56),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_36),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_32),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_108),
.Y(n_174)
);

BUFx2_ASAP7_75t_SL g175 ( 
.A(n_58),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_26),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_83),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_71),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_49),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_21),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_66),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_2),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_53),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_80),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_152),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_34),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

BUFx8_ASAP7_75t_SL g188 ( 
.A(n_13),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_31),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_31),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_0),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_42),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g194 ( 
.A(n_44),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_20),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_10),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_62),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_81),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_16),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_39),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_4),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_92),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_54),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_119),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_111),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_21),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_67),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_26),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_63),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_34),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_74),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_139),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_96),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_148),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_93),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_77),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_129),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_39),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_8),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_124),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_87),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_99),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_29),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_146),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_16),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_142),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_85),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_127),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_59),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_134),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_145),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_135),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_110),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_6),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_114),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_79),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_45),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_78),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_95),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_1),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_22),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_13),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_143),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_41),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_88),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_70),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_29),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_28),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_25),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_104),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_12),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_140),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_98),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_68),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_76),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_64),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_136),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_22),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_84),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_35),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_73),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_12),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_101),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_72),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_4),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_137),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_47),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_69),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_86),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_123),
.Y(n_275)
);

INVxp33_ASAP7_75t_R g276 ( 
.A(n_133),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_126),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_128),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_18),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_43),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_38),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_122),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_10),
.Y(n_283)
);

BUFx2_ASAP7_75t_SL g284 ( 
.A(n_30),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_61),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_38),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_40),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_42),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_151),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_19),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_103),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_106),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_102),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_113),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_27),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_17),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_51),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_7),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_57),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_188),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_222),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_168),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_180),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_229),
.Y(n_305)
);

INVxp33_ASAP7_75t_SL g306 ( 
.A(n_193),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_191),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_182),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_195),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_247),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_198),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_201),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_212),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_177),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_291),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_155),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_300),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_155),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_156),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_220),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_156),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_199),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_228),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_232),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_205),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_239),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_246),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_206),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_254),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_194),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_157),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_256),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_157),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_208),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_210),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_159),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_190),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_159),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_222),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_272),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_279),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_162),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_211),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_162),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_164),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_164),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_296),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_213),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_170),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_272),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_165),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_153),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_166),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_167),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_172),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_173),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_179),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_183),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_284),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_184),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_204),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_197),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_217),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_170),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_236),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_203),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_302),
.B(n_200),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_185),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_367),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_200),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_355),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_308),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_357),
.Y(n_383)
);

NAND2x1_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_185),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_248),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_315),
.B(n_194),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_248),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_303),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_209),
.B(n_190),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_282),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_312),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_309),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_282),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_310),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_314),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_321),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_324),
.B(n_325),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

CKINVDCx8_ASAP7_75t_R g408 ( 
.A(n_371),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_209),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_334),
.B(n_249),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_338),
.B(n_249),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_244),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

AND2x4_ASAP7_75t_SL g417 ( 
.A(n_317),
.B(n_194),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_320),
.A2(n_299),
.B1(n_176),
.B2(n_171),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_352),
.B(n_187),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_307),
.A2(n_263),
.B(n_187),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_323),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_332),
.B(n_263),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_326),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_318),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_330),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_336),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_337),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_346),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_306),
.A2(n_299),
.B1(n_176),
.B2(n_171),
.Y(n_431)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_305),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_311),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_322),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_322),
.A2(n_252),
.B1(n_230),
.B2(n_253),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_421),
.A2(n_306),
.B1(n_354),
.B2(n_319),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_378),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_189),
.C(n_186),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_376),
.B(n_192),
.Y(n_442)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_423),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_378),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_378),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_381),
.B(n_214),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_422),
.A2(n_354),
.B1(n_319),
.B2(n_223),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_175),
.Y(n_449)
);

INVx8_ASAP7_75t_L g450 ( 
.A(n_426),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_378),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_395),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_393),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_333),
.Y(n_454)
);

OR2x6_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_276),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_381),
.B(n_215),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_426),
.B(n_154),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_216),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_373),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_333),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_373),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_426),
.B(n_154),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_388),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_421),
.A2(n_380),
.B1(n_395),
.B2(n_415),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_395),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_391),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_426),
.B(n_158),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_421),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_377),
.Y(n_473)
);

CKINVDCx6p67_ASAP7_75t_R g474 ( 
.A(n_426),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_380),
.B(n_218),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_339),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g479 ( 
.A(n_419),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_402),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_388),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_428),
.B(n_153),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_L g487 ( 
.A(n_428),
.B(n_153),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_388),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_382),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_383),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_414),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_426),
.B(n_160),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_431),
.B(n_196),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_401),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_421),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_404),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_427),
.B(n_339),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_374),
.B(n_238),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_375),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_421),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_417),
.B(n_311),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_374),
.A2(n_266),
.B1(n_153),
.B2(n_262),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_375),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_407),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_SL g511 ( 
.A(n_387),
.B(n_230),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_427),
.B(n_341),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_379),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_390),
.B(n_219),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_379),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_414),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_401),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_419),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_390),
.B(n_224),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_401),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_428),
.B(n_160),
.Y(n_522)
);

OR2x6_ASAP7_75t_L g523 ( 
.A(n_433),
.B(n_266),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_432),
.B(n_341),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_384),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_401),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_374),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_397),
.A2(n_234),
.B1(n_261),
.B2(n_369),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_389),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_386),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_401),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_401),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_428),
.B(n_430),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_390),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_390),
.Y(n_535)
);

INVxp67_ASAP7_75t_SL g536 ( 
.A(n_384),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_L g538 ( 
.A(n_428),
.B(n_153),
.Y(n_538)
);

AOI21x1_ASAP7_75t_L g539 ( 
.A1(n_385),
.A2(n_271),
.B(n_269),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_414),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_389),
.A2(n_262),
.B1(n_274),
.B2(n_258),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_389),
.B(n_225),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_414),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_432),
.A2(n_253),
.B1(n_270),
.B2(n_252),
.Y(n_544)
);

NOR2x1p5_ASAP7_75t_L g545 ( 
.A(n_429),
.B(n_265),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_403),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_SL g547 ( 
.A(n_436),
.B(n_265),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_389),
.B(n_227),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_396),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_396),
.B(n_231),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_396),
.B(n_242),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_403),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_396),
.B(n_233),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_403),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_405),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_405),
.Y(n_556)
);

AND2x2_ASAP7_75t_SL g557 ( 
.A(n_417),
.B(n_262),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_405),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_400),
.B(n_260),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_431),
.B(n_202),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_409),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_409),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_409),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_432),
.B(n_345),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_432),
.B(n_348),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_430),
.B(n_161),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_411),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_430),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_430),
.A2(n_283),
.B1(n_221),
.B2(n_226),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_418),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_430),
.B(n_348),
.Y(n_572)
);

NAND2x1_ASAP7_75t_L g573 ( 
.A(n_400),
.B(n_262),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_459),
.A2(n_430),
.B1(n_278),
.B2(n_290),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_489),
.B(n_408),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_459),
.B(n_433),
.Y(n_576)
);

O2A1O1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_461),
.A2(n_385),
.B(n_416),
.C(n_406),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_453),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_437),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_461),
.B(n_433),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_568),
.Y(n_581)
);

INVxp67_ASAP7_75t_SL g582 ( 
.A(n_452),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_443),
.B(n_349),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_443),
.B(n_350),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_568),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_447),
.B(n_350),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_525),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_525),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_437),
.B(n_435),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_473),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_471),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_527),
.B(n_420),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_472),
.A2(n_420),
.B1(n_410),
.B2(n_413),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_551),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_529),
.B(n_420),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_465),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_442),
.B(n_435),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_546),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_546),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_465),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_529),
.B(n_420),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_503),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_549),
.B(n_498),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_549),
.B(n_418),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_557),
.B(n_438),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_498),
.B(n_410),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_557),
.B(n_408),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_442),
.B(n_435),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_480),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_SL g611 ( 
.A(n_528),
.B(n_369),
.C(n_316),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_472),
.B(n_412),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_504),
.B(n_412),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_456),
.B(n_161),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_571),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_504),
.B(n_466),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_452),
.A2(n_413),
.B1(n_270),
.B2(n_207),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_570),
.B(n_408),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_455),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_533),
.B(n_534),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_481),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_477),
.B(n_163),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_464),
.B(n_235),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_458),
.B(n_163),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_572),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_535),
.B(n_237),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_441),
.B(n_169),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_551),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_499),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_464),
.B(n_240),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_559),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_522),
.B(n_169),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_500),
.Y(n_633)
);

OAI221xp5_ASAP7_75t_L g634 ( 
.A1(n_541),
.A2(n_406),
.B1(n_286),
.B2(n_287),
.C(n_297),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_467),
.B(n_241),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_524),
.B(n_372),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_566),
.B(n_174),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_571),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_505),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_510),
.B(n_243),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_512),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_502),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_571),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_495),
.B(n_372),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_495),
.B(n_425),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_503),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_509),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_560),
.B(n_174),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_509),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_559),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_491),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_515),
.B(n_520),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_463),
.B(n_250),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_514),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_537),
.B(n_543),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_514),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_516),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_463),
.B(n_251),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_489),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_463),
.B(n_280),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_516),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_468),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_460),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_468),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_537),
.B(n_285),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_470),
.Y(n_666)
);

A2O1A1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_502),
.A2(n_292),
.B(n_293),
.C(n_294),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_449),
.A2(n_295),
.B1(n_298),
.B2(n_178),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_470),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_448),
.B(n_544),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_560),
.B(n_178),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_543),
.B(n_268),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_476),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_476),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_542),
.B(n_181),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_478),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_482),
.Y(n_677)
);

NOR3xp33_ASAP7_75t_L g678 ( 
.A(n_547),
.B(n_181),
.C(n_255),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_475),
.B(n_255),
.Y(n_679)
);

BUFx6f_ASAP7_75t_SL g680 ( 
.A(n_455),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_482),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_506),
.B(n_434),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_548),
.B(n_257),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_564),
.B(n_316),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_502),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_475),
.B(n_257),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_484),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_455),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_484),
.B(n_277),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_449),
.A2(n_277),
.B1(n_275),
.B2(n_273),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_SL g692 ( 
.A(n_565),
.B(n_301),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_550),
.B(n_259),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_449),
.A2(n_275),
.B1(n_273),
.B2(n_268),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_485),
.Y(n_695)
);

BUFx8_ASAP7_75t_L g696 ( 
.A(n_506),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_485),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_475),
.B(n_483),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_483),
.B(n_259),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_493),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_493),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_483),
.B(n_264),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_494),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_494),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_497),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_497),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_488),
.B(n_264),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_488),
.B(n_52),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_488),
.B(n_490),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_556),
.B(n_301),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_513),
.B(n_2),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_553),
.B(n_3),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_486),
.A2(n_7),
.B(n_9),
.C(n_11),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_490),
.B(n_82),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_556),
.B(n_65),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_511),
.B(n_9),
.C(n_14),
.Y(n_716)
);

AOI22x1_ASAP7_75t_L g717 ( 
.A1(n_490),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_508),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_552),
.B(n_100),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_558),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_449),
.B(n_23),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_558),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_554),
.B(n_91),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_562),
.Y(n_724)
);

BUFx5_ASAP7_75t_L g725 ( 
.A(n_507),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_479),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_479),
.A2(n_24),
.B1(n_33),
.B2(n_35),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_473),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_555),
.B(n_115),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_562),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_563),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_511),
.A2(n_523),
.B1(n_457),
.B2(n_462),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_486),
.A2(n_36),
.B(n_37),
.C(n_40),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_536),
.B(n_46),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_561),
.B(n_50),
.Y(n_735)
);

CKINVDCx8_ASAP7_75t_R g736 ( 
.A(n_659),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_SL g737 ( 
.A(n_575),
.B(n_711),
.Y(n_737)
);

INVx6_ASAP7_75t_L g738 ( 
.A(n_696),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_656),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_582),
.B(n_561),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_646),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_686),
.B(n_455),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_625),
.B(n_519),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_663),
.B(n_676),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_602),
.Y(n_745)
);

AO22x2_ASAP7_75t_L g746 ( 
.A1(n_606),
.A2(n_519),
.B1(n_547),
.B2(n_573),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_728),
.B(n_579),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_721),
.B(n_523),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_625),
.A2(n_538),
.B(n_487),
.C(n_492),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_582),
.B(n_616),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_600),
.B(n_569),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_589),
.Y(n_752)
);

NOR2xp67_ASAP7_75t_L g753 ( 
.A(n_663),
.B(n_563),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_619),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_647),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_648),
.A2(n_573),
.B(n_567),
.C(n_569),
.Y(n_756)
);

INVx4_ASAP7_75t_L g757 ( 
.A(n_596),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_596),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_676),
.B(n_469),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_611),
.B(n_487),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_649),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_636),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_609),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_597),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_642),
.B(n_594),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_642),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_654),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_682),
.B(n_545),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_657),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_661),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_602),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_628),
.B(n_507),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_614),
.B(n_530),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_578),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_696),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_614),
.B(n_517),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_622),
.B(n_474),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_596),
.B(n_450),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_622),
.B(n_474),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_662),
.Y(n_780)
);

OR2x2_ASAP7_75t_SL g781 ( 
.A(n_644),
.B(n_540),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_583),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_586),
.A2(n_532),
.B1(n_531),
.B2(n_526),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_624),
.B(n_518),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_591),
.Y(n_785)
);

CKINVDCx6p67_ASAP7_75t_R g786 ( 
.A(n_680),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_682),
.B(n_539),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_651),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_624),
.B(n_521),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_600),
.B(n_593),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_666),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_651),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_712),
.A2(n_538),
.B1(n_491),
.B2(n_446),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_593),
.B(n_446),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_610),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_586),
.A2(n_491),
.B1(n_439),
.B2(n_451),
.Y(n_796)
);

BUFx12f_ASAP7_75t_L g797 ( 
.A(n_689),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_607),
.B(n_451),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_603),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_621),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_629),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_583),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_590),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_648),
.A2(n_491),
.B1(n_444),
.B2(n_440),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_685),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_584),
.B(n_444),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_613),
.B(n_440),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_603),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_584),
.B(n_450),
.Y(n_809)
);

OR2x2_ASAP7_75t_SL g810 ( 
.A(n_645),
.B(n_89),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_633),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_612),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_612),
.B(n_496),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_726),
.A2(n_496),
.B1(n_445),
.B2(n_450),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_674),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_631),
.B(n_90),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_639),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_612),
.B(n_496),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_587),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_641),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_605),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_664),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_688),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_669),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_612),
.B(n_496),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_588),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_650),
.B(n_588),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_675),
.B(n_445),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_673),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_677),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_681),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_612),
.B(n_445),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_695),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_700),
.Y(n_834)
);

BUFx12f_ASAP7_75t_SL g835 ( 
.A(n_734),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_671),
.B(n_107),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_604),
.B(n_445),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_734),
.B(n_576),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_697),
.Y(n_839)
);

OAI22x1_ASAP7_75t_SL g840 ( 
.A1(n_683),
.A2(n_112),
.B1(n_118),
.B2(n_121),
.Y(n_840)
);

OR2x2_ASAP7_75t_SL g841 ( 
.A(n_716),
.B(n_692),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_701),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_617),
.B(n_130),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_617),
.B(n_652),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_675),
.B(n_131),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_SL g846 ( 
.A1(n_726),
.A2(n_141),
.B1(n_147),
.B2(n_149),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_727),
.A2(n_718),
.B1(n_671),
.B2(n_670),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_652),
.B(n_698),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_725),
.B(n_592),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_L g850 ( 
.A(n_694),
.B(n_627),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_684),
.A2(n_693),
.B1(n_627),
.B2(n_732),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_710),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_684),
.B(n_693),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_710),
.B(n_632),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_632),
.A2(n_637),
.B1(n_601),
.B2(n_595),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_703),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_640),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_725),
.B(n_709),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_725),
.B(n_577),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_704),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_637),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_705),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_580),
.B(n_608),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_725),
.B(n_580),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_678),
.B(n_618),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_725),
.B(n_706),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_R g867 ( 
.A(n_680),
.B(n_679),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_690),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_651),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_725),
.B(n_720),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_691),
.B(n_626),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_581),
.B(n_585),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_678),
.B(n_721),
.Y(n_873)
);

BUFx4f_ASAP7_75t_L g874 ( 
.A(n_651),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_581),
.B(n_585),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_687),
.B(n_699),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_702),
.B(n_707),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_623),
.B(n_630),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_722),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_626),
.B(n_668),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_653),
.B(n_658),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_660),
.B(n_724),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_598),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_730),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_731),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_672),
.B(n_690),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_635),
.A2(n_634),
.B1(n_717),
.B2(n_718),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_599),
.B(n_643),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_615),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_672),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_715),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_638),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_713),
.B(n_733),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_708),
.A2(n_620),
.B(n_655),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_655),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_620),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_574),
.B(n_665),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_665),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_715),
.B(n_735),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_719),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_667),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_727),
.A2(n_723),
.B1(n_729),
.B2(n_714),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_586),
.A2(n_625),
.B1(n_606),
.B2(n_734),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_698),
.A2(n_504),
.B(n_498),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_SL g905 ( 
.A(n_611),
.B(n_547),
.C(n_436),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_659),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_582),
.B(n_616),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_582),
.B(n_616),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_861),
.B(n_744),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_906),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_778),
.A2(n_849),
.B(n_878),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_765),
.B(n_742),
.Y(n_912)
);

INVxp33_ASAP7_75t_L g913 ( 
.A(n_803),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_774),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_853),
.B(n_763),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_765),
.B(n_742),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_758),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_847),
.A2(n_743),
.B(n_802),
.C(n_782),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_736),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_775),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_849),
.A2(n_874),
.B(n_740),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_805),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_747),
.B(n_797),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_752),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_R g925 ( 
.A(n_799),
.B(n_808),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_758),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_847),
.A2(n_851),
.B1(n_846),
.B2(n_903),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_821),
.B(n_750),
.Y(n_928)
);

BUFx4f_ASAP7_75t_L g929 ( 
.A(n_786),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_874),
.A2(n_740),
.B(n_881),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_871),
.A2(n_854),
.B(n_844),
.C(n_843),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_844),
.A2(n_843),
.B(n_863),
.C(n_759),
.Y(n_932)
);

O2A1O1Ixp5_ASAP7_75t_L g933 ( 
.A1(n_828),
.A2(n_779),
.B(n_777),
.C(n_836),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_780),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_855),
.A2(n_902),
.B1(n_838),
.B2(n_908),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_907),
.A2(n_908),
.B(n_877),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_788),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_SL g938 ( 
.A1(n_810),
.A2(n_841),
.B1(n_781),
.B2(n_747),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_754),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_757),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_880),
.A2(n_850),
.B(n_890),
.C(n_886),
.Y(n_941)
);

OAI21xp33_ASAP7_75t_L g942 ( 
.A1(n_737),
.A2(n_887),
.B(n_865),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_886),
.A2(n_898),
.B(n_868),
.C(n_876),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_747),
.B(n_738),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_873),
.A2(n_746),
.B1(n_838),
.B2(n_893),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_806),
.B(n_857),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_753),
.B(n_827),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_790),
.A2(n_859),
.B(n_794),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_859),
.A2(n_864),
.B1(n_812),
.B2(n_897),
.Y(n_949)
);

NOR2xp67_ASAP7_75t_L g950 ( 
.A(n_773),
.B(n_784),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_864),
.A2(n_812),
.B1(n_776),
.B2(n_789),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_858),
.A2(n_814),
.B(n_866),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_827),
.B(n_848),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_785),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_738),
.Y(n_955)
);

NOR2xp67_ASAP7_75t_SL g956 ( 
.A(n_812),
.B(n_757),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_848),
.B(n_795),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_812),
.A2(n_858),
.B1(n_896),
.B2(n_900),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_788),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_791),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_819),
.A2(n_826),
.B1(n_870),
.B2(n_866),
.Y(n_961)
);

NAND2xp33_ASAP7_75t_L g962 ( 
.A(n_891),
.B(n_760),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_815),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_766),
.B(n_800),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_814),
.A2(n_870),
.B(n_904),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_882),
.A2(n_751),
.B(n_798),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_768),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_751),
.A2(n_807),
.B(n_798),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_801),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_894),
.A2(n_807),
.B(n_837),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_811),
.B(n_817),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_820),
.B(n_787),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_772),
.B(n_764),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_788),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_737),
.B(n_852),
.Y(n_975)
);

AOI222xp33_ASAP7_75t_L g976 ( 
.A1(n_840),
.A2(n_845),
.B1(n_746),
.B2(n_748),
.C1(n_905),
.C2(n_816),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_822),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_816),
.B(n_792),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_792),
.Y(n_979)
);

CKINVDCx6p67_ASAP7_75t_R g980 ( 
.A(n_901),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_748),
.B(n_867),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_813),
.A2(n_825),
.B(n_818),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_813),
.A2(n_825),
.B(n_832),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_893),
.A2(n_739),
.B(n_756),
.C(n_839),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_832),
.A2(n_875),
.B(n_872),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_823),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_893),
.A2(n_741),
.B1(n_770),
.B2(n_769),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_749),
.A2(n_899),
.B(n_809),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_835),
.B(n_772),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_819),
.B(n_826),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_755),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_761),
.B(n_767),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_833),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_892),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_824),
.Y(n_995)
);

NAND2x1_ASAP7_75t_L g996 ( 
.A(n_869),
.B(n_792),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_891),
.B(n_783),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_891),
.B(n_745),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_829),
.B(n_842),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_771),
.B(n_869),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_830),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_883),
.B(n_860),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_834),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_831),
.B(n_856),
.Y(n_1004)
);

AND2x6_ASAP7_75t_L g1005 ( 
.A(n_895),
.B(n_796),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_888),
.A2(n_793),
.B(n_804),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_884),
.A2(n_885),
.B1(n_862),
.B2(n_879),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_889),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_847),
.A2(n_853),
.B(n_743),
.C(n_802),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_906),
.B(n_659),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_780),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_765),
.B(n_742),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_851),
.A2(n_903),
.B1(n_847),
.B2(n_855),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_747),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_853),
.B(n_625),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_788),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_780),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_861),
.B(n_663),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_851),
.B(n_861),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_758),
.Y(n_1020)
);

CKINVDCx11_ASAP7_75t_R g1021 ( 
.A(n_736),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_853),
.B(n_625),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_762),
.B(n_752),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_851),
.A2(n_903),
.B1(n_847),
.B2(n_855),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_774),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_853),
.B(n_625),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_861),
.B(n_663),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_803),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_SL g1029 ( 
.A1(n_853),
.A2(n_843),
.B(n_606),
.C(n_845),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_762),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_851),
.A2(n_871),
.B(n_847),
.C(n_880),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_861),
.B(n_663),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_778),
.A2(n_582),
.B(n_600),
.Y(n_1033)
);

AND2x2_ASAP7_75t_SL g1034 ( 
.A(n_836),
.B(n_557),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_861),
.B(n_663),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_853),
.B(n_625),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_906),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_758),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_778),
.A2(n_582),
.B(n_600),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_851),
.A2(n_871),
.B(n_847),
.C(n_880),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_847),
.A2(n_851),
.B1(n_853),
.B2(n_846),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_851),
.B(n_861),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_1010),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1031),
.A2(n_1040),
.B(n_931),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_936),
.A2(n_988),
.B(n_911),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_932),
.A2(n_935),
.B(n_1041),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_982),
.A2(n_983),
.B(n_970),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_946),
.B(n_928),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_1041),
.A2(n_927),
.B(n_942),
.C(n_1009),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_909),
.B(n_1019),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_974),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_965),
.A2(n_1039),
.B(n_1033),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1042),
.B(n_1015),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_914),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1013),
.A2(n_1024),
.B(n_952),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_954),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_969),
.Y(n_1057)
);

CKINVDCx11_ASAP7_75t_R g1058 ( 
.A(n_1021),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_L g1059 ( 
.A(n_927),
.B(n_942),
.C(n_918),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1025),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_925),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_941),
.A2(n_943),
.B(n_984),
.C(n_1034),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1018),
.B(n_1027),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_930),
.A2(n_933),
.B(n_948),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_939),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_950),
.A2(n_1006),
.B(n_921),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_1032),
.B(n_1035),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1022),
.B(n_1026),
.Y(n_1068)
);

AO31x2_ASAP7_75t_L g1069 ( 
.A1(n_951),
.A2(n_949),
.A3(n_958),
.B(n_968),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_961),
.A2(n_966),
.A3(n_985),
.B(n_972),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_997),
.A2(n_998),
.B(n_990),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1036),
.B(n_953),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_SL g1073 ( 
.A(n_1014),
.B(n_910),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_957),
.B(n_950),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_976),
.A2(n_975),
.B(n_962),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_924),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_919),
.B(n_920),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1030),
.B(n_913),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_947),
.B(n_987),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_977),
.Y(n_1080)
);

NAND3x1_ASAP7_75t_L g1081 ( 
.A(n_989),
.B(n_1023),
.C(n_915),
.Y(n_1081)
);

AO31x2_ASAP7_75t_L g1082 ( 
.A1(n_999),
.A2(n_1004),
.A3(n_1001),
.B(n_995),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_971),
.B(n_973),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1002),
.A2(n_1007),
.B(n_1000),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_1029),
.A2(n_963),
.A3(n_1017),
.B(n_960),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_978),
.A2(n_987),
.B(n_981),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_974),
.Y(n_1087)
);

OAI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_945),
.A2(n_964),
.B(n_967),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_956),
.B(n_940),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_934),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_992),
.A2(n_1003),
.B(n_993),
.C(n_986),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1011),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1005),
.A2(n_992),
.B(n_994),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_978),
.A2(n_980),
.B1(n_1012),
.B2(n_991),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1012),
.B(n_1008),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1020),
.A2(n_996),
.B(n_959),
.C(n_937),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_959),
.Y(n_1097)
);

OAI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_944),
.A2(n_923),
.B1(n_929),
.B2(n_1037),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_974),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1005),
.A2(n_917),
.B(n_1038),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_1016),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1005),
.B(n_938),
.Y(n_1102)
);

INVx4_ASAP7_75t_L g1103 ( 
.A(n_1016),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_1005),
.A2(n_1016),
.B(n_926),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_979),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_979),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_944),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_1021),
.Y(n_1108)
);

OAI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1031),
.A2(n_851),
.B(n_1040),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_SL g1110 ( 
.A1(n_1013),
.A2(n_853),
.B(n_1024),
.C(n_625),
.Y(n_1110)
);

AOI211x1_ASAP7_75t_L g1111 ( 
.A1(n_942),
.A2(n_847),
.B(n_1024),
.C(n_1013),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_914),
.Y(n_1112)
);

CKINVDCx11_ASAP7_75t_R g1113 ( 
.A(n_1021),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1031),
.A2(n_1040),
.A3(n_1013),
.B(n_1024),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_1031),
.B(n_851),
.C(n_1040),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1010),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_940),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_936),
.A2(n_878),
.B(n_988),
.Y(n_1118)
);

NOR2xp67_ASAP7_75t_SL g1119 ( 
.A(n_955),
.B(n_736),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_982),
.A2(n_983),
.B(n_970),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_946),
.B(n_625),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_914),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1031),
.A2(n_1040),
.B(n_851),
.C(n_1041),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1031),
.A2(n_1040),
.B(n_851),
.C(n_1041),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_1031),
.A2(n_1040),
.A3(n_1013),
.B(n_1024),
.Y(n_1125)
);

AOI221x1_ASAP7_75t_L g1126 ( 
.A1(n_1031),
.A2(n_1040),
.B1(n_1013),
.B2(n_1024),
.C(n_847),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_914),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_974),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_936),
.A2(n_878),
.B(n_988),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_982),
.A2(n_983),
.B(n_970),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1031),
.A2(n_851),
.B(n_1040),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_909),
.B(n_663),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_SL g1133 ( 
.A1(n_1031),
.A2(n_1040),
.B(n_931),
.Y(n_1133)
);

AOI21xp33_ASAP7_75t_L g1134 ( 
.A1(n_1031),
.A2(n_851),
.B(n_847),
.Y(n_1134)
);

AOI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_1031),
.A2(n_851),
.B(n_847),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1031),
.A2(n_851),
.B(n_1040),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_912),
.B(n_916),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_922),
.B(n_752),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_946),
.B(n_625),
.Y(n_1139)
);

AO221x1_ASAP7_75t_L g1140 ( 
.A1(n_1013),
.A2(n_847),
.B1(n_846),
.B2(n_1024),
.C(n_676),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_940),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_974),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_936),
.A2(n_878),
.B(n_988),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_982),
.A2(n_983),
.B(n_970),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1028),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_946),
.B(n_625),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_982),
.A2(n_983),
.B(n_970),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_936),
.A2(n_878),
.B(n_988),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_1031),
.A2(n_1040),
.A3(n_1013),
.B(n_1024),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_936),
.A2(n_878),
.B(n_988),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_982),
.A2(n_983),
.B(n_970),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1031),
.A2(n_1040),
.A3(n_1013),
.B(n_1024),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_946),
.B(n_625),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1031),
.A2(n_1040),
.B(n_851),
.C(n_1041),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_914),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_946),
.B(n_625),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_982),
.A2(n_983),
.B(n_970),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_982),
.A2(n_983),
.B(n_970),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_914),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_988),
.A2(n_1040),
.B(n_1031),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_914),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1031),
.A2(n_851),
.B(n_1040),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_909),
.B(n_663),
.Y(n_1163)
);

AO21x1_ASAP7_75t_L g1164 ( 
.A1(n_1046),
.A2(n_1135),
.B(n_1134),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1064),
.A2(n_1066),
.B(n_1045),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1115),
.A2(n_1109),
.B1(n_1136),
.B2(n_1162),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1068),
.B(n_1053),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1058),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_1044),
.A2(n_1129),
.B(n_1118),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_1089),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_1103),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1065),
.Y(n_1172)
);

INVx6_ASAP7_75t_L g1173 ( 
.A(n_1103),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1082),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1143),
.A2(n_1150),
.B(n_1148),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1083),
.B(n_1072),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1137),
.B(n_1095),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1048),
.B(n_1067),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1124),
.A2(n_1154),
.B(n_1049),
.C(n_1059),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1144),
.A2(n_1151),
.B(n_1158),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1163),
.B(n_1121),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1079),
.B(n_1086),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1080),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1147),
.A2(n_1157),
.B(n_1052),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1140),
.A2(n_1059),
.B1(n_1055),
.B2(n_1160),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1055),
.A2(n_1160),
.B1(n_1088),
.B2(n_1063),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_SL g1188 ( 
.A1(n_1062),
.A2(n_1091),
.B(n_1074),
.C(n_1102),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1071),
.A2(n_1100),
.B(n_1110),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1084),
.A2(n_1093),
.B(n_1126),
.Y(n_1190)
);

NOR2xp67_ASAP7_75t_L g1191 ( 
.A(n_1061),
.B(n_1043),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_1051),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1117),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1133),
.A2(n_1104),
.B(n_1081),
.Y(n_1194)
);

OAI211xp5_ASAP7_75t_L g1195 ( 
.A1(n_1111),
.A2(n_1139),
.B(n_1156),
.C(n_1153),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1145),
.Y(n_1196)
);

OR2x2_ASAP7_75t_L g1197 ( 
.A(n_1146),
.B(n_1138),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1088),
.A2(n_1096),
.B(n_1094),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_1077),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1054),
.Y(n_1200)
);

AOI222xp33_ASAP7_75t_L g1201 ( 
.A1(n_1076),
.A2(n_1078),
.B1(n_1098),
.B2(n_1107),
.C1(n_1161),
.C2(n_1159),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1056),
.A2(n_1155),
.B(n_1060),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1085),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1085),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1090),
.A2(n_1092),
.B1(n_1112),
.B2(n_1127),
.Y(n_1205)
);

INVx6_ASAP7_75t_L g1206 ( 
.A(n_1051),
.Y(n_1206)
);

AO21x2_ASAP7_75t_L g1207 ( 
.A1(n_1122),
.A2(n_1097),
.B(n_1070),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1111),
.A2(n_1116),
.B1(n_1105),
.B2(n_1106),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1082),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1082),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_SL g1211 ( 
.A1(n_1114),
.A2(n_1152),
.B(n_1149),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1069),
.A2(n_1070),
.B(n_1149),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1141),
.Y(n_1213)
);

AO21x2_ASAP7_75t_L g1214 ( 
.A1(n_1070),
.A2(n_1069),
.B(n_1152),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1113),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1125),
.A2(n_1149),
.B(n_1073),
.Y(n_1216)
);

INVx6_ASAP7_75t_L g1217 ( 
.A(n_1087),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1108),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1125),
.B(n_1119),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1099),
.Y(n_1220)
);

INVx6_ASAP7_75t_L g1221 ( 
.A(n_1101),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1069),
.A2(n_1101),
.B(n_1128),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1128),
.B(n_1142),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1065),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1047),
.A2(n_1130),
.B(n_1120),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1123),
.A2(n_1040),
.B(n_1031),
.C(n_1041),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1058),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1067),
.A2(n_676),
.B1(n_682),
.B2(n_663),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1057),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1047),
.A2(n_1130),
.B(n_1120),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1115),
.A2(n_847),
.B1(n_1131),
.B2(n_1109),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1047),
.A2(n_1130),
.B(n_1120),
.Y(n_1232)
);

CKINVDCx11_ASAP7_75t_R g1233 ( 
.A(n_1058),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1057),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1047),
.A2(n_1130),
.B(n_1120),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1137),
.B(n_1095),
.Y(n_1236)
);

OR2x6_ASAP7_75t_SL g1237 ( 
.A(n_1043),
.B(n_799),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1047),
.A2(n_1130),
.B(n_1120),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_1138),
.Y(n_1239)
);

AOI21xp33_ASAP7_75t_L g1240 ( 
.A1(n_1115),
.A2(n_851),
.B(n_853),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1082),
.Y(n_1241)
);

NOR2xp67_ASAP7_75t_L g1242 ( 
.A(n_1061),
.B(n_659),
.Y(n_1242)
);

AOI22x1_ASAP7_75t_L g1243 ( 
.A1(n_1086),
.A2(n_836),
.B1(n_711),
.B2(n_663),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1050),
.B(n_663),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1140),
.A2(n_847),
.B1(n_846),
.B2(n_417),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1057),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1140),
.A2(n_847),
.B1(n_846),
.B2(n_417),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1140),
.A2(n_847),
.B1(n_846),
.B2(n_417),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1137),
.B(n_1095),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1057),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1047),
.A2(n_1130),
.B(n_1120),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1086),
.B(n_1093),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1089),
.Y(n_1253)
);

CKINVDCx20_ASAP7_75t_R g1254 ( 
.A(n_1058),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1123),
.A2(n_851),
.B(n_1031),
.Y(n_1255)
);

NAND3xp33_ASAP7_75t_L g1256 ( 
.A(n_1123),
.B(n_851),
.C(n_1031),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1123),
.A2(n_851),
.B(n_1031),
.Y(n_1257)
);

OR2x2_ASAP7_75t_L g1258 ( 
.A(n_1068),
.B(n_1053),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1051),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1118),
.A2(n_1143),
.B(n_1129),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1050),
.B(n_663),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1126),
.A2(n_847),
.B1(n_1041),
.B2(n_927),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1064),
.A2(n_1045),
.B(n_1046),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_1233),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1197),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1239),
.Y(n_1266)
);

AOI21x1_ASAP7_75t_SL g1267 ( 
.A1(n_1219),
.A2(n_1178),
.B(n_1182),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1180),
.A2(n_1179),
.B1(n_1166),
.B2(n_1231),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1260),
.A2(n_1166),
.B(n_1165),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_SL g1270 ( 
.A1(n_1180),
.A2(n_1244),
.B1(n_1261),
.B2(n_1245),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1179),
.A2(n_1231),
.B1(n_1226),
.B2(n_1262),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1200),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1176),
.B(n_1167),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1255),
.A2(n_1257),
.B(n_1226),
.C(n_1256),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1262),
.A2(n_1261),
.B(n_1244),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1258),
.B(n_1195),
.Y(n_1276)
);

OAI31xp33_ASAP7_75t_L g1277 ( 
.A1(n_1240),
.A2(n_1228),
.A3(n_1195),
.B(n_1208),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1202),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1189),
.A2(n_1190),
.B(n_1243),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_R g1280 ( 
.A(n_1254),
.B(n_1168),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1172),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1196),
.B(n_1177),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1245),
.A2(n_1247),
.B1(n_1248),
.B2(n_1186),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1201),
.B(n_1177),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1236),
.B(n_1249),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1209),
.A2(n_1210),
.B(n_1185),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1183),
.A2(n_1198),
.B(n_1216),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1187),
.B(n_1186),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1247),
.A2(n_1248),
.B1(n_1205),
.B2(n_1252),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1172),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1196),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1224),
.Y(n_1292)
);

AOI221x1_ASAP7_75t_SL g1293 ( 
.A1(n_1184),
.A2(n_1234),
.B1(n_1250),
.B2(n_1229),
.C(n_1246),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1188),
.A2(n_1183),
.B(n_1164),
.C(n_1252),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1233),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1174),
.A2(n_1241),
.B1(n_1237),
.B2(n_1263),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1263),
.A2(n_1199),
.B1(n_1170),
.B2(n_1253),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1254),
.A2(n_1218),
.B1(n_1227),
.B2(n_1215),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1222),
.A2(n_1170),
.B(n_1253),
.C(n_1211),
.Y(n_1299)
);

OAI31xp33_ASAP7_75t_L g1300 ( 
.A1(n_1220),
.A2(n_1213),
.A3(n_1193),
.B(n_1223),
.Y(n_1300)
);

AOI221xp5_ASAP7_75t_L g1301 ( 
.A1(n_1214),
.A2(n_1224),
.B1(n_1207),
.B2(n_1204),
.C(n_1203),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1193),
.B(n_1213),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1214),
.B(n_1212),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1194),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1169),
.A2(n_1242),
.B1(n_1173),
.B2(n_1212),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1206),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1218),
.A2(n_1173),
.B1(n_1192),
.B2(n_1221),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1169),
.A2(n_1175),
.B(n_1191),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1171),
.B(n_1259),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1206),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1173),
.A2(n_1221),
.B1(n_1217),
.B2(n_1175),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1217),
.B(n_1181),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1217),
.A2(n_1225),
.B1(n_1230),
.B2(n_1232),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1235),
.B(n_1238),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1251),
.Y(n_1315)
);

O2A1O1Ixp5_ASAP7_75t_L g1316 ( 
.A1(n_1180),
.A2(n_1046),
.B(n_1164),
.C(n_1262),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1197),
.B(n_1239),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1180),
.A2(n_726),
.B1(n_727),
.B2(n_847),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1180),
.A2(n_1262),
.B1(n_847),
.B2(n_671),
.C(n_648),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1233),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1179),
.A2(n_1040),
.B(n_1031),
.Y(n_1321)
);

O2A1O1Ixp5_ASAP7_75t_L g1322 ( 
.A1(n_1180),
.A2(n_1046),
.B(n_1164),
.C(n_1262),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1172),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1259),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1180),
.B(n_434),
.Y(n_1325)
);

O2A1O1Ixp5_ASAP7_75t_L g1326 ( 
.A1(n_1180),
.A2(n_1046),
.B(n_1164),
.C(n_1262),
.Y(n_1326)
);

OAI221xp5_ASAP7_75t_L g1327 ( 
.A1(n_1180),
.A2(n_851),
.B1(n_1040),
.B2(n_1031),
.C(n_676),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1180),
.A2(n_726),
.B1(n_727),
.B2(n_847),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1312),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1269),
.B(n_1278),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1315),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1286),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1286),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1303),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1287),
.A2(n_1288),
.B(n_1289),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1319),
.A2(n_1328),
.B1(n_1318),
.B2(n_1268),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1279),
.B(n_1311),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1268),
.B(n_1274),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1288),
.A2(n_1289),
.B(n_1283),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1308),
.B(n_1321),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1315),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1279),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1304),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1314),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1272),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1313),
.A2(n_1305),
.B(n_1283),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1318),
.A2(n_1328),
.B1(n_1270),
.B2(n_1271),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1301),
.B(n_1296),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1297),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1271),
.B(n_1294),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1293),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1316),
.A2(n_1326),
.B(n_1322),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1276),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1266),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1327),
.A2(n_1275),
.B1(n_1325),
.B2(n_1284),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1277),
.B(n_1293),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1302),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1317),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1299),
.Y(n_1359)
);

CKINVDCx16_ASAP7_75t_R g1360 ( 
.A(n_1307),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1265),
.B(n_1273),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1353),
.B(n_1291),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1334),
.B(n_1310),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1343),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1341),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1331),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1337),
.B(n_1324),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1332),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1345),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1353),
.B(n_1300),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1343),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1344),
.B(n_1282),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_SL g1373 ( 
.A(n_1340),
.B(n_1323),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1333),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1353),
.B(n_1309),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1353),
.B(n_1323),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1344),
.B(n_1323),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1342),
.A2(n_1267),
.B(n_1285),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1357),
.B(n_1290),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1330),
.B(n_1290),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1369),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1363),
.B(n_1358),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1370),
.A2(n_1347),
.B1(n_1336),
.B2(n_1355),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1370),
.A2(n_1355),
.B(n_1347),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1368),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1380),
.A2(n_1339),
.B1(n_1336),
.B2(n_1335),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1364),
.Y(n_1387)
);

AND2x4_ASAP7_75t_SL g1388 ( 
.A(n_1372),
.B(n_1340),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1375),
.B(n_1358),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1378),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1364),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1369),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1369),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1373),
.B(n_1329),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1363),
.B(n_1358),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1376),
.Y(n_1396)
);

INVx5_ASAP7_75t_L g1397 ( 
.A(n_1371),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1362),
.B(n_1347),
.C(n_1355),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1371),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1380),
.B(n_1358),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1373),
.A2(n_1350),
.B1(n_1338),
.B2(n_1339),
.Y(n_1401)
);

NOR3xp33_ASAP7_75t_L g1402 ( 
.A(n_1362),
.B(n_1356),
.C(n_1338),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1380),
.B(n_1358),
.Y(n_1403)
);

OAI321xp33_ASAP7_75t_L g1404 ( 
.A1(n_1379),
.A2(n_1338),
.A3(n_1356),
.B1(n_1336),
.B2(n_1350),
.C(n_1346),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1373),
.A2(n_1350),
.B1(n_1339),
.B2(n_1335),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1378),
.A2(n_1339),
.B1(n_1335),
.B2(n_1350),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1363),
.Y(n_1407)
);

INVx4_ASAP7_75t_R g1408 ( 
.A(n_1366),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1367),
.B(n_1329),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1365),
.B(n_1329),
.Y(n_1410)
);

OAI31xp33_ASAP7_75t_L g1411 ( 
.A1(n_1375),
.A2(n_1350),
.A3(n_1356),
.B(n_1359),
.Y(n_1411)
);

CKINVDCx16_ASAP7_75t_R g1412 ( 
.A(n_1377),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1397),
.B(n_1367),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1381),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1381),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1392),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1392),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1402),
.Y(n_1418)
);

OR2x6_ASAP7_75t_L g1419 ( 
.A(n_1394),
.B(n_1340),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1393),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1393),
.Y(n_1421)
);

INVx4_ASAP7_75t_SL g1422 ( 
.A(n_1394),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1394),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1385),
.Y(n_1424)
);

INVxp67_ASAP7_75t_SL g1425 ( 
.A(n_1387),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1385),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1407),
.B(n_1374),
.Y(n_1427)
);

AOI21xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1383),
.A2(n_1360),
.B(n_1264),
.Y(n_1428)
);

INVx4_ASAP7_75t_SL g1429 ( 
.A(n_1394),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1397),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1391),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1397),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1397),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1399),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1424),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1431),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1424),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1430),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1422),
.B(n_1412),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1422),
.B(n_1412),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1422),
.B(n_1409),
.Y(n_1441)
);

AOI33xp33_ASAP7_75t_L g1442 ( 
.A1(n_1418),
.A2(n_1406),
.A3(n_1386),
.B1(n_1405),
.B2(n_1401),
.B3(n_1348),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1427),
.B(n_1407),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1418),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1427),
.B(n_1382),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1414),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1428),
.B(n_1411),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1427),
.B(n_1425),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1422),
.B(n_1409),
.Y(n_1449)
);

AND3x2_ASAP7_75t_L g1450 ( 
.A(n_1430),
.B(n_1411),
.C(n_1396),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1425),
.B(n_1382),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1431),
.B(n_1395),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1422),
.B(n_1400),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1422),
.B(n_1400),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1434),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1414),
.Y(n_1456)
);

NAND2x1_ASAP7_75t_L g1457 ( 
.A(n_1430),
.B(n_1408),
.Y(n_1457)
);

OR2x6_ASAP7_75t_L g1458 ( 
.A(n_1432),
.B(n_1340),
.Y(n_1458)
);

AOI21xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1428),
.A2(n_1320),
.B(n_1295),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1434),
.B(n_1403),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1432),
.B(n_1384),
.C(n_1398),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1415),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1429),
.B(n_1403),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1429),
.B(n_1388),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1424),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1416),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1416),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1417),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1429),
.B(n_1388),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1417),
.Y(n_1470)
);

NAND4xp25_ASAP7_75t_L g1471 ( 
.A(n_1423),
.B(n_1398),
.C(n_1359),
.D(n_1351),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1426),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1423),
.Y(n_1473)
);

AOI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1419),
.A2(n_1404),
.B(n_1335),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1429),
.B(n_1410),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1466),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1473),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1444),
.B(n_1461),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1446),
.Y(n_1479)
);

NOR4xp25_ASAP7_75t_L g1480 ( 
.A(n_1447),
.B(n_1404),
.C(n_1432),
.D(n_1433),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1446),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1439),
.B(n_1429),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1471),
.B(n_1361),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1473),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1456),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1448),
.B(n_1420),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1448),
.B(n_1420),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1439),
.B(n_1429),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1440),
.B(n_1464),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1440),
.B(n_1423),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1456),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1442),
.B(n_1361),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1450),
.B(n_1361),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1462),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1455),
.B(n_1421),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1469),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1474),
.B(n_1390),
.C(n_1352),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1436),
.B(n_1361),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1469),
.B(n_1419),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1462),
.Y(n_1500)
);

OAI21xp33_ASAP7_75t_L g1501 ( 
.A1(n_1460),
.A2(n_1348),
.B(n_1419),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1443),
.B(n_1389),
.Y(n_1502)
);

NOR3xp33_ASAP7_75t_L g1503 ( 
.A(n_1438),
.B(n_1298),
.C(n_1390),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1467),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1467),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1457),
.B(n_1432),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1441),
.B(n_1419),
.Y(n_1507)
);

AOI31xp33_ASAP7_75t_L g1508 ( 
.A1(n_1459),
.A2(n_1413),
.A3(n_1354),
.B(n_1359),
.Y(n_1508)
);

NAND2x1_ASAP7_75t_L g1509 ( 
.A(n_1438),
.B(n_1408),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1457),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1479),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1484),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1489),
.B(n_1441),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1490),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1481),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1480),
.A2(n_1437),
.B(n_1435),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1489),
.B(n_1482),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1485),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1482),
.B(n_1449),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1491),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1488),
.B(n_1449),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1478),
.B(n_1468),
.Y(n_1522)
);

INVxp67_ASAP7_75t_L g1523 ( 
.A(n_1484),
.Y(n_1523)
);

NAND2x1_ASAP7_75t_SL g1524 ( 
.A(n_1488),
.B(n_1438),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1477),
.B(n_1459),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1492),
.A2(n_1339),
.B1(n_1335),
.B2(n_1352),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1494),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1476),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1495),
.B(n_1443),
.Y(n_1530)
);

NAND2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1509),
.B(n_1432),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1490),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1508),
.B(n_1483),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1486),
.Y(n_1535)
);

OAI221xp5_ASAP7_75t_L g1536 ( 
.A1(n_1523),
.A2(n_1503),
.B1(n_1497),
.B2(n_1493),
.C(n_1510),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1523),
.B(n_1500),
.Y(n_1537)
);

NAND3xp33_ASAP7_75t_L g1538 ( 
.A(n_1529),
.B(n_1505),
.C(n_1504),
.Y(n_1538)
);

AOI32xp33_ASAP7_75t_L g1539 ( 
.A1(n_1534),
.A2(n_1501),
.A3(n_1507),
.B1(n_1499),
.B2(n_1510),
.Y(n_1539)
);

NAND2x1_ASAP7_75t_L g1540 ( 
.A(n_1513),
.B(n_1507),
.Y(n_1540)
);

AOI222xp33_ASAP7_75t_L g1541 ( 
.A1(n_1529),
.A2(n_1390),
.B1(n_1498),
.B2(n_1499),
.C1(n_1349),
.C2(n_1348),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1514),
.B(n_1532),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1524),
.A2(n_1433),
.B(n_1495),
.C(n_1451),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1512),
.B(n_1292),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1524),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1514),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1535),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1517),
.B(n_1486),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1517),
.B(n_1487),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1535),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1513),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1516),
.B(n_1487),
.Y(n_1552)
);

AO221x1_ASAP7_75t_L g1553 ( 
.A1(n_1514),
.A2(n_1433),
.B1(n_1470),
.B2(n_1468),
.C(n_1506),
.Y(n_1553)
);

OAI32xp33_ASAP7_75t_L g1554 ( 
.A1(n_1516),
.A2(n_1506),
.A3(n_1390),
.B1(n_1433),
.B2(n_1360),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1540),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1542),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1546),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1551),
.B(n_1512),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1545),
.B(n_1519),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1536),
.A2(n_1527),
.B1(n_1522),
.B2(n_1532),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1547),
.B(n_1516),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1550),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1548),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1544),
.B(n_1519),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1552),
.B(n_1516),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1544),
.Y(n_1566)
);

NOR4xp25_ASAP7_75t_L g1567 ( 
.A(n_1565),
.B(n_1561),
.C(n_1557),
.D(n_1558),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1565),
.A2(n_1554),
.B(n_1543),
.Y(n_1568)
);

NAND4xp25_ASAP7_75t_L g1569 ( 
.A(n_1559),
.B(n_1526),
.C(n_1512),
.D(n_1539),
.Y(n_1569)
);

AOI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1560),
.A2(n_1538),
.B1(n_1522),
.B2(n_1553),
.C(n_1537),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1560),
.A2(n_1549),
.B(n_1532),
.Y(n_1571)
);

NAND4xp25_ASAP7_75t_L g1572 ( 
.A(n_1564),
.B(n_1541),
.C(n_1521),
.D(n_1527),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1561),
.A2(n_1530),
.B(n_1531),
.Y(n_1573)
);

NOR3x1_ASAP7_75t_L g1574 ( 
.A(n_1555),
.B(n_1515),
.C(n_1511),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1563),
.A2(n_1521),
.B1(n_1533),
.B2(n_1525),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1567),
.A2(n_1556),
.B(n_1562),
.C(n_1566),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1575),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1569),
.A2(n_1531),
.B1(n_1530),
.B2(n_1360),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1570),
.A2(n_1520),
.B1(n_1511),
.B2(n_1515),
.C(n_1528),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1574),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1576),
.A2(n_1571),
.B(n_1568),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1577),
.B(n_1580),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1579),
.B(n_1525),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1578),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1580),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1577),
.B(n_1533),
.Y(n_1586)
);

NOR2xp67_ASAP7_75t_L g1587 ( 
.A(n_1585),
.B(n_1573),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1581),
.A2(n_1572),
.B1(n_1535),
.B2(n_1518),
.Y(n_1588)
);

O2A1O1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1581),
.A2(n_1528),
.B(n_1520),
.C(n_1518),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1584),
.B(n_1531),
.Y(n_1590)
);

AOI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1583),
.A2(n_1433),
.B1(n_1470),
.B2(n_1472),
.C(n_1435),
.Y(n_1591)
);

AOI211xp5_ASAP7_75t_L g1592 ( 
.A1(n_1590),
.A2(n_1586),
.B(n_1582),
.C(n_1280),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1587),
.B(n_1502),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1589),
.Y(n_1594)
);

AND3x4_ASAP7_75t_L g1595 ( 
.A(n_1592),
.B(n_1588),
.C(n_1591),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1595),
.Y(n_1596)
);

OAI22x1_ASAP7_75t_L g1597 ( 
.A1(n_1596),
.A2(n_1594),
.B1(n_1593),
.B2(n_1472),
.Y(n_1597)
);

XNOR2x1_ASAP7_75t_SL g1598 ( 
.A(n_1597),
.B(n_1453),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1598),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1599),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1599),
.B(n_1437),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1600),
.A2(n_1465),
.B1(n_1452),
.B2(n_1451),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1601),
.A2(n_1281),
.B(n_1458),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1603),
.B(n_1465),
.Y(n_1604)
);

NAND2xp33_ASAP7_75t_R g1605 ( 
.A(n_1602),
.B(n_1458),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1604),
.A2(n_1458),
.B1(n_1453),
.B2(n_1454),
.Y(n_1606)
);

AOI22x1_ASAP7_75t_L g1607 ( 
.A1(n_1605),
.A2(n_1360),
.B1(n_1452),
.B2(n_1463),
.Y(n_1607)
);

AOI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1606),
.A2(n_1463),
.B1(n_1454),
.B2(n_1458),
.Y(n_1608)
);

AOI211xp5_ASAP7_75t_L g1609 ( 
.A1(n_1608),
.A2(n_1607),
.B(n_1306),
.C(n_1445),
.Y(n_1609)
);


endmodule