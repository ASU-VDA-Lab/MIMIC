module fake_jpeg_23237_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_45),
.Y(n_57)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_28),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_19),
.B1(n_22),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_31),
.B1(n_34),
.B2(n_23),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_65),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_19),
.B1(n_18),
.B2(n_38),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_31),
.B1(n_27),
.B2(n_23),
.Y(n_110)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_29),
.Y(n_65)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_19),
.Y(n_88)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_28),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_89),
.B(n_91),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_45),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_43),
.B1(n_38),
.B2(n_46),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_92),
.A2(n_55),
.B1(n_35),
.B2(n_36),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_105),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_96),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_53),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_38),
.B1(n_49),
.B2(n_46),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_107),
.B1(n_110),
.B2(n_113),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_34),
.B1(n_31),
.B2(n_38),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_49),
.B1(n_30),
.B2(n_32),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_40),
.Y(n_115)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_51),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_51),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_55),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_63),
.B(n_40),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_51),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_77),
.B(n_27),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_24),
.B(n_17),
.C(n_21),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_154),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_131),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_24),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_130),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_40),
.B(n_35),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_114),
.C(n_111),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_21),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_95),
.A2(n_67),
.B1(n_80),
.B2(n_79),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_94),
.B(n_17),
.Y(n_138)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_146),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_151),
.B1(n_86),
.B2(n_101),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_28),
.B1(n_25),
.B2(n_36),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_152),
.B1(n_101),
.B2(n_86),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_25),
.Y(n_147)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_92),
.A2(n_39),
.B1(n_37),
.B2(n_28),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_110),
.A2(n_37),
.B1(n_82),
.B2(n_84),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_156),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_10),
.B(n_16),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_10),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_106),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_140),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_159),
.A2(n_164),
.B1(n_7),
.B2(n_14),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_90),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_174),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_169),
.B(n_184),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_0),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_114),
.C(n_99),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_176),
.C(n_188),
.Y(n_219)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_108),
.C(n_59),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_182),
.B1(n_187),
.B2(n_189),
.Y(n_192)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_96),
.B1(n_109),
.B2(n_104),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_96),
.B(n_109),
.C(n_76),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_125),
.A2(n_118),
.B1(n_97),
.B2(n_108),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_56),
.C(n_97),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_125),
.A2(n_106),
.B1(n_1),
.B2(n_2),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_106),
.A3(n_8),
.B1(n_9),
.B2(n_15),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_133),
.B(n_0),
.C(n_1),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_123),
.B1(n_145),
.B2(n_152),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_202),
.B1(n_220),
.B2(n_192),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_198),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_210),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_123),
.B1(n_129),
.B2(n_153),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_150),
.B(n_124),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_215),
.B(n_216),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_140),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_186),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_149),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_144),
.B1(n_126),
.B2(n_143),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

INVx5_ASAP7_75t_SL g214 ( 
.A(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_168),
.A2(n_131),
.B(n_138),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_170),
.A2(n_132),
.B(n_142),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_137),
.B1(n_8),
.B2(n_9),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_160),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_160),
.C(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_15),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_246),
.C(n_221),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_159),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_247),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_231),
.B(n_237),
.Y(n_249)
);

AO21x2_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_189),
.B(n_162),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_233),
.A2(n_239),
.B1(n_245),
.B2(n_196),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_166),
.B(n_162),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_236),
.B(n_210),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_175),
.B(n_183),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_205),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_205),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_242),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_161),
.B1(n_173),
.B2(n_2),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_0),
.Y(n_243)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_198),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_1),
.C(n_3),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_7),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_244),
.B(n_231),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_260),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_219),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_223),
.B(n_228),
.Y(n_273)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_257),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_225),
.C(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_199),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_224),
.A2(n_233),
.B1(n_241),
.B2(n_230),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_245),
.B1(n_201),
.B2(n_206),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_199),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_216),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_247),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_236),
.B(n_209),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_228),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_278),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_233),
.B1(n_244),
.B2(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_273),
.A2(n_249),
.B(n_248),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_279),
.C(n_256),
.Y(n_287)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_232),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_283),
.B1(n_229),
.B2(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_252),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_242),
.B1(n_215),
.B2(n_195),
.Y(n_283)
);

BUFx12f_ASAP7_75t_SL g286 ( 
.A(n_277),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_287),
.B(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_269),
.B(n_262),
.Y(n_291)
);

XOR2x1_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_298),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_251),
.C(n_254),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_294),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_258),
.C(n_263),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_296),
.A2(n_297),
.B1(n_284),
.B2(n_276),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_268),
.A2(n_275),
.B1(n_285),
.B2(n_283),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_252),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_259),
.C(n_200),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_299),
.B(n_270),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_304),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_288),
.A2(n_292),
.B1(n_271),
.B2(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_303),
.C(n_309),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_285),
.B1(n_281),
.B2(n_284),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_281),
.CI(n_278),
.CON(n_304),
.SN(n_304)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_274),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_SL g320 ( 
.A(n_310),
.B(n_317),
.C(n_304),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_309),
.A2(n_293),
.B1(n_291),
.B2(n_212),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.C(n_316),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_306),
.A2(n_294),
.B(n_208),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_207),
.B1(n_200),
.B2(n_3),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_307),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_314),
.Y(n_323)
);

AOI21xp33_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_304),
.B(n_303),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_320),
.B1(n_317),
.B2(n_11),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_313),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_324),
.A2(n_325),
.B(n_321),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_325),
.B(n_11),
.Y(n_328)
);

A2O1A1O1Ixp25_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_7),
.B(n_8),
.C(n_12),
.D(n_14),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_326),
.C(n_3),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_4),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_4),
.Y(n_332)
);


endmodule