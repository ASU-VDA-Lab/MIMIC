module real_jpeg_8445_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_1),
.A2(n_25),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_1),
.A2(n_38),
.B1(n_66),
.B2(n_67),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_1),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_3),
.A2(n_66),
.B1(n_67),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_90),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_90),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_3),
.A2(n_25),
.B1(n_35),
.B2(n_90),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g92 ( 
.A(n_4),
.Y(n_92)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_51),
.B(n_64),
.C(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_51),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_30),
.B(n_49),
.C(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_9),
.A2(n_51),
.B1(n_52),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_9),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_102),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_102),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_9),
.A2(n_25),
.B1(n_35),
.B2(n_102),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_10),
.A2(n_25),
.B1(n_35),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_10),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_10),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_59),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_59),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_11),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_150),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_150),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_11),
.A2(n_25),
.B1(n_35),
.B2(n_150),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_12),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_131),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_131),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_12),
.A2(n_25),
.B1(n_35),
.B2(n_131),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_13),
.A2(n_25),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_13),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_13),
.A2(n_34),
.B1(n_66),
.B2(n_67),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_15),
.A2(n_51),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_15),
.B(n_51),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_15),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_15),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_15),
.A2(n_30),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_15),
.B(n_30),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_15),
.B(n_32),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_15),
.A2(n_27),
.B(n_31),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_15),
.A2(n_25),
.B1(n_35),
.B2(n_115),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_16),
.A2(n_25),
.B1(n_35),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_16),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_16),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_61),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_17),
.A2(n_66),
.B1(n_67),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_17),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_17),
.A2(n_51),
.B1(n_52),
.B2(n_95),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_95),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_17),
.A2(n_25),
.B1(n_35),
.B2(n_95),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B(n_33),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_23),
.A2(n_32),
.B1(n_37),
.B2(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_23),
.A2(n_32),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_24),
.A2(n_29),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_24),
.A2(n_29),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_24),
.A2(n_29),
.B1(n_213),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_24),
.A2(n_29),
.B1(n_238),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_24),
.A2(n_29),
.B1(n_256),
.B2(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_24),
.A2(n_29),
.B1(n_58),
.B2(n_282),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_25),
.A2(n_26),
.B(n_115),
.C(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_36),
.B(n_43),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_77),
.B(n_334),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_70),
.C(n_72),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_44),
.A2(n_45),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_56),
.C(n_62),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_46),
.A2(n_47),
.B1(n_62),
.B2(n_309),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_48),
.A2(n_50),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_48),
.A2(n_50),
.B1(n_141),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_48),
.A2(n_50),
.B1(n_158),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_48),
.A2(n_50),
.B1(n_198),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_48),
.A2(n_50),
.B1(n_209),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_48),
.A2(n_50),
.B1(n_235),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_308),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_49),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_50),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_51),
.B(n_53),
.Y(n_145)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_52),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_56),
.A2(n_57),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_62),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_62),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_65),
.B(n_69),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_65),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_63),
.A2(n_65),
.B1(n_101),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_63),
.A2(n_65),
.B1(n_128),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_63),
.A2(n_65),
.B1(n_137),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_63),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_63),
.A2(n_65),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_63),
.A2(n_65),
.B1(n_221),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_63),
.A2(n_65),
.B1(n_230),
.B2(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_65),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_68),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_66),
.B(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_69),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_330),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_70),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_74),
.A2(n_75),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_327),
.B(n_333),
.Y(n_77)
);

OAI321xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_300),
.A3(n_320),
.B1(n_325),
.B2(n_326),
.C(n_336),
.Y(n_78)
);

AOI321xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_246),
.A3(n_288),
.B1(n_294),
.B2(n_299),
.C(n_337),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_203),
.C(n_242),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_173),
.B(n_202),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_152),
.B(n_172),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_133),
.B(n_151),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_122),
.B(n_132),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_108),
.B(n_121),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_96),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_96),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_91),
.A2(n_92),
.B1(n_149),
.B2(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_112),
.B1(n_113),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_103),
.B2(n_107),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_107),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_116),
.B(n_120),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_114),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_113),
.B1(n_130),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_112),
.A2(n_113),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_112),
.A2(n_113),
.B1(n_184),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_112),
.A2(n_113),
.B1(n_218),
.B2(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_112),
.A2(n_113),
.B(n_228),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_115),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_124),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_127),
.C(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_135),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_138),
.CI(n_142),
.CON(n_135),
.SN(n_135)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_140),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_147),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_165),
.B2(n_166),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_168),
.C(n_170),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_160),
.B2(n_164),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_162),
.C(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_167),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_168),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_174),
.B(n_175),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_188),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_177),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_177),
.B(n_187),
.C(n_188),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_182),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_199),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_196),
.B2(n_197),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_196),
.C(n_199),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_193),
.A2(n_195),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_201),
.Y(n_212)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_204),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_223),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_205),
.B(n_223),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_216),
.C(n_222),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_215),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_210),
.B1(n_211),
.B2(n_214),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_214),
.C(n_215),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_222),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_219),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_240),
.B2(n_241),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_226),
.B(n_231),
.C(n_241),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_229),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_236),
.C(n_239),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_234),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_240),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_243),
.B(n_244),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_265),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_247),
.B(n_265),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_258),
.C(n_264),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_248),
.A2(n_249),
.B1(n_258),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_254),
.C(n_257),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_252),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_253),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_258),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_260),
.B1(n_281),
.B2(n_283),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_259),
.A2(n_281),
.B(n_284),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_261),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_261),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_262),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_286),
.B2(n_287),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_277),
.B2(n_278),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_268),
.B(n_278),
.C(n_287),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_273),
.B(n_276),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_275),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_276),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_276),
.A2(n_302),
.B1(n_311),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_284),
.B2(n_285),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_281),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_289),
.A2(n_295),
.B(n_298),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_291),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_313),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_313),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_311),
.C(n_312),
.Y(n_301)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_302),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_304),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_309),
.C(n_310),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_315),
.C(n_319),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_307),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_332),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_329),
.Y(n_331)
);


endmodule