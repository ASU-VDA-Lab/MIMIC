module fake_jpeg_16215_n_80 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_80);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_7),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_31),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_34),
.C(n_16),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_13),
.B1(n_27),
.B2(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_57),
.Y(n_68)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_1),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_2),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_17),
.B1(n_24),
.B2(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B(n_4),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_3),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_67),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_65),
.Y(n_71)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_59),
.B1(n_11),
.B2(n_12),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_9),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_72),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_10),
.C(n_18),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_68),
.B(n_64),
.C(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_68),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_74),
.C(n_69),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_19),
.B(n_22),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);


endmodule