module fake_ariane_432_n_641 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_641);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_641;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_616;
wire n_617;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_544;
wire n_216;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_25),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_20),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_8),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_35),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_90),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_73),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_47),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_38),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_24),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_16),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_43),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_8),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_101),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_29),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_15),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_40),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_107),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_116),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_21),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_56),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_58),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_114),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_44),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_76),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_106),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_32),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_41),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_59),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_57),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_19),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_39),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_99),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_61),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_34),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_122),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_91),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_54),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_64),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_113),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_42),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_85),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_46),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_11),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_28),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_9),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_109),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_23),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_138),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_183),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_141),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_0),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_151),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_151),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_203),
.Y(n_224)
);

NOR2xp67_ASAP7_75t_L g225 ( 
.A(n_154),
.B(n_0),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_146),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_148),
.B(n_150),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_139),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_140),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_143),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_144),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_196),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_196),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_147),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_154),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_149),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

NAND2xp33_ASAP7_75t_R g244 ( 
.A(n_153),
.B(n_2),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_165),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_155),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_165),
.B(n_2),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_248),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_161),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_209),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_204),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_188),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_210),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_215),
.B(n_188),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_211),
.B(n_175),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_250),
.B(n_202),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_223),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_216),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_221),
.B(n_190),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_212),
.Y(n_290)
);

AND3x1_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_244),
.C(n_242),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

NAND2xp33_ASAP7_75t_SL g296 ( 
.A(n_237),
.B(n_177),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_206),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_224),
.A2(n_195),
.B1(n_200),
.B2(n_193),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_237),
.B(n_157),
.Y(n_301)
);

CKINVDCx8_ASAP7_75t_R g302 ( 
.A(n_242),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_259),
.B(n_158),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_262),
.Y(n_305)
);

AND3x4_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_244),
.C(n_4),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_301),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_160),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_162),
.Y(n_312)
);

AND3x4_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_3),
.C(n_4),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_252),
.B(n_177),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_163),
.Y(n_316)
);

INVx4_ASAP7_75t_SL g317 ( 
.A(n_292),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_252),
.B(n_177),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_292),
.B(n_166),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_264),
.B(n_177),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_13),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_253),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_3),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_192),
.B(n_191),
.Y(n_332)
);

AND2x6_ASAP7_75t_L g333 ( 
.A(n_295),
.B(n_14),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_167),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_17),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_R g340 ( 
.A(n_298),
.B(n_170),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_283),
.B(n_172),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_267),
.B(n_173),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_270),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_267),
.B(n_176),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_282),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_289),
.B(n_5),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_293),
.B(n_178),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_265),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_266),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_268),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_298),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_286),
.B(n_5),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_297),
.A2(n_186),
.B1(n_182),
.B2(n_181),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_280),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_272),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_278),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_284),
.Y(n_362)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_299),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_263),
.B(n_279),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_269),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_251),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_279),
.B(n_6),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_269),
.B(n_6),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_288),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_329),
.A2(n_349),
.B1(n_275),
.B2(n_296),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_305),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_311),
.Y(n_373)
);

AO22x2_ASAP7_75t_L g374 ( 
.A1(n_306),
.A2(n_275),
.B1(n_290),
.B2(n_302),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_309),
.B(n_251),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

AO22x2_ASAP7_75t_L g378 ( 
.A1(n_313),
.A2(n_287),
.B1(n_296),
.B2(n_300),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

OAI221xp5_ASAP7_75t_L g380 ( 
.A1(n_355),
.A2(n_258),
.B1(n_281),
.B2(n_273),
.C(n_11),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_366),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_303),
.B(n_258),
.Y(n_382)
);

AO22x2_ASAP7_75t_L g383 ( 
.A1(n_329),
.A2(n_281),
.B1(n_273),
.B2(n_276),
.Y(n_383)
);

AO22x2_ASAP7_75t_L g384 ( 
.A1(n_349),
.A2(n_276),
.B1(n_9),
.B2(n_10),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_7),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_317),
.B(n_7),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_354),
.Y(n_389)
);

OAI221xp5_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_10),
.B1(n_12),
.B2(n_18),
.C(n_22),
.Y(n_390)
);

OAI221xp5_ASAP7_75t_L g391 ( 
.A1(n_364),
.A2(n_12),
.B1(n_26),
.B2(n_27),
.C(n_30),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_137),
.Y(n_394)
);

AO22x2_ASAP7_75t_L g395 ( 
.A1(n_368),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_134),
.Y(n_396)
);

AO22x2_ASAP7_75t_L g397 ( 
.A1(n_368),
.A2(n_37),
.B1(n_45),
.B2(n_48),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_308),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_331),
.B(n_49),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_50),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_308),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_337),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_351),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_307),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_411)
);

AO22x2_ASAP7_75t_L g412 ( 
.A1(n_365),
.A2(n_55),
.B1(n_60),
.B2(n_63),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_348),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_360),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_351),
.B(n_131),
.Y(n_416)
);

AO22x2_ASAP7_75t_L g417 ( 
.A1(n_324),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_363),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_321),
.B(n_69),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_314),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_314),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_318),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_310),
.B(n_71),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_312),
.B(n_129),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_319),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_304),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_304),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_L g429 ( 
.A(n_316),
.B(n_72),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_318),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_376),
.B(n_363),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_350),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_382),
.B(n_332),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_SL g434 ( 
.A(n_419),
.B(n_347),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_373),
.B(n_304),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_373),
.B(n_345),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_388),
.B(n_345),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_388),
.B(n_386),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_385),
.B(n_343),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_370),
.B(n_344),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_369),
.B(n_345),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_369),
.B(n_334),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_SL g443 ( 
.A(n_379),
.B(n_322),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_SL g444 ( 
.A(n_387),
.B(n_334),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_420),
.B(n_401),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_420),
.B(n_401),
.Y(n_446)
);

NAND2xp33_ASAP7_75t_SL g447 ( 
.A(n_392),
.B(n_389),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_400),
.B(n_334),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_372),
.B(n_356),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_393),
.B(n_326),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_326),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_408),
.B(n_328),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_409),
.B(n_338),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_371),
.B(n_330),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_410),
.B(n_325),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_413),
.B(n_315),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_339),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_426),
.B(n_339),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_374),
.B(n_333),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_381),
.B(n_333),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_398),
.B(n_333),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_381),
.B(n_333),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_375),
.B(n_327),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_377),
.B(n_327),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_415),
.B(n_327),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_421),
.B(n_327),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_422),
.B(n_74),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_423),
.B(n_75),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_399),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_394),
.B(n_402),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_469),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_463),
.A2(n_396),
.B(n_416),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_418),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_433),
.A2(n_403),
.B(n_404),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_405),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_455),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_446),
.B(n_414),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_432),
.A2(n_380),
.B(n_411),
.C(n_390),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_428),
.Y(n_479)
);

OAI22x1_ASAP7_75t_L g480 ( 
.A1(n_459),
.A2(n_378),
.B1(n_384),
.B2(n_374),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_464),
.A2(n_425),
.B(n_427),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_456),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_470),
.A2(n_429),
.B(n_395),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_457),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_451),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_457),
.A2(n_397),
.B1(n_412),
.B2(n_378),
.Y(n_487)
);

AOI221x1_ASAP7_75t_L g488 ( 
.A1(n_439),
.A2(n_412),
.B1(n_417),
.B2(n_384),
.C(n_383),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_447),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_457),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_454),
.B(n_417),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_466),
.A2(n_391),
.B(n_78),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_443),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g494 ( 
.A1(n_461),
.A2(n_77),
.B(n_79),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_435),
.B(n_80),
.Y(n_495)
);

A2O1A1Ixp33_ASAP7_75t_L g496 ( 
.A1(n_452),
.A2(n_81),
.B(n_82),
.C(n_83),
.Y(n_496)
);

INVx3_ASAP7_75t_SL g497 ( 
.A(n_460),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_450),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_126),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_431),
.Y(n_500)
);

OA21x2_ASAP7_75t_L g501 ( 
.A1(n_483),
.A2(n_465),
.B(n_458),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_481),
.A2(n_472),
.B(n_494),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_473),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_468),
.B(n_467),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_436),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_474),
.A2(n_453),
.B(n_442),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_482),
.Y(n_507)
);

AOI222xp33_ASAP7_75t_L g508 ( 
.A1(n_487),
.A2(n_434),
.B1(n_448),
.B2(n_441),
.C1(n_444),
.C2(n_92),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_473),
.B(n_125),
.Y(n_509)
);

OAI22xp33_ASAP7_75t_L g510 ( 
.A1(n_488),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_489),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_479),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_495),
.A2(n_95),
.B(n_97),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_497),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_475),
.A2(n_98),
.B(n_100),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_477),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_477),
.Y(n_518)
);

OR2x6_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_102),
.Y(n_519)
);

INVx8_ASAP7_75t_L g520 ( 
.A(n_499),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_475),
.A2(n_103),
.B(n_105),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_108),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_489),
.B(n_111),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_478),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_486),
.Y(n_525)
);

CKINVDCx11_ASAP7_75t_R g526 ( 
.A(n_515),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_517),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_519),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_518),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_506),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_520),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_524),
.A2(n_493),
.B(n_496),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_520),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_501),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_511),
.B(n_491),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_511),
.B(n_490),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_513),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_498),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_502),
.A2(n_476),
.B(n_485),
.Y(n_539)
);

AO21x2_ASAP7_75t_L g540 ( 
.A1(n_510),
.A2(n_492),
.B(n_484),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_484),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_492),
.Y(n_542)
);

OAI221xp5_ASAP7_75t_L g543 ( 
.A1(n_522),
.A2(n_508),
.B1(n_524),
.B2(n_500),
.C(n_512),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_501),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_522),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g546 ( 
.A(n_520),
.B(n_505),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_525),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_123),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_507),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_508),
.A2(n_124),
.B(n_504),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_509),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_523),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_516),
.A2(n_521),
.B(n_514),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_525),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_525),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_520),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_531),
.B(n_526),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_537),
.Y(n_558)
);

XOR2x2_ASAP7_75t_SL g559 ( 
.A(n_552),
.B(n_551),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_535),
.B(n_536),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_526),
.Y(n_561)
);

CKINVDCx8_ASAP7_75t_R g562 ( 
.A(n_531),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_533),
.B(n_546),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_533),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_R g565 ( 
.A(n_545),
.B(n_538),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_545),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_R g567 ( 
.A(n_538),
.B(n_541),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_535),
.B(n_536),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_528),
.B(n_538),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_R g570 ( 
.A(n_541),
.B(n_542),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_537),
.Y(n_571)
);

OR2x4_ASAP7_75t_L g572 ( 
.A(n_528),
.B(n_548),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_556),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_R g574 ( 
.A(n_542),
.B(n_546),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_547),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_546),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_549),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_527),
.B(n_529),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_575),
.B(n_527),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_542),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_566),
.B(n_578),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_579),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_544),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_571),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_579),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_544),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_557),
.Y(n_588)
);

NOR2x1p5_ASAP7_75t_L g589 ( 
.A(n_561),
.B(n_528),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_568),
.B(n_530),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_558),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_563),
.B(n_569),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_564),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_559),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_577),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_593),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_534),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_594),
.A2(n_543),
.B1(n_550),
.B2(n_565),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_584),
.B(n_580),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_590),
.B(n_529),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_587),
.Y(n_601)
);

AO21x2_ASAP7_75t_L g602 ( 
.A1(n_585),
.A2(n_555),
.B(n_554),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_602),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_597),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_601),
.B(n_587),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_599),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_600),
.B(n_591),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_601),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_596),
.B(n_588),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_605),
.B(n_595),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_608),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_607),
.B(n_598),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_606),
.B(n_594),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_604),
.B(n_583),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_612),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_611),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_610),
.Y(n_617)
);

AOI21xp33_ASAP7_75t_L g618 ( 
.A1(n_613),
.A2(n_603),
.B(n_609),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_614),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_615),
.B(n_608),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_616),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_617),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g623 ( 
.A(n_621),
.B(n_618),
.C(n_619),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_622),
.B(n_617),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_624),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_625),
.B(n_623),
.C(n_620),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_626),
.A2(n_532),
.B(n_572),
.Y(n_627)
);

NOR2x1_ASAP7_75t_L g628 ( 
.A(n_627),
.B(n_589),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_R g629 ( 
.A(n_628),
.B(n_562),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_629),
.B(n_573),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_630),
.B(n_592),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_631),
.B(n_587),
.C(n_592),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_632),
.A2(n_540),
.B1(n_576),
.B2(n_539),
.Y(n_633)
);

NAND4xp25_ASAP7_75t_L g634 ( 
.A(n_633),
.B(n_567),
.C(n_592),
.D(n_570),
.Y(n_634)
);

OAI322xp33_ASAP7_75t_L g635 ( 
.A1(n_633),
.A2(n_530),
.A3(n_574),
.B1(n_586),
.B2(n_583),
.C1(n_534),
.C2(n_539),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_634),
.B(n_581),
.Y(n_636)
);

INVxp67_ASAP7_75t_L g637 ( 
.A(n_635),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_637),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_636),
.Y(n_639)
);

AOI221xp5_ASAP7_75t_L g640 ( 
.A1(n_638),
.A2(n_530),
.B1(n_540),
.B2(n_581),
.C(n_534),
.Y(n_640)
);

AOI211xp5_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_639),
.B(n_553),
.C(n_581),
.Y(n_641)
);


endmodule