module fake_jpeg_15575_n_121 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_8),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_21),
.B1(n_19),
.B2(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_38),
.B1(n_23),
.B2(n_26),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_5),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_23),
.A2(n_20),
.B1(n_22),
.B2(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_48),
.B1(n_53),
.B2(n_61),
.Y(n_64)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_49),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_25),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_52),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_25),
.Y(n_52)
);

AND2x6_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_4),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_29),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_28),
.A2(n_22),
.B1(n_21),
.B2(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_41),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_60),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_38),
.B1(n_28),
.B2(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_71),
.B1(n_59),
.B2(n_50),
.Y(n_89)
);

OAI22x1_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_28),
.B1(n_36),
.B2(n_30),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_52),
.B(n_44),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_79),
.B(n_60),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_36),
.C(n_5),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_48),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_78),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_73),
.B(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_61),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_40),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_42),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_53),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_90),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_88),
.B(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_47),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_64),
.B1(n_74),
.B2(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_64),
.B1(n_69),
.B2(n_79),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_103),
.B1(n_90),
.B2(n_89),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_79),
.B(n_77),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_77),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_93),
.C(n_67),
.Y(n_111)
);

AO221x1_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_70),
.B1(n_63),
.B2(n_43),
.C(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_70),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_SL g106 ( 
.A(n_94),
.B(n_84),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_108),
.B1(n_98),
.B2(n_102),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_87),
.B(n_86),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_109),
.B(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_97),
.A3(n_98),
.B1(n_103),
.B2(n_95),
.C1(n_101),
.C2(n_96),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_115),
.A3(n_116),
.B1(n_112),
.B2(n_111),
.C1(n_105),
.C2(n_9),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_118),
.A2(n_119),
.B(n_116),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

OAI321xp33_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_6),
.A3(n_13),
.B1(n_117),
.B2(n_106),
.C(n_108),
.Y(n_121)
);


endmodule