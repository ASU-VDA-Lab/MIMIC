module real_aes_628_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g465 ( .A(n_0), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_1), .B(n_261), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_2), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g138 ( .A(n_3), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_4), .B(n_507), .Y(n_539) );
NAND2xp33_ASAP7_75t_SL g533 ( .A(n_5), .B(n_150), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_6), .B(n_157), .Y(n_253) );
INVx1_ASAP7_75t_L g526 ( .A(n_7), .Y(n_526) );
INVx1_ASAP7_75t_L g166 ( .A(n_8), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_9), .Y(n_794) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_10), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_11), .Y(n_183) );
AND2x2_ASAP7_75t_L g537 ( .A(n_12), .B(n_210), .Y(n_537) );
INVx2_ASAP7_75t_L g127 ( .A(n_13), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_14), .Y(n_108) );
INVx1_ASAP7_75t_L g262 ( .A(n_15), .Y(n_262) );
AOI221x1_ASAP7_75t_L g529 ( .A1(n_16), .A2(n_124), .B1(n_506), .B2(n_530), .C(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_17), .B(n_507), .Y(n_515) );
INVx1_ASAP7_75t_L g112 ( .A(n_18), .Y(n_112) );
INVx1_ASAP7_75t_L g259 ( .A(n_19), .Y(n_259) );
INVx1_ASAP7_75t_SL g224 ( .A(n_20), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_21), .B(n_144), .Y(n_245) );
AOI33xp33_ASAP7_75t_L g195 ( .A1(n_22), .A2(n_52), .A3(n_133), .B1(n_142), .B2(n_196), .B3(n_197), .Y(n_195) );
AOI221xp5_ASAP7_75t_SL g505 ( .A1(n_23), .A2(n_41), .B1(n_506), .B2(n_507), .C(n_508), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_24), .A2(n_506), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_25), .B(n_261), .Y(n_542) );
INVx1_ASAP7_75t_L g175 ( .A(n_26), .Y(n_175) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_27), .A2(n_90), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g158 ( .A(n_27), .B(n_90), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_28), .B(n_264), .Y(n_519) );
INVxp67_ASAP7_75t_L g528 ( .A(n_29), .Y(n_528) );
AND2x2_ASAP7_75t_L g573 ( .A(n_30), .B(n_209), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_31), .B(n_152), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_32), .A2(n_506), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_33), .B(n_264), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_34), .A2(n_44), .B1(n_784), .B2(n_785), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_34), .Y(n_784) );
INVx1_ASAP7_75t_L g132 ( .A(n_35), .Y(n_132) );
AND2x2_ASAP7_75t_L g150 ( .A(n_35), .B(n_138), .Y(n_150) );
AND2x2_ASAP7_75t_L g156 ( .A(n_35), .B(n_135), .Y(n_156) );
OR2x6_ASAP7_75t_L g110 ( .A(n_36), .B(n_111), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_37), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_38), .B(n_152), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_39), .A2(n_125), .B1(n_157), .B2(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_40), .B(n_247), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_42), .A2(n_81), .B1(n_130), .B2(n_506), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_43), .B(n_144), .Y(n_225) );
INVx1_ASAP7_75t_L g785 ( .A(n_44), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_45), .B(n_261), .Y(n_571) );
AOI222xp33_ASAP7_75t_L g101 ( .A1(n_46), .A2(n_102), .B1(n_467), .B2(n_472), .C1(n_481), .C2(n_797), .Y(n_101) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_46), .A2(n_115), .B1(n_463), .B2(n_464), .Y(n_114) );
INVx1_ASAP7_75t_L g463 ( .A(n_46), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_47), .B(n_163), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_48), .B(n_144), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_49), .Y(n_242) );
AND2x2_ASAP7_75t_L g587 ( .A(n_50), .B(n_209), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_51), .B(n_209), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_53), .B(n_144), .Y(n_207) );
INVx1_ASAP7_75t_L g137 ( .A(n_54), .Y(n_137) );
INVx1_ASAP7_75t_L g146 ( .A(n_54), .Y(n_146) );
AND2x2_ASAP7_75t_L g208 ( .A(n_55), .B(n_209), .Y(n_208) );
AOI221xp5_ASAP7_75t_L g164 ( .A1(n_56), .A2(n_74), .B1(n_130), .B2(n_152), .C(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_57), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_58), .B(n_507), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_59), .B(n_125), .Y(n_185) );
AOI21xp5_ASAP7_75t_SL g129 ( .A1(n_60), .A2(n_130), .B(n_139), .Y(n_129) );
AND2x2_ASAP7_75t_L g552 ( .A(n_61), .B(n_209), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_62), .B(n_264), .Y(n_585) );
INVx1_ASAP7_75t_L g256 ( .A(n_63), .Y(n_256) );
AND2x2_ASAP7_75t_SL g520 ( .A(n_64), .B(n_210), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_65), .B(n_261), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_66), .A2(n_506), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g206 ( .A(n_67), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_68), .B(n_264), .Y(n_543) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_69), .B(n_163), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g460 ( .A1(n_70), .A2(n_89), .B1(n_461), .B2(n_462), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_70), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_71), .A2(n_130), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g135 ( .A(n_72), .Y(n_135) );
INVx1_ASAP7_75t_L g148 ( .A(n_72), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_73), .B(n_152), .Y(n_198) );
AND2x2_ASAP7_75t_L g226 ( .A(n_75), .B(n_124), .Y(n_226) );
INVx1_ASAP7_75t_L g257 ( .A(n_76), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_77), .A2(n_130), .B(n_223), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_78), .A2(n_130), .B(n_190), .C(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_79), .B(n_507), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_80), .A2(n_84), .B1(n_152), .B2(n_507), .Y(n_556) );
INVx1_ASAP7_75t_L g113 ( .A(n_82), .Y(n_113) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_83), .B(n_124), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_85), .A2(n_130), .B1(n_193), .B2(n_194), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_86), .B(n_261), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_87), .B(n_261), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_88), .A2(n_506), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g462 ( .A(n_89), .Y(n_462) );
NOR2xp33_ASAP7_75t_SL g486 ( .A(n_89), .B(n_487), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_89), .A2(n_490), .B(n_491), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_89), .A2(n_487), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_92), .B(n_264), .Y(n_549) );
AND2x2_ASAP7_75t_L g199 ( .A(n_93), .B(n_124), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_94), .A2(n_173), .B(n_174), .C(n_177), .Y(n_172) );
INVxp67_ASAP7_75t_L g531 ( .A(n_95), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_96), .B(n_507), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_97), .B(n_264), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_98), .A2(n_506), .B(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g471 ( .A(n_99), .Y(n_471) );
BUFx2_ASAP7_75t_SL g478 ( .A(n_99), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_100), .B(n_144), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_114), .B(n_465), .Y(n_102) );
CKINVDCx11_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g466 ( .A(n_106), .Y(n_466) );
AND2x2_ASAP7_75t_L g799 ( .A(n_106), .B(n_800), .Y(n_799) );
BUFx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g480 ( .A(n_107), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x6_ASAP7_75t_SL g497 ( .A(n_108), .B(n_110), .Y(n_497) );
OR2x6_ASAP7_75t_SL g782 ( .A(n_108), .B(n_109), .Y(n_782) );
OR2x2_ASAP7_75t_L g796 ( .A(n_108), .B(n_110), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVx2_ASAP7_75t_L g464 ( .A(n_115), .Y(n_464) );
XOR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_459), .Y(n_115) );
NAND3x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_349), .C(n_414), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_303), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_248), .B(n_276), .Y(n_118) );
AOI21xp33_ASAP7_75t_SL g488 ( .A1(n_119), .A2(n_248), .B(n_276), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_211), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_159), .Y(n_120) );
AOI21xp33_ASAP7_75t_L g350 ( .A1(n_121), .A2(n_351), .B(n_362), .Y(n_350) );
AND2x2_ASAP7_75t_SL g385 ( .A(n_121), .B(n_292), .Y(n_385) );
AND2x2_ASAP7_75t_L g400 ( .A(n_121), .B(n_401), .Y(n_400) );
OR2x6_ASAP7_75t_L g410 ( .A(n_121), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g412 ( .A(n_121), .B(n_402), .Y(n_412) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g286 ( .A(n_122), .Y(n_286) );
AND2x2_ASAP7_75t_L g299 ( .A(n_122), .B(n_300), .Y(n_299) );
INVx4_ASAP7_75t_L g318 ( .A(n_122), .Y(n_318) );
AND2x2_ASAP7_75t_L g321 ( .A(n_122), .B(n_237), .Y(n_321) );
NOR2x1_ASAP7_75t_SL g324 ( .A(n_122), .B(n_252), .Y(n_324) );
AND2x4_ASAP7_75t_L g336 ( .A(n_122), .B(n_334), .Y(n_336) );
OR2x2_ASAP7_75t_L g346 ( .A(n_122), .B(n_218), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_122), .B(n_358), .Y(n_363) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_128), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_124), .A2(n_172), .B1(n_178), .B2(n_179), .Y(n_171) );
INVx3_ASAP7_75t_L g179 ( .A(n_124), .Y(n_179) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_125), .B(n_182), .Y(n_181) );
AOI21x1_ASAP7_75t_L g580 ( .A1(n_125), .A2(n_581), .B(n_587), .Y(n_580) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
AND2x4_ASAP7_75t_L g157 ( .A(n_127), .B(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_127), .B(n_158), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_151), .B(n_157), .Y(n_128) );
INVxp67_ASAP7_75t_L g184 ( .A(n_130), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_130), .A2(n_152), .B1(n_525), .B2(n_527), .Y(n_524) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
NOR2x1p5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g197 ( .A(n_133), .Y(n_197) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x6_ASAP7_75t_L g141 ( .A(n_134), .B(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x6_ASAP7_75t_L g261 ( .A(n_135), .B(n_145), .Y(n_261) );
AND2x6_ASAP7_75t_L g506 ( .A(n_136), .B(n_156), .Y(n_506) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
INVx2_ASAP7_75t_L g142 ( .A(n_137), .Y(n_142) );
AND2x4_ASAP7_75t_L g264 ( .A(n_137), .B(n_147), .Y(n_264) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_141), .B(n_143), .C(n_149), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_SL g165 ( .A1(n_141), .A2(n_149), .B(n_166), .C(n_167), .Y(n_165) );
INVxp67_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_141), .A2(n_149), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_141), .A2(n_149), .B(n_224), .C(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g247 ( .A(n_141), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_141), .A2(n_176), .B1(n_256), .B2(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g153 ( .A(n_142), .B(n_154), .Y(n_153) );
INVxp33_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
INVx1_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
AND2x4_ASAP7_75t_L g507 ( .A(n_144), .B(n_150), .Y(n_507) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g193 ( .A(n_149), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_149), .A2(n_245), .B(n_246), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_149), .B(n_157), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_149), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_149), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_149), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_149), .A2(n_549), .B(n_550), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_149), .A2(n_570), .B(n_571), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_149), .A2(n_584), .B(n_585), .Y(n_583) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_150), .Y(n_177) );
INVx1_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx1_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_155), .Y(n_241) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_157), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_157), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_157), .B(n_531), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g532 ( .A(n_157), .B(n_176), .C(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_157), .A2(n_539), .B(n_540), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_159), .A2(n_292), .B1(n_387), .B2(n_388), .Y(n_386) );
INVx1_ASAP7_75t_SL g430 ( .A(n_159), .Y(n_430) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_187), .Y(n_159) );
INVx2_ASAP7_75t_L g361 ( .A(n_160), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_160), .B(n_307), .Y(n_433) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_169), .Y(n_160) );
BUFx3_ASAP7_75t_L g279 ( .A(n_161), .Y(n_279) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g272 ( .A(n_162), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_162), .B(n_189), .Y(n_294) );
AND2x4_ASAP7_75t_L g311 ( .A(n_162), .B(n_312), .Y(n_311) );
INVxp67_ASAP7_75t_L g327 ( .A(n_162), .Y(n_327) );
INVx2_ASAP7_75t_L g384 ( .A(n_162), .Y(n_384) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_168), .Y(n_162) );
INVx2_ASAP7_75t_SL g190 ( .A(n_163), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_163), .A2(n_515), .B(n_516), .Y(n_514) );
AND2x2_ASAP7_75t_L g302 ( .A(n_169), .B(n_268), .Y(n_302) );
NOR2xp67_ASAP7_75t_L g348 ( .A(n_169), .B(n_271), .Y(n_348) );
AND2x2_ASAP7_75t_L g367 ( .A(n_169), .B(n_271), .Y(n_367) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g229 ( .A(n_170), .Y(n_229) );
INVx1_ASAP7_75t_L g310 ( .A(n_170), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_170), .B(n_201), .Y(n_329) );
AND2x4_ASAP7_75t_L g383 ( .A(n_170), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_180), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_179), .A2(n_202), .B(n_208), .Y(n_201) );
AO21x2_ASAP7_75t_L g271 ( .A1(n_179), .A2(n_202), .B(n_208), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g342 ( .A(n_187), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_187), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g187 ( .A(n_188), .B(n_200), .Y(n_187) );
AND2x2_ASAP7_75t_L g326 ( .A(n_188), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g366 ( .A(n_188), .Y(n_366) );
AND2x2_ASAP7_75t_L g371 ( .A(n_188), .B(n_271), .Y(n_371) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_189), .B(n_201), .Y(n_231) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_199), .Y(n_189) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_190), .A2(n_191), .B(n_199), .Y(n_268) );
AOI21x1_ASAP7_75t_L g554 ( .A1(n_190), .A2(n_555), .B(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_192), .B(n_198), .Y(n_191) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g307 ( .A(n_200), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_200), .B(n_279), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_200), .B(n_229), .Y(n_446) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_201), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_209), .Y(n_219) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_209), .A2(n_505), .B(n_511), .Y(n_504) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OAI21xp33_ASAP7_75t_SL g211 ( .A1(n_212), .A2(n_227), .B(n_232), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_214), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g284 ( .A(n_215), .Y(n_284) );
AND2x2_ASAP7_75t_L g298 ( .A(n_215), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g332 ( .A(n_215), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g398 ( .A(n_215), .B(n_316), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g444 ( .A(n_215), .B(n_445), .C(n_446), .Y(n_444) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_216), .Y(n_275) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g291 ( .A(n_218), .Y(n_291) );
AND2x2_ASAP7_75t_L g297 ( .A(n_218), .B(n_252), .Y(n_297) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_218), .Y(n_308) );
AND2x2_ASAP7_75t_L g353 ( .A(n_218), .B(n_251), .Y(n_353) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_218), .Y(n_376) );
INVx1_ASAP7_75t_L g393 ( .A(n_218), .Y(n_393) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_226), .Y(n_218) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_219), .A2(n_546), .B(n_552), .Y(n_545) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_219), .A2(n_567), .B(n_573), .Y(n_566) );
AO21x2_ASAP7_75t_L g630 ( .A1(n_219), .A2(n_567), .B(n_573), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g435 ( .A(n_227), .Y(n_435) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_228), .B(n_306), .Y(n_407) );
INVx1_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g269 ( .A(n_229), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AOI211x1_ASAP7_75t_L g303 ( .A1(n_233), .A2(n_304), .B(n_313), .C(n_330), .Y(n_303) );
INVx2_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_SL g296 ( .A(n_234), .B(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g356 ( .A(n_234), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g292 ( .A(n_236), .B(n_251), .Y(n_292) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x4_ASAP7_75t_L g250 ( .A(n_237), .B(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_237), .Y(n_317) );
INVx1_ASAP7_75t_L g334 ( .A(n_237), .Y(n_334) );
AND2x2_ASAP7_75t_L g402 ( .A(n_237), .B(n_252), .Y(n_402) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_243), .Y(n_237) );
NOR3xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .C(n_242), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_266), .B(n_273), .Y(n_248) );
NOR2x1_ASAP7_75t_L g421 ( .A(n_249), .B(n_318), .Y(n_421) );
INVx2_ASAP7_75t_L g453 ( .A(n_249), .Y(n_453) );
INVx4_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g285 ( .A(n_250), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g358 ( .A(n_251), .Y(n_358) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g300 ( .A(n_252), .Y(n_300) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_258), .B(n_265), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B1(n_262), .B2(n_263), .Y(n_258) );
INVxp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVxp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
OR2x2_ASAP7_75t_L g360 ( .A(n_267), .B(n_361), .Y(n_360) );
NAND2x1_ASAP7_75t_SL g382 ( .A(n_267), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x4_ASAP7_75t_L g282 ( .A(n_268), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
INVx1_ASAP7_75t_L g436 ( .A(n_269), .Y(n_436) );
AND2x2_ASAP7_75t_L g301 ( .A(n_270), .B(n_302), .Y(n_301) );
NOR2x1_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g283 ( .A(n_271), .Y(n_283) );
INVxp33_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g340 ( .A(n_275), .B(n_333), .Y(n_340) );
OAI211xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_287), .C(n_295), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g364 ( .A(n_278), .B(n_365), .Y(n_364) );
NOR2xp67_ASAP7_75t_SL g369 ( .A(n_278), .B(n_370), .Y(n_369) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_279), .B(n_366), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_281), .B(n_285), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
AND2x2_ASAP7_75t_L g413 ( .A(n_282), .B(n_383), .Y(n_413) );
AOI222xp33_ASAP7_75t_L g431 ( .A1(n_285), .A2(n_432), .B1(n_434), .B2(n_437), .C1(n_438), .C2(n_441), .Y(n_431) );
INVx1_ASAP7_75t_L g395 ( .A(n_286), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_293), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_291), .Y(n_322) );
AND2x4_ASAP7_75t_SL g357 ( .A(n_291), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g411 ( .A(n_292), .Y(n_411) );
AND2x2_ASAP7_75t_L g456 ( .A(n_292), .B(n_308), .Y(n_456) );
AND2x2_ASAP7_75t_L g337 ( .A(n_293), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g450 ( .A(n_294), .B(n_329), .Y(n_450) );
OAI21xp33_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_298), .B(n_301), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_296), .A2(n_316), .B(n_357), .Y(n_417) );
AND2x2_ASAP7_75t_L g441 ( .A(n_297), .B(n_318), .Y(n_441) );
NOR2xp33_ASAP7_75t_SL g451 ( .A(n_297), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g389 ( .A(n_300), .Y(n_389) );
NOR2x1_ASAP7_75t_L g394 ( .A(n_300), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g424 ( .A(n_302), .Y(n_424) );
INVx1_ASAP7_75t_L g487 ( .A(n_303), .Y(n_487) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_309), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g427 ( .A(n_307), .B(n_311), .Y(n_427) );
BUFx2_ASAP7_75t_L g315 ( .A(n_308), .Y(n_315) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g338 ( .A(n_310), .Y(n_338) );
INVx2_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
AND2x2_ASAP7_75t_L g380 ( .A(n_310), .B(n_371), .Y(n_380) );
AND2x4_ASAP7_75t_L g347 ( .A(n_311), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g387 ( .A(n_311), .B(n_344), .Y(n_387) );
AND2x2_ASAP7_75t_L g438 ( .A(n_311), .B(n_439), .Y(n_438) );
AOI31xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_319), .A3(n_323), .B(n_325), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g335 ( .A(n_315), .B(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_SL g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x4_ASAP7_75t_L g333 ( .A(n_318), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_321), .A2(n_373), .B1(n_404), .B2(n_407), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_321), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g458 ( .A(n_321), .B(n_374), .Y(n_458) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g373 ( .A(n_324), .B(n_374), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g396 ( .A(n_326), .B(n_367), .Y(n_396) );
INVx1_ASAP7_75t_L g406 ( .A(n_328), .Y(n_406) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_339), .Y(n_330) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B(n_337), .Y(n_331) );
INVx1_ASAP7_75t_L g429 ( .A(n_332), .Y(n_429) );
AND2x2_ASAP7_75t_L g437 ( .A(n_333), .B(n_389), .Y(n_437) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_333), .Y(n_443) );
AND2x2_ASAP7_75t_L g388 ( .A(n_336), .B(n_389), .Y(n_388) );
AOI22xp33_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_341), .B1(n_345), .B2(n_347), .Y(n_339) );
NOR2xp33_ASAP7_75t_SL g341 ( .A(n_342), .B(n_343), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_342), .A2(n_361), .B1(n_455), .B2(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g354 ( .A(n_347), .Y(n_354) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_349), .B(n_414), .C(n_486), .D(n_488), .Y(n_485) );
INVxp67_ASAP7_75t_L g490 ( .A(n_349), .Y(n_490) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_377), .Y(n_349) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_354), .B(n_355), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
OAI21xp33_ASAP7_75t_L g355 ( .A1(n_353), .A2(n_356), .B(n_359), .Y(n_355) );
AOI22xp33_ASAP7_75t_SL g379 ( .A1(n_356), .A2(n_380), .B1(n_381), .B2(n_385), .Y(n_379) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_368), .B2(n_372), .Y(n_362) );
INVx1_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2xp67_ASAP7_75t_L g377 ( .A(n_378), .B(n_390), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_386), .Y(n_378) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
NAND2xp33_ASAP7_75t_SL g432 ( .A(n_382), .B(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g405 ( .A(n_383), .Y(n_405) );
INVx3_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
INVxp67_ASAP7_75t_L g448 ( .A(n_388), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_391), .B(n_399), .C(n_403), .D(n_408), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_396), .B1(n_397), .B2(n_398), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g401 ( .A(n_393), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g449 ( .A(n_397), .Y(n_449) );
NAND2xp33_ASAP7_75t_SL g404 ( .A(n_405), .B(n_406), .Y(n_404) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B(n_413), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g493 ( .A(n_414), .Y(n_493) );
AND3x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_431), .C(n_442), .Y(n_414) );
AOI221x1_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B1(n_420), .B2(n_422), .C(n_428), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp33_ASAP7_75t_SL g422 ( .A(n_423), .B(n_426), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
NAND2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI211xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_447), .C(n_454), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_447) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_SL g468 ( .A(n_469), .B(n_471), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_469), .A2(n_476), .B(n_479), .Y(n_475) );
INVx2_ASAP7_75t_L g802 ( .A(n_469), .Y(n_802) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_471), .B(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
CKINVDCx11_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
CKINVDCx8_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_783), .B(n_786), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_484), .A2(n_494), .B1(n_498), .B2(n_780), .Y(n_483) );
INVx1_ASAP7_75t_L g788 ( .A(n_484), .Y(n_788) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_489), .C(n_492), .Y(n_484) );
INVx1_ASAP7_75t_L g491 ( .A(n_488), .Y(n_491) );
OAI21x1_ASAP7_75t_L g787 ( .A1(n_494), .A2(n_788), .B(n_789), .Y(n_787) );
CKINVDCx6p67_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
INVx3_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
NAND2x1_ASAP7_75t_SL g789 ( .A(n_498), .B(n_790), .Y(n_789) );
INVx4_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_693), .Y(n_499) );
NAND3xp33_ASAP7_75t_SL g500 ( .A(n_501), .B(n_603), .C(n_643), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_521), .B(n_534), .C(n_559), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_502), .B(n_608), .Y(n_642) );
NOR2x1p5_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
INVx2_ASAP7_75t_L g594 ( .A(n_504), .Y(n_594) );
OR2x2_ASAP7_75t_L g606 ( .A(n_504), .B(n_513), .Y(n_606) );
AND2x2_ASAP7_75t_L g620 ( .A(n_504), .B(n_579), .Y(n_620) );
INVx1_ASAP7_75t_L g648 ( .A(n_504), .Y(n_648) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_504), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_504), .B(n_513), .Y(n_754) );
OR2x2_ASAP7_75t_L g575 ( .A(n_512), .B(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_512), .Y(n_710) );
AND2x2_ASAP7_75t_L g715 ( .A(n_512), .B(n_577), .Y(n_715) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g521 ( .A(n_513), .B(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g574 ( .A(n_513), .B(n_523), .Y(n_574) );
OR2x2_ASAP7_75t_L g593 ( .A(n_513), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g622 ( .A(n_513), .Y(n_622) );
AND2x4_ASAP7_75t_SL g661 ( .A(n_513), .B(n_523), .Y(n_661) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_513), .Y(n_665) );
OR2x2_ASAP7_75t_L g682 ( .A(n_513), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g692 ( .A(n_513), .B(n_599), .Y(n_692) );
INVx1_ASAP7_75t_L g721 ( .A(n_513), .Y(n_721) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_520), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_521), .B(n_650), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_522), .B(n_579), .Y(n_596) );
AND2x2_ASAP7_75t_L g608 ( .A(n_522), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g626 ( .A(n_522), .B(n_593), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_522), .B(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g599 ( .A(n_523), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g621 ( .A(n_523), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g656 ( .A(n_523), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_523), .B(n_579), .Y(n_680) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .Y(n_523) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_535), .B(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g629 ( .A(n_535), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_535), .B(n_545), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_535), .B(n_650), .C(n_651), .Y(n_649) );
AND2x2_ASAP7_75t_L g697 ( .A(n_535), .B(n_602), .Y(n_697) );
INVx5_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g564 ( .A(n_536), .B(n_565), .Y(n_564) );
AND2x4_ASAP7_75t_SL g601 ( .A(n_536), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g617 ( .A(n_536), .Y(n_617) );
OR2x2_ASAP7_75t_L g640 ( .A(n_536), .B(n_630), .Y(n_640) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_536), .Y(n_657) );
AND2x2_ASAP7_75t_SL g675 ( .A(n_536), .B(n_563), .Y(n_675) );
AND2x4_ASAP7_75t_L g690 ( .A(n_536), .B(n_566), .Y(n_690) );
AND2x2_ASAP7_75t_L g704 ( .A(n_536), .B(n_545), .Y(n_704) );
OR2x2_ASAP7_75t_L g725 ( .A(n_536), .B(n_553), .Y(n_725) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g779 ( .A(n_544), .B(n_657), .Y(n_779) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .Y(n_544) );
AND2x4_ASAP7_75t_L g602 ( .A(n_545), .B(n_565), .Y(n_602) );
INVx2_ASAP7_75t_L g613 ( .A(n_545), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_545), .B(n_563), .Y(n_618) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_545), .Y(n_651) );
OR2x2_ASAP7_75t_L g674 ( .A(n_545), .B(n_566), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_545), .B(n_566), .Y(n_677) );
INVx1_ASAP7_75t_L g686 ( .A(n_545), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
AND2x2_ASAP7_75t_L g589 ( .A(n_553), .B(n_566), .Y(n_589) );
BUFx2_ASAP7_75t_L g638 ( .A(n_553), .Y(n_638) );
AND2x2_ASAP7_75t_L g733 ( .A(n_553), .B(n_613), .Y(n_733) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_554), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_574), .B1(n_575), .B2(n_588), .C(n_590), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_562), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_562), .B(n_629), .Y(n_669) );
OR2x2_ASAP7_75t_L g681 ( .A(n_562), .B(n_677), .Y(n_681) );
OR2x2_ASAP7_75t_L g684 ( .A(n_562), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g773 ( .A(n_562), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g612 ( .A(n_563), .B(n_613), .Y(n_612) );
OA33x2_ASAP7_75t_L g645 ( .A1(n_563), .A2(n_606), .A3(n_646), .B1(n_649), .B2(n_652), .B3(n_655), .Y(n_645) );
OR2x2_ASAP7_75t_L g676 ( .A(n_563), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g700 ( .A(n_563), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g708 ( .A(n_563), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g728 ( .A(n_563), .B(n_602), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_563), .B(n_617), .Y(n_766) );
INVx2_ASAP7_75t_L g636 ( .A(n_564), .Y(n_636) );
AOI322xp5_ASAP7_75t_L g706 ( .A1(n_564), .A2(n_619), .A3(n_707), .B1(n_710), .B2(n_711), .C1(n_713), .C2(n_715), .Y(n_706) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_566), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
OR2x2_ASAP7_75t_L g688 ( .A(n_574), .B(n_667), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_574), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g761 ( .A(n_574), .Y(n_761) );
INVx1_ASAP7_75t_SL g627 ( .A(n_575), .Y(n_627) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g660 ( .A(n_577), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx2_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
INVx1_ASAP7_75t_L g609 ( .A(n_579), .Y(n_609) );
INVx1_ASAP7_75t_L g650 ( .A(n_579), .Y(n_650) );
OR2x2_ASAP7_75t_L g667 ( .A(n_579), .B(n_594), .Y(n_667) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_579), .Y(n_742) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .Y(n_581) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_589), .B(n_712), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_597), .B(n_601), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_591), .A2(n_665), .B(n_666), .C(n_668), .Y(n_664) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g729 ( .A(n_593), .B(n_730), .Y(n_729) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_594), .Y(n_598) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g753 ( .A(n_596), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_SL g722 ( .A(n_599), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g730 ( .A(n_599), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_599), .B(n_721), .Y(n_738) );
INVx3_ASAP7_75t_SL g663 ( .A(n_602), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_610), .B1(n_614), .B2(n_619), .C(n_623), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_609), .Y(n_654) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_612), .A2(n_639), .B(n_711), .Y(n_717) );
AND2x2_ASAP7_75t_L g743 ( .A(n_612), .B(n_690), .Y(n_743) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_613), .Y(n_631) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_617), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g752 ( .A(n_617), .B(n_674), .Y(n_752) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g701 ( .A(n_620), .Y(n_701) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_628), .B(n_632), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx2_ASAP7_75t_L g774 ( .A(n_629), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_630), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g703 ( .A(n_630), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_631), .B(n_653), .Y(n_652) );
OAI31xp33_ASAP7_75t_SL g632 ( .A1(n_633), .A2(n_635), .A3(n_637), .B(n_641), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_636), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OR2x2_ASAP7_75t_L g714 ( .A(n_638), .B(n_640), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_638), .B(n_690), .Y(n_769) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NOR5xp2_ASAP7_75t_L g643 ( .A(n_644), .B(n_658), .C(n_670), .D(n_679), .E(n_687), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_648), .B(n_650), .Y(n_683) );
INVx1_ASAP7_75t_L g723 ( .A(n_648), .Y(n_723) );
INVxp67_ASAP7_75t_SL g760 ( .A(n_648), .Y(n_760) );
INVx1_ASAP7_75t_L g712 ( .A(n_651), .Y(n_712) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp33_ASAP7_75t_SL g655 ( .A(n_656), .B(n_657), .Y(n_655) );
OAI321xp33_ASAP7_75t_L g695 ( .A1(n_656), .A2(n_696), .A3(n_698), .B1(n_702), .B2(n_705), .C(n_706), .Y(n_695) );
INVx1_ASAP7_75t_L g749 ( .A(n_657), .Y(n_749) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B(n_664), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_660), .A2(n_733), .B1(n_740), .B2(n_743), .Y(n_739) );
AND2x2_ASAP7_75t_L g768 ( .A(n_661), .B(n_742), .Y(n_768) );
INVx1_ASAP7_75t_L g678 ( .A(n_666), .Y(n_678) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_676), .B(n_678), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_677), .A2(n_688), .B1(n_689), .B2(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g750 ( .A(n_677), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B1(n_682), .B2(n_684), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_686), .B(n_690), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_688), .A2(n_765), .B1(n_767), .B2(n_769), .C(n_770), .Y(n_764) );
INVx1_ASAP7_75t_L g771 ( .A(n_688), .Y(n_771) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_689), .A2(n_746), .B1(n_753), .B2(n_755), .C(n_756), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g716 ( .A1(n_691), .A2(n_717), .B(n_718), .Y(n_716) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_744), .Y(n_693) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_716), .C(n_734), .Y(n_694) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_697), .Y(n_763) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g762 ( .A(n_705), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_707), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g755 ( .A(n_715), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_724), .B(n_726), .Y(n_718) );
INVxp67_ASAP7_75t_L g776 ( .A(n_719), .Y(n_776) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_SL g731 ( .A(n_722), .Y(n_731) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_729), .B1(n_731), .B2(n_732), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B(n_739), .Y(n_734) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g777 ( .A(n_740), .Y(n_777) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_764), .C(n_775), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_751), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI21xp5_ASAP7_75t_SL g756 ( .A1(n_757), .A2(n_762), .B(n_763), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVxp67_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_768), .A2(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AOI21xp33_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B(n_778), .Y(n_775) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_781), .Y(n_792) );
CKINVDCx11_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_783), .A2(n_787), .B(n_793), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
BUFx4f_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
BUFx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVxp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
endmodule