module fake_jpeg_3522_n_113 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_113);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_113;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_30),
.A2(n_26),
.B1(n_27),
.B2(n_11),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_3),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_40),
.Y(n_48)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_7),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_49),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_39),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_30),
.A2(n_27),
.B1(n_23),
.B2(n_21),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_56),
.B1(n_19),
.B2(n_11),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_8),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_61),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_57),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_65),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_31),
.C(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_10),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_69),
.Y(n_81)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_10),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_51),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp67_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_82),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_45),
.Y(n_80)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_63),
.C(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_71),
.B1(n_79),
.B2(n_76),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_96),
.B1(n_87),
.B2(n_65),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_77),
.B(n_71),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_97),
.Y(n_101)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_78),
.A3(n_76),
.B1(n_80),
.B2(n_75),
.C(n_61),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_75),
.B(n_61),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_100),
.B(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_94),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_103),
.C(n_45),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_84),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_64),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_105),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_101),
.B(n_55),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_102),
.B(n_100),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_51),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_107),
.B(n_55),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_68),
.C(n_54),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_19),
.Y(n_113)
);


endmodule