module fake_jpeg_3930_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_5),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_0),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_17),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_18),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_3),
.Y(n_18)
);

AO22x2_ASAP7_75t_L g19 ( 
.A1(n_11),
.A2(n_3),
.B1(n_4),
.B2(n_13),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_12),
.B(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_SL g33 ( 
.A1(n_32),
.A2(n_19),
.B(n_22),
.C(n_7),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_SL g37 ( 
.A1(n_33),
.A2(n_19),
.B(n_9),
.C(n_17),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_23),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_29),
.A3(n_27),
.B1(n_18),
.B2(n_24),
.C1(n_26),
.C2(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_37),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_33),
.B(n_35),
.Y(n_39)
);


endmodule