module real_jpeg_1570_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_1),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_1),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_1),
.B(n_32),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_1),
.B(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_68),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_1),
.Y(n_150)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_2),
.B(n_39),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_2),
.B(n_70),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_46),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_2),
.B(n_42),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_2),
.B(n_68),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_3),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_3),
.B(n_42),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_3),
.B(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_3),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_3),
.B(n_68),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_35),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_5),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_5),
.B(n_42),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_5),
.B(n_27),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_68),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_5),
.B(n_32),
.Y(n_265)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_6),
.B(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_6),
.B(n_46),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_70),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_10),
.B(n_27),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_10),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_10),
.B(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_10),
.B(n_42),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_46),
.Y(n_153)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_12),
.B(n_39),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_12),
.B(n_70),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_12),
.B(n_46),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_12),
.B(n_42),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_14),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_14),
.B(n_46),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_14),
.B(n_42),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_14),
.B(n_68),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_14),
.B(n_27),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_14),
.B(n_32),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_169),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_167),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_19),
.B(n_133),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_81),
.C(n_114),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_20),
.A2(n_21),
.B1(n_114),
.B2(n_115),
.Y(n_173)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_58),
.B2(n_80),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_22),
.B(n_59),
.C(n_73),
.Y(n_134)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.C(n_47),
.Y(n_23)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_24),
.B(n_37),
.CI(n_47),
.CON(n_199),
.SN(n_199)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_26),
.B(n_31),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_26),
.A2(n_33),
.B1(n_185),
.B2(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_28),
.B(n_63),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_30),
.A2(n_31),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_30),
.A2(n_33),
.B(n_34),
.C(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_30),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_30),
.A2(n_31),
.B1(n_253),
.B2(n_254),
.Y(n_266)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_31),
.B(n_118),
.C(n_120),
.Y(n_162)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_32),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_33),
.B(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.C(n_45),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_38),
.A2(n_45),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_38),
.Y(n_197)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_41),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_41),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_41),
.A2(n_154),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_45),
.Y(n_196)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_46),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_53),
.C(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_50),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_55),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_55),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_67),
.C(n_69),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_60),
.A2(n_61),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.C(n_66),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_65),
.A2(n_66),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_66),
.A2(n_87),
.B1(n_118),
.B2(n_119),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_69),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_67),
.Y(n_112)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_74),
.B(n_77),
.C(n_78),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_77),
.A2(n_79),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_81),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_99),
.C(n_109),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_82),
.A2(n_83),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.C(n_92),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_84),
.B(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_89),
.A2(n_90),
.B(n_91),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_92),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.C(n_97),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_95),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_99),
.B(n_109),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_107),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_100),
.B(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.C(n_104),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_101),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_102),
.B(n_186),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_102),
.B(n_106),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_103),
.A2(n_104),
.B1(n_128),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_128),
.B1(n_129),
.B2(n_132),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_130),
.C(n_131),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_105),
.B(n_107),
.Y(n_191)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_124),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_125),
.C(n_127),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_119),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_126),
.A2(n_208),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_157),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_145),
.B2(n_156),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_188),
.C(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_143),
.A2(n_144),
.B1(n_188),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_153),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_157),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.CI(n_160),
.CON(n_157),
.SN(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_200),
.B(n_321),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_172),
.B(n_174),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_198),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_175),
.A2(n_198),
.B1(n_199),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_175),
.Y(n_316)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_178),
.B(n_315),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_190),
.C(n_192),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_187),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_181),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_188),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_190),
.A2(n_192),
.B1(n_193),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_199),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_318),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_312),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_237),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_229),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_205),
.B(n_229),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_215),
.C(n_219),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_206),
.B(n_309),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_206),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_211),
.CI(n_212),
.CON(n_206),
.SN(n_206)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_211),
.C(n_212),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.C(n_210),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_209),
.B(n_210),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_215),
.B(n_219),
.Y(n_309)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.C(n_227),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_220),
.B(n_223),
.CI(n_227),
.CON(n_299),
.SN(n_299)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.C(n_226),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_226),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_248),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_229),
.Y(n_329)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.CI(n_234),
.CON(n_229),
.SN(n_229)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_230),
.B(n_233),
.C(n_234),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_307),
.B(n_311),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_295),
.B(n_306),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_267),
.B(n_294),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_258),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_258),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_251),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_243),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.C(n_246),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_245),
.CI(n_246),
.CON(n_259),
.SN(n_259)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_247),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_249),
.C(n_251),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_256),
.C(n_257),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.C(n_266),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_291),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_259),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_261),
.B1(n_266),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_288),
.B(n_293),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_279),
.B(n_287),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_275),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_275),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_273),
.C(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_282),
.B(n_286),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_302),
.C(n_303),
.Y(n_310)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_299),
.Y(n_328)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_310),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_313),
.A2(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);


endmodule