module fake_jpeg_14566_n_82 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_82);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_82;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx5_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_9),
.A2(n_7),
.B(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_1),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_17),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_20),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_10),
.B1(n_21),
.B2(n_25),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_26),
.B1(n_15),
.B2(n_17),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_49),
.C(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_5),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_31),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_16),
.B(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_18),
.B1(n_28),
.B2(n_16),
.Y(n_50)
);

A2O1A1O1Ixp25_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_28),
.B(n_18),
.C(n_9),
.D(n_8),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_28),
.B(n_5),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_41),
.B(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_40),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_46),
.C(n_50),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_59),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_55),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_71),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_32),
.B1(n_39),
.B2(n_42),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_63),
.C(n_62),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_71),
.C(n_67),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_59),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

AOI321xp33_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_76),
.A3(n_78),
.B1(n_8),
.B2(n_32),
.C(n_39),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_32),
.Y(n_82)
);


endmodule