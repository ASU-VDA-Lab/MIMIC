module fake_netlist_1_519_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
NAND2xp5_ASAP7_75t_SL g3 ( .A(n_0), .B(n_1), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
INVx8_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
HB1xp67_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
OAI21xp5_ASAP7_75t_L g7 ( .A1(n_4), .A2(n_2), .B(n_0), .Y(n_7) );
AOI21x1_ASAP7_75t_L g8 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_6), .B(n_5), .Y(n_10) );
OR2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_7), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_9), .B(n_7), .Y(n_12) );
AOI221xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_2), .C(n_11), .Y(n_13) );
NAND3xp33_ASAP7_75t_SL g14 ( .A(n_13), .B(n_1), .C(n_6), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
OR2x2_ASAP7_75t_L g16 ( .A(n_15), .B(n_1), .Y(n_16) );
endmodule