module fake_jpeg_19096_n_181 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_25),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_29),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g30 ( 
.A(n_17),
.B(n_10),
.CON(n_30),
.SN(n_30)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_11),
.B1(n_18),
.B2(n_15),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_31),
.B(n_27),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_20),
.B1(n_12),
.B2(n_15),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_22),
.B1(n_20),
.B2(n_12),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_49),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_25),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_20),
.B(n_14),
.C(n_24),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_50),
.B(n_45),
.Y(n_65)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_13),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_23),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_54),
.B1(n_40),
.B2(n_50),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_26),
.B1(n_12),
.B2(n_35),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_61),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_65),
.B(n_62),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

OA21x2_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_48),
.B(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_73),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_57),
.B(n_62),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_41),
.B1(n_50),
.B2(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_75),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_56),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_82),
.C(n_90),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_86),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_46),
.B(n_52),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_94),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_40),
.B1(n_57),
.B2(n_61),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_89),
.B1(n_93),
.B2(n_50),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_57),
.B1(n_63),
.B2(n_53),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_63),
.C(n_68),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_50),
.B(n_49),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_43),
.C(n_44),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_42),
.B(n_43),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_97),
.B(n_64),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_108),
.B1(n_111),
.B2(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_86),
.C(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_107),
.C(n_110),
.Y(n_120)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_80),
.Y(n_117)
);

XOR2x1_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_70),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_78),
.C(n_70),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_79),
.B1(n_76),
.B2(n_50),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_44),
.C(n_67),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_69),
.B1(n_67),
.B2(n_43),
.Y(n_111)
);

NAND2xp67_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_81),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_19),
.C(n_7),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_121),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_98),
.B1(n_99),
.B2(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_51),
.B1(n_64),
.B2(n_55),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_127),
.B1(n_108),
.B2(n_47),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_16),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_51),
.B1(n_64),
.B2(n_55),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_33),
.C(n_35),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_120),
.C(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_140),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_96),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_136),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_96),
.B(n_110),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_9),
.B(n_8),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_140),
.C(n_118),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_125),
.B1(n_122),
.B2(n_14),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_19),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_19),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_141),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_33),
.C(n_47),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_16),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_149),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_144),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_124),
.C(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_132),
.B1(n_138),
.B2(n_141),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_10),
.B1(n_9),
.B2(n_8),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_150),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_21),
.C(n_14),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_21),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_154),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_139),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_157),
.B(n_0),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_136),
.B(n_9),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_0),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_0),
.B(n_1),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_148),
.C(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_162),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_158),
.B(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_153),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_161),
.B(n_2),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_164),
.B(n_165),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_21),
.C(n_1),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_166),
.B(n_1),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_171),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_170),
.B(n_172),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_21),
.C(n_3),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_160),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_175),
.B(n_174),
.Y(n_177)
);

AOI21x1_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_3),
.B(n_4),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_3),
.B(n_5),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_177),
.A2(n_5),
.B(n_6),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_178),
.B(n_5),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);


endmodule