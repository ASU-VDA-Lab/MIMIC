module real_jpeg_15207_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_98),
.B1(n_101),
.B2(n_106),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_0),
.A2(n_106),
.B1(n_144),
.B2(n_149),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_0),
.A2(n_106),
.B1(n_261),
.B2(n_264),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_0),
.A2(n_106),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_509),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_1),
.B(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_2),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_4),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_5),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_5),
.A2(n_180),
.B1(n_226),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_5),
.A2(n_180),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_5),
.A2(n_180),
.B1(n_325),
.B2(n_328),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_7),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_7),
.A2(n_55),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_7),
.A2(n_55),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_7),
.A2(n_299),
.A3(n_302),
.B1(n_305),
.B2(n_309),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_7),
.B(n_42),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_7),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_7),
.B(n_57),
.Y(n_363)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_8),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_8),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_8),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_9),
.A2(n_25),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_9),
.A2(n_25),
.B1(n_336),
.B2(n_339),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

BUFx4f_ASAP7_75t_L g200 ( 
.A(n_12),
.Y(n_200)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_13),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_168),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_166),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_156),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_18),
.B(n_156),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.C(n_140),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_19),
.A2(n_132),
.B1(n_155),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_19),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_88),
.B1(n_89),
.B2(n_131),
.Y(n_19)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_20),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_56),
.B2(n_87),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_22),
.B(n_56),
.C(n_88),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

AND2x4_ASAP7_75t_SL g291 ( 
.A(n_23),
.B(n_292),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_23),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_24),
.B(n_42),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_25),
.B(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_29),
.Y(n_148)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_30),
.Y(n_281)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_33),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_33),
.B(n_177),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_42),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_38),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_38),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_40),
.Y(n_222)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_42),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_42),
.B(n_177),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_42),
.A2(n_468),
.B(n_469),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_45),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AND2x4_ASAP7_75t_SL g401 ( 
.A(n_49),
.B(n_176),
.Y(n_401)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_50),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_53),
.A2(n_219),
.A3(n_223),
.B1(n_228),
.B2(n_232),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_55),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_55),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_R g216 ( 
.A(n_55),
.B(n_90),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_55),
.B(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_55),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_R g141 ( 
.A(n_56),
.B(n_142),
.C(n_155),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_56),
.A2(n_87),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_56),
.A2(n_87),
.B1(n_142),
.B2(n_495),
.Y(n_494)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_68),
.B(n_80),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_57),
.B(n_80),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_57),
.B(n_250),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_57),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_57),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_66),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_61),
.Y(n_264)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_61),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_70),
.B1(n_73),
.B2(n_76),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_68),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_68),
.B(n_80),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_68),
.B(n_335),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_68),
.Y(n_447)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_72),
.Y(n_338)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_72),
.Y(n_342)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_79),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_86),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_87),
.B(n_283),
.C(n_291),
.Y(n_431)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_97),
.B(n_107),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_90),
.A2(n_159),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_90),
.A2(n_159),
.B(n_454),
.Y(n_475)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_90)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_91),
.Y(n_271)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_95),
.Y(n_179)
);

OAI21x1_ASAP7_75t_R g158 ( 
.A1(n_97),
.A2(n_133),
.B(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_100),
.Y(n_288)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_108),
.B(n_284),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_126),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_109),
.B(n_285),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_115),
.B1(n_119),
.B2(n_123),
.Y(n_110)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_114),
.Y(n_276)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g286 ( 
.A(n_130),
.Y(n_286)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_132),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_133),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_134),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_135),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_136),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_138),
.A2(n_269),
.B1(n_272),
.B2(n_281),
.Y(n_268)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_141),
.B(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_142),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_153),
.B(n_154),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_143),
.Y(n_468)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

AOI21x1_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g383 ( 
.A(n_153),
.B(n_162),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_154),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_158),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_160),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_160),
.A2(n_164),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_164),
.B(n_419),
.C(n_425),
.Y(n_441)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_488),
.B(n_506),
.Y(n_169)
);

AO221x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_395),
.B1(n_481),
.B2(n_486),
.C(n_487),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_293),
.B(n_394),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_253),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_173),
.B(n_253),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_217),
.C(n_245),
.Y(n_173)
);

XOR2x1_ASAP7_75t_L g389 ( 
.A(n_174),
.B(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_183),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_175),
.B(n_184),
.C(n_216),
.Y(n_256)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_215),
.B2(n_216),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_205),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_186),
.B(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_196),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_187),
.B(n_209),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_187),
.B(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_187),
.A2(n_260),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_191),
.Y(n_304)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_192),
.Y(n_322)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_195),
.Y(n_360)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_199),
.Y(n_308)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_203),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_204),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_205),
.B(n_323),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_205),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_209),
.B(n_211),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_217),
.A2(n_245),
.B1(n_246),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_217),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_238),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_218),
.A2(n_238),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_218),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_226),
.Y(n_301)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_238),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_238),
.A2(n_385),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_238),
.A2(n_385),
.B1(n_475),
.B2(n_476),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_238),
.B(n_445),
.Y(n_477)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_243),
.B(n_244),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_241),
.Y(n_355)
);

INVx4_ASAP7_75t_SL g409 ( 
.A(n_241),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g320 ( 
.A1(n_244),
.A2(n_321),
.B(n_323),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_244),
.A2(n_267),
.B(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_248),
.B(n_379),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_249),
.B(n_334),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_282),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_255),
.B(n_258),
.C(n_282),
.Y(n_434)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_268),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_259),
.B(n_268),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_265),
.B(n_266),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_266),
.B(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_277),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_289),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_285),
.Y(n_453)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_292),
.B(n_382),
.Y(n_381)
);

AOI21x1_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_388),
.B(n_393),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_371),
.B(n_387),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_346),
.B(n_370),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_319),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_297),
.B(n_319),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_316),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_298),
.B(n_316),
.Y(n_368)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx5_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_318),
.B(n_334),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_332),
.Y(n_319)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_332)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_333),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_334),
.A2(n_446),
.B(n_447),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_337),
.Y(n_413)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_343),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_344),
.C(n_373),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_365),
.B(n_369),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_361),
.B(n_364),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_356),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_363),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_368),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_374),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_384),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_380),
.B2(n_381),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_381),
.C(n_384),
.Y(n_392)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_379),
.Y(n_417)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g450 ( 
.A(n_383),
.B(n_451),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_385),
.A2(n_478),
.B(n_498),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_392),
.Y(n_393)
);

NOR3xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_437),
.C(n_458),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_433),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_397),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_426),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_398),
.B(n_426),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_405),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_399),
.B(n_406),
.C(n_439),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.C(n_402),
.Y(n_399)
);

XOR2x1_ASAP7_75t_SL g428 ( 
.A(n_400),
.B(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_401),
.A2(n_402),
.B1(n_403),
.B2(n_430),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_401),
.Y(n_430)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_418),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_410),
.Y(n_406)
);

AOI21x1_ASAP7_75t_SL g455 ( 
.A1(n_407),
.A2(n_411),
.B(n_417),
.Y(n_455)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_417),
.Y(n_410)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_412),
.Y(n_446)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_418),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_423),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_421),
.Y(n_432)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_424),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_431),
.C(n_432),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_432),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_434),
.B(n_435),
.Y(n_484)
);

A2O1A1Ixp33_ASAP7_75t_L g481 ( 
.A1(n_437),
.A2(n_482),
.B(n_483),
.C(n_485),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_438),
.B(n_440),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_441),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_448),
.B1(n_456),
.B2(n_457),
.Y(n_442)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_456),
.C(n_460),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_448),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_455),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.Y(n_449)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_450),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_452),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_463),
.C(n_464),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_458),
.Y(n_486)
);

NOR2x1_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_461),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_461),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_465),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_466),
.C(n_500),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_466),
.A2(n_472),
.B1(n_479),
.B2(n_480),
.Y(n_465)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

OA21x2_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_470),
.B(n_471),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_470),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_471),
.A2(n_492),
.B1(n_493),
.B2(n_496),
.Y(n_491)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_471),
.Y(n_496)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_472),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_474),
.B1(n_477),
.B2(n_478),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_475),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_475),
.Y(n_498)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_477),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_480),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_501),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_499),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_499),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_497),
.Y(n_490)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_496),
.C(n_497),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_501),
.A2(n_507),
.B(n_508),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_505),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_505),
.Y(n_508)
);


endmodule