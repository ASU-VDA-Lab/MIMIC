module real_jpeg_32344_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_SL g125 ( 
.A(n_0),
.Y(n_125)
);

OAI22x1_ASAP7_75t_SL g151 ( 
.A1(n_0),
.A2(n_125),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

AOI22x1_ASAP7_75t_L g209 ( 
.A1(n_0),
.A2(n_125),
.B1(n_210),
.B2(n_213),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_0),
.B(n_110),
.Y(n_289)
);

OAI22x1_ASAP7_75t_SL g306 ( 
.A1(n_0),
.A2(n_125),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_0),
.A2(n_316),
.A3(n_321),
.B1(n_325),
.B2(n_332),
.Y(n_315)
);

NAND2xp67_ASAP7_75t_SL g415 ( 
.A(n_0),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_0),
.B(n_237),
.Y(n_420)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_1),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_1),
.Y(n_295)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_1),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_2),
.B(n_498),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_2),
.B(n_497),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_5),
.Y(n_301)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_5),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_6),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_7),
.A2(n_55),
.B1(n_87),
.B2(n_90),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_55),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_7),
.A2(n_55),
.B1(n_504),
.B2(n_508),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_8),
.A2(n_48),
.B(n_51),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_8),
.B(n_52),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_8),
.A2(n_164),
.B1(n_169),
.B2(n_171),
.Y(n_163)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_8),
.A2(n_171),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_8),
.A2(n_171),
.B1(n_256),
.B2(n_259),
.Y(n_255)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_12),
.A2(n_116),
.B1(n_118),
.B2(n_122),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_12),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_12),
.A2(n_122),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_12),
.A2(n_122),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

OAI22x1_ASAP7_75t_L g297 ( 
.A1(n_12),
.A2(n_122),
.B1(n_298),
.B2(n_302),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_13),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_496),
.B(n_513),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_175),
.B(n_493),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_16),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_157),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_17),
.B(n_157),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.C(n_144),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_18),
.A2(n_19),
.B1(n_138),
.B2(n_139),
.Y(n_278)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_96),
.B2(n_134),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_67),
.B2(n_95),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_23),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_47),
.B1(n_54),
.B2(n_65),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_24),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_24),
.Y(n_161)
);

AOI22x1_ASAP7_75t_L g243 ( 
.A1(n_24),
.A2(n_149),
.B1(n_151),
.B2(n_228),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_33),
.Y(n_349)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_34),
.Y(n_156)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_37),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_38),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_38),
.B(n_125),
.Y(n_392)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_39),
.Y(n_403)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_41),
.Y(n_253)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_47),
.Y(n_147)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_49),
.Y(n_331)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_50),
.Y(n_232)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_54),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_64),
.Y(n_320)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21x1_ASAP7_75t_L g444 ( 
.A1(n_66),
.A2(n_161),
.B(n_226),
.Y(n_444)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_67),
.B(n_134),
.C(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_86),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_68),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_77),
.Y(n_68)
);

OAI21x1_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_78),
.B(n_81),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_69),
.Y(n_206)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_69),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_69),
.A2(n_77),
.B1(n_209),
.B2(n_248),
.Y(n_247)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_70),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_71),
.Y(n_418)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_76),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_76),
.Y(n_190)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_76),
.Y(n_258)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_76),
.Y(n_261)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_76),
.Y(n_304)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_77),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_SL g406 ( 
.A1(n_78),
.A2(n_125),
.B(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NOR2xp67_ASAP7_75t_R g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_85),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_85),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_86),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_234)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_94),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_139),
.C(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_95),
.B(n_146),
.Y(n_271)
);

AO22x1_ASAP7_75t_L g468 ( 
.A1(n_96),
.A2(n_242),
.B1(n_243),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_96),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_115),
.B1(n_123),
.B2(n_133),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_115),
.B1(n_123),
.B2(n_133),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_97),
.B(n_133),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_97),
.A2(n_133),
.B1(n_163),
.B2(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_124),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_105),
.B2(n_107),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_101),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_101),
.Y(n_356)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_106),
.Y(n_507)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_111),
.Y(n_359)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_113),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_133),
.B(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_117),
.Y(n_170)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_121),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_125),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_125),
.B(n_401),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_127),
.Y(n_509)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_128),
.A2(n_344),
.A3(n_347),
.B1(n_350),
.B2(n_353),
.Y(n_343)
);

OAI32xp33_ASAP7_75t_L g365 ( 
.A1(n_128),
.A2(n_344),
.A3(n_347),
.B1(n_350),
.B2(n_353),
.Y(n_365)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_163),
.B(n_172),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_134),
.B(n_241),
.C(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_134),
.B(n_312),
.C(n_436),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_135),
.B(n_224),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g366 ( 
.A(n_139),
.B(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_139),
.B(n_473),
.C(n_474),
.Y(n_472)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_140),
.B(n_271),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_141),
.B(n_241),
.C(n_368),
.Y(n_450)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_142),
.B(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_144),
.Y(n_277)
);

INVxp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B(n_150),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_161),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_148),
.A2(n_161),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_157),
.Y(n_518)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_162),
.CI(n_173),
.CON(n_157),
.SN(n_157)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_158),
.B(n_162),
.C(n_173),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_176),
.A2(n_514),
.B(n_515),
.C(n_516),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_279),
.B(n_489),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_273),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_266),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_179),
.B(n_266),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_222),
.C(n_239),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XOR2x1_ASAP7_75t_L g462 ( 
.A(n_181),
.B(n_222),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_214),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_182),
.A2(n_215),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_198),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_183),
.Y(n_215)
);

XOR2x2_ASAP7_75t_L g470 ( 
.A(n_183),
.B(n_198),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_191),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_184),
.Y(n_265)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_191),
.B(n_306),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_192),
.A2(n_255),
.B1(n_262),
.B2(n_265),
.Y(n_254)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_193),
.B(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_193),
.A2(n_297),
.B1(n_306),
.B2(n_362),
.Y(n_361)
);

NOR2x1_ASAP7_75t_R g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g197 ( 
.A(n_194),
.Y(n_197)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22x1_ASAP7_75t_L g377 ( 
.A1(n_208),
.A2(n_237),
.B1(n_369),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_209),
.Y(n_369)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B(n_219),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_238),
.Y(n_222)
);

NAND2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_233),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_224),
.A2(n_286),
.B1(n_287),
.B2(n_312),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_224),
.B(n_288),
.C(n_311),
.Y(n_340)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_234),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_225),
.Y(n_312)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_238),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_239),
.B(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_240),
.B(n_464),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_241),
.A2(n_242),
.B1(n_368),
.B2(n_370),
.Y(n_367)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_241),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_241),
.A2(n_242),
.B1(n_376),
.B2(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g467 ( 
.A(n_245),
.B(n_468),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_284),
.C(n_313),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_246),
.A2(n_313),
.B1(n_314),
.B2(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_246),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_246),
.B(n_360),
.C(n_392),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_246),
.A2(n_247),
.B1(n_392),
.B2(n_427),
.Y(n_426)
);

AO22x1_ASAP7_75t_L g438 ( 
.A1(n_246),
.A2(n_254),
.B1(n_382),
.B2(n_439),
.Y(n_438)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_248),
.Y(n_378)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_254),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_255),
.A2(n_262),
.B(n_305),
.Y(n_442)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_258),
.Y(n_307)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx4f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_270),
.C(n_272),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_274),
.A2(n_491),
.B(n_492),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_275),
.B(n_276),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_457),
.B(n_486),
.Y(n_279)
);

AOI211x1_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_383),
.B(n_431),
.C(n_456),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_371),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_338),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_283),
.B(n_338),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_285),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_311),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_290),
.B(n_414),
.Y(n_413)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_296),
.B(n_305),
.Y(n_290)
);

INVx3_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_295),
.Y(n_416)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_301),
.Y(n_411)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_311),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_311),
.B(n_397),
.Y(n_422)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_337),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_315),
.B(n_337),
.Y(n_379)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_366),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_340),
.B(n_366),
.C(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_341),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_360),
.B1(n_361),
.B2(n_365),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_343),
.B(n_360),
.Y(n_436)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_360),
.B(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_R g419 ( 
.A(n_361),
.B(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_361),
.B(n_420),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_368),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_380),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_380),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.C(n_379),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_376),
.A2(n_390),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_399),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_376),
.B(n_442),
.Y(n_441)
);

XOR2x2_ASAP7_75t_L g449 ( 
.A(n_376),
.B(n_442),
.Y(n_449)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_393),
.B(n_429),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_388),
.B(n_391),
.Y(n_430)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_392),
.Y(n_427)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_423),
.B(n_428),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_396),
.A2(n_412),
.B(n_422),
.Y(n_395)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_404),
.B(n_406),
.Y(n_399)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

AOI21x1_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_419),
.B(n_421),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_SL g428 ( 
.A(n_424),
.B(n_425),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_451),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_459),
.Y(n_458)
);

NAND2x1_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_445),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_437),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_437),
.Y(n_476)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_448),
.Y(n_447)
);

XNOR2x1_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_438),
.B(n_480),
.C(n_482),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_441),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_444),
.Y(n_473)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_445),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_449),
.C(n_450),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_455),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_450),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_454),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_454),
.Y(n_459)
);

NAND4xp25_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.C(n_475),
.D(n_478),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_460),
.A2(n_487),
.B(n_488),
.Y(n_486)
);

AO21x1_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_463),
.B(n_465),
.Y(n_460)
);

AND3x1_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_463),
.C(n_465),
.Y(n_487)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_462),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_470),
.C(n_471),
.Y(n_465)
);

OAI22x1_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_467),
.B1(n_470),
.B2(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_483),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_483),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_490),
.Y(n_489)
);

NOR3xp33_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_497),
.C(n_500),
.Y(n_515)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_499),
.Y(n_496)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_511),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_510),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_502),
.B(n_510),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);


endmodule