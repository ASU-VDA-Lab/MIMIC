module fake_ariane_1612_n_1678 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1678);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1678;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_24),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_33),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_25),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_18),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_28),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_61),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_10),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_32),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_79),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_88),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_93),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_74),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_16),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_71),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_51),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_2),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_91),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_17),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_115),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_123),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_55),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_48),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_107),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_41),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_82),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_17),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_97),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_12),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_120),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_24),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_81),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_63),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_67),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_80),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_19),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_19),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_52),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_69),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_15),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_45),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_73),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_26),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_125),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_13),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_29),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_84),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_16),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_43),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_5),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_53),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_70),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_4),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_127),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_43),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_129),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_75),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_14),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_57),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_30),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_89),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_132),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_108),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_98),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_65),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_101),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_44),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_119),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_111),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_59),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_117),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_78),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_48),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_146),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_31),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_47),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_52),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_56),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_135),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_40),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_33),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_38),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_27),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_6),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_124),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_106),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_60),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g260 ( 
.A(n_44),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_31),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_39),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_109),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_114),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_77),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_149),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_62),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_8),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_49),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_12),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_15),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_151),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_50),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_7),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_102),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_30),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_18),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_66),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_22),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_50),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_35),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_130),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_90),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_64),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_143),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_4),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_133),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_49),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_41),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_46),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_2),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_27),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_26),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_72),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_94),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_51),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_20),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_39),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_7),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_83),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_131),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_118),
.Y(n_304)
);

BUFx2_ASAP7_75t_SL g305 ( 
.A(n_122),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_11),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_165),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_236),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_241),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_259),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_175),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_280),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_284),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_303),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_215),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_260),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_260),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_165),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_246),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_245),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_306),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_250),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_175),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_225),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_190),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_225),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_154),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_156),
.B(n_0),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_156),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_155),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_162),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_281),
.B(n_0),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_278),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_162),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_178),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_157),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_178),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_186),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_248),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_186),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_159),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_160),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_188),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_205),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_188),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_205),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_166),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_170),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_172),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_248),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_174),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_179),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_163),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_195),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_195),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_196),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_196),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_197),
.B(n_1),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_249),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_197),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_200),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_210),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_163),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_200),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_163),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_201),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_163),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_201),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_281),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_311),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_299),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_316),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_333),
.B(n_299),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_318),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_329),
.Y(n_389)
);

NAND2xp33_ASAP7_75t_L g390 ( 
.A(n_341),
.B(n_299),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_318),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_L g392 ( 
.A(n_341),
.B(n_299),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_317),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_321),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_331),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_321),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_333),
.B(n_299),
.Y(n_398)
);

AND3x1_ASAP7_75t_L g399 ( 
.A(n_337),
.B(n_219),
.C(n_210),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_344),
.B(n_235),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_322),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_331),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_322),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_334),
.Y(n_405)
);

BUFx8_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_334),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_338),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_344),
.Y(n_410)
);

AND2x2_ASAP7_75t_SL g411 ( 
.A(n_342),
.B(n_161),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

BUFx12f_ASAP7_75t_L g413 ( 
.A(n_324),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_345),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_347),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_313),
.B(n_330),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_350),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_353),
.B(n_207),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_364),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_364),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

OA21x2_ASAP7_75t_L g430 ( 
.A1(n_365),
.A2(n_209),
.B(n_207),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_366),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_366),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_367),
.B(n_209),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_370),
.B(n_211),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_370),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_371),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_374),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_328),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_308),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_376),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_415),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_335),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_442),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_369),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_411),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_363),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_410),
.B(n_336),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_413),
.Y(n_454)
);

NAND2x1p5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_376),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_387),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_411),
.B(n_349),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_L g459 ( 
.A(n_410),
.B(n_340),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_349),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_368),
.B1(n_354),
.B2(n_356),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_410),
.Y(n_462)
);

BUFx10_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_369),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_393),
.B(n_326),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_387),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_422),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_394),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_430),
.A2(n_372),
.B1(n_342),
.B2(n_378),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_380),
.Y(n_471)
);

AOI21x1_ASAP7_75t_L g472 ( 
.A1(n_381),
.A2(n_223),
.B(n_211),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_L g473 ( 
.A(n_410),
.B(n_351),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_426),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_352),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_400),
.B(n_357),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_413),
.B(n_335),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_430),
.A2(n_377),
.B1(n_375),
.B2(n_373),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_399),
.A2(n_362),
.B1(n_361),
.B2(n_359),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_387),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_414),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_413),
.Y(n_485)
);

BUFx10_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_416),
.B(n_428),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_380),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_389),
.Y(n_489)
);

CKINVDCx6p67_ASAP7_75t_R g490 ( 
.A(n_440),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_431),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_387),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_400),
.B(n_358),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_393),
.B(n_346),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_407),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_385),
.A2(n_360),
.B1(n_255),
.B2(n_282),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_416),
.B(n_309),
.Y(n_499)
);

OAI22xp33_ASAP7_75t_L g500 ( 
.A1(n_423),
.A2(n_247),
.B1(n_199),
.B2(n_254),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_379),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_416),
.B(n_310),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_416),
.B(n_307),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_431),
.B(n_323),
.Y(n_505)
);

BUFx8_ASAP7_75t_SL g506 ( 
.A(n_379),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_387),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_381),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_414),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_432),
.B(n_312),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_432),
.B(n_332),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g512 ( 
.A(n_379),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_414),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_437),
.B(n_314),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_407),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_437),
.B(n_332),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_423),
.B(n_315),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_430),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_385),
.B(n_223),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_430),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_383),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_438),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_407),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_438),
.B(n_319),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_443),
.B(n_264),
.Y(n_525)
);

NOR2x1p5_ASAP7_75t_L g526 ( 
.A(n_434),
.B(n_219),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_396),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_L g528 ( 
.A1(n_434),
.A2(n_212),
.B1(n_183),
.B2(n_185),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_396),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_394),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_396),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_383),
.B(n_164),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_385),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_435),
.B(n_230),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_396),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_394),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_385),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_412),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_384),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_414),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_406),
.B(n_189),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_412),
.Y(n_544)
);

OAI21xp33_ASAP7_75t_SL g545 ( 
.A1(n_435),
.A2(n_418),
.B(n_419),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_406),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_418),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_394),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_414),
.B(n_224),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_406),
.B(n_230),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_418),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_402),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_406),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_414),
.B(n_193),
.C(n_191),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_385),
.B(n_224),
.Y(n_555)
);

BUFx10_ASAP7_75t_L g556 ( 
.A(n_398),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_414),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_394),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_419),
.B(n_237),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_384),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_419),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_402),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_420),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_398),
.A2(n_279),
.B1(n_275),
.B2(n_237),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_386),
.B(n_234),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_420),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_398),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_386),
.B(n_164),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_406),
.B(n_202),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_419),
.B(n_251),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_388),
.B(n_234),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_421),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_421),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_402),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_420),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_394),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_388),
.B(n_238),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_391),
.B(n_238),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_398),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_421),
.B(n_251),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_398),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_420),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_421),
.B(n_273),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_394),
.Y(n_584)
);

INVx2_ASAP7_75t_SL g585 ( 
.A(n_425),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_420),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_425),
.Y(n_587)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_425),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_508),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_550),
.B(n_425),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_458),
.B(n_391),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_460),
.B(n_463),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_463),
.B(n_395),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_448),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_471),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_508),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_448),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_450),
.B(n_395),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_490),
.B(n_320),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_450),
.B(n_397),
.Y(n_600)
);

NAND2x1_ASAP7_75t_L g601 ( 
.A(n_563),
.B(n_429),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_521),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_451),
.B(n_429),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_550),
.B(n_429),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_471),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_470),
.B(n_397),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_484),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_461),
.B(n_401),
.Y(n_608)
);

BUFx8_ASAP7_75t_L g609 ( 
.A(n_465),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_446),
.A2(n_429),
.B1(n_439),
.B2(n_433),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_463),
.B(n_401),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_464),
.B(n_420),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_521),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_502),
.A2(n_273),
.B1(n_279),
.B2(n_295),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_517),
.B(n_403),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_449),
.B(n_403),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_510),
.A2(n_439),
.B1(n_433),
.B2(n_408),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_484),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_517),
.B(n_405),
.Y(n_619)
);

BUFx8_ASAP7_75t_L g620 ( 
.A(n_465),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_516),
.B(n_405),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_455),
.B(n_408),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_490),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_446),
.A2(n_520),
.B1(n_518),
.B2(n_452),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_506),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_541),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_525),
.B(n_409),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_488),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_560),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_455),
.B(n_420),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_504),
.B(n_433),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_446),
.A2(n_433),
.B1(n_439),
.B2(n_436),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_514),
.B(n_420),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_447),
.B(n_325),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_588),
.B(n_439),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_588),
.B(n_424),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_448),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_502),
.B(n_424),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_499),
.B(n_424),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_481),
.B(n_477),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_518),
.A2(n_441),
.B1(n_436),
.B2(n_427),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_494),
.B(n_424),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_445),
.B(n_424),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_457),
.B(n_424),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_520),
.A2(n_441),
.B1(n_436),
.B2(n_427),
.Y(n_646)
);

BUFx5_ASAP7_75t_L g647 ( 
.A(n_486),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_560),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_535),
.A2(n_441),
.B1(n_436),
.B2(n_427),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_468),
.Y(n_650)
);

BUFx8_ASAP7_75t_L g651 ( 
.A(n_454),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_474),
.B(n_424),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_535),
.A2(n_567),
.B1(n_579),
.B2(n_519),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_512),
.B(n_424),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_489),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_475),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_512),
.B(n_441),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_478),
.B(n_275),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_491),
.B(n_427),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_495),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_492),
.B(n_522),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_531),
.B(n_427),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_567),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_505),
.B(n_427),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_487),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_455),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_503),
.B(n_427),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_550),
.A2(n_441),
.B1(n_436),
.B2(n_427),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_511),
.B(n_585),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_545),
.A2(n_240),
.B(n_296),
.C(n_268),
.Y(n_670)
);

OAI22xp33_ASAP7_75t_L g671 ( 
.A1(n_550),
.A2(n_295),
.B1(n_301),
.B2(n_300),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_506),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_583),
.A2(n_441),
.B1(n_436),
.B2(n_404),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_478),
.B(n_327),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_585),
.B(n_436),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_478),
.B(n_300),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_559),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_526),
.B(n_436),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_485),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_559),
.B(n_441),
.Y(n_680)
);

INVxp33_ASAP7_75t_L g681 ( 
.A(n_496),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_579),
.A2(n_441),
.B1(n_240),
.B2(n_296),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_579),
.B(n_402),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_570),
.B(n_404),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_570),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_580),
.B(n_404),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_580),
.Y(n_687)
);

INVx8_ASAP7_75t_L g688 ( 
.A(n_478),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_533),
.B(n_404),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_498),
.B(n_343),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_568),
.B(n_239),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_SL g692 ( 
.A1(n_553),
.A2(n_546),
.B1(n_555),
.B2(n_519),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_536),
.A2(n_268),
.B(n_239),
.C(n_244),
.Y(n_693)
);

AND2x2_ASAP7_75t_SL g694 ( 
.A(n_479),
.B(n_161),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_539),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_497),
.B(n_244),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_528),
.B(n_203),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_497),
.B(n_258),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_501),
.B(n_258),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_501),
.B(n_287),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_448),
.B(n_287),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_527),
.Y(n_702)
);

NOR2xp67_ASAP7_75t_L g703 ( 
.A(n_485),
.B(n_158),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_536),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_515),
.B(n_301),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_515),
.B(n_206),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_523),
.B(n_208),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_523),
.B(n_214),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_448),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_540),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_544),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_547),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_553),
.B(n_216),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_551),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_519),
.B(n_217),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_527),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_579),
.B(n_221),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_529),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_561),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_565),
.A2(n_392),
.B(n_390),
.C(n_382),
.Y(n_720)
);

NAND3xp33_ASAP7_75t_L g721 ( 
.A(n_453),
.B(n_272),
.C(n_228),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_519),
.B(n_226),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_538),
.B(n_233),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_538),
.B(n_243),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_572),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_519),
.B(n_252),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_538),
.B(n_233),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_524),
.B(n_253),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_538),
.B(n_270),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_573),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_529),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_519),
.B(n_555),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_539),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_543),
.B(n_190),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_532),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_500),
.B(n_256),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_569),
.B(n_583),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_583),
.B(n_261),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_539),
.B(n_262),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_583),
.A2(n_267),
.B1(n_305),
.B2(n_285),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_537),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_555),
.B(n_265),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_556),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_555),
.B(n_265),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_587),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_556),
.B(n_263),
.Y(n_746)
);

AND2x6_ASAP7_75t_L g747 ( 
.A(n_538),
.B(n_270),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_555),
.B(n_269),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_555),
.A2(n_267),
.B1(n_305),
.B2(n_297),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_537),
.B(n_271),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_552),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_622),
.A2(n_530),
.B(n_469),
.Y(n_752)
);

OAI321xp33_ASAP7_75t_L g753 ( 
.A1(n_671),
.A2(n_564),
.A3(n_577),
.B1(n_578),
.B2(n_571),
.C(n_472),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_622),
.A2(n_576),
.B(n_548),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_640),
.A2(n_459),
.B(n_453),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_615),
.B(n_556),
.Y(n_756)
);

BUFx8_ASAP7_75t_L g757 ( 
.A(n_625),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_615),
.A2(n_552),
.B(n_562),
.C(n_574),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_631),
.A2(n_476),
.B(n_459),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_631),
.A2(n_480),
.B(n_462),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_619),
.B(n_581),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_702),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_635),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_590),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_650),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_592),
.B(n_558),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_716),
.Y(n_767)
);

BUFx4f_ASAP7_75t_L g768 ( 
.A(n_688),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_694),
.A2(n_562),
.B1(n_574),
.B2(n_549),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_619),
.B(n_581),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_594),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_675),
.A2(n_632),
.B(n_612),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_664),
.A2(n_473),
.B(n_476),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_616),
.B(n_581),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_689),
.A2(n_473),
.B(n_462),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_713),
.B(n_276),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_594),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_651),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_656),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_637),
.A2(n_467),
.B(n_480),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_623),
.B(n_599),
.Y(n_781)
);

CKINVDCx10_ASAP7_75t_R g782 ( 
.A(n_658),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_590),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_593),
.B(n_563),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_738),
.B(n_283),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_593),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_628),
.A2(n_467),
.B(n_582),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_665),
.A2(n_483),
.B(n_582),
.Y(n_788)
);

NOR2x1p5_ASAP7_75t_SL g789 ( 
.A(n_647),
.B(n_472),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_611),
.B(n_563),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_611),
.A2(n_624),
.B1(n_592),
.B2(n_704),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_591),
.B(n_586),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_695),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_718),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_636),
.A2(n_483),
.B(n_557),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_647),
.B(n_558),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_661),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_731),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_695),
.Y(n_799)
);

O2A1O1Ixp33_ASAP7_75t_SL g800 ( 
.A1(n_670),
.A2(n_557),
.B(n_566),
.C(n_586),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_591),
.A2(n_549),
.B(n_444),
.C(n_509),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_669),
.A2(n_507),
.B(n_482),
.Y(n_802)
);

AOI22x1_ASAP7_75t_L g803 ( 
.A1(n_719),
.A2(n_586),
.B1(n_542),
.B2(n_444),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_621),
.B(n_444),
.Y(n_804)
);

BUFx4f_ASAP7_75t_L g805 ( 
.A(n_688),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_680),
.A2(n_507),
.B(n_482),
.Y(n_806)
);

OAI21xp33_ASAP7_75t_L g807 ( 
.A1(n_691),
.A2(n_292),
.B(n_288),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_704),
.A2(n_534),
.B(n_509),
.C(n_566),
.Y(n_808)
);

CKINVDCx10_ASAP7_75t_R g809 ( 
.A(n_658),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_641),
.B(n_509),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_642),
.A2(n_534),
.B(n_542),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_642),
.A2(n_534),
.B(n_542),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_697),
.A2(n_566),
.B(n_392),
.C(n_390),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_666),
.A2(n_584),
.B(n_558),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_624),
.A2(n_466),
.B1(n_584),
.B2(n_558),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_646),
.A2(n_554),
.B(n_466),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_651),
.Y(n_817)
);

AO21x2_ASAP7_75t_L g818 ( 
.A1(n_723),
.A2(n_382),
.B(n_558),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_647),
.B(n_653),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_666),
.A2(n_584),
.B(n_466),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_646),
.A2(n_584),
.B(n_575),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_610),
.B(n_584),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_639),
.A2(n_575),
.B(n_513),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_717),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_634),
.A2(n_601),
.B(n_644),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_735),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_645),
.A2(n_493),
.B(n_456),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_677),
.A2(n_290),
.B(n_291),
.C(n_293),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_685),
.B(n_456),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_609),
.Y(n_830)
);

OAI321xp33_ASAP7_75t_L g831 ( 
.A1(n_671),
.A2(n_294),
.A3(n_298),
.B1(n_267),
.B2(n_9),
.C(n_11),
.Y(n_831)
);

BUFx12f_ASAP7_75t_L g832 ( 
.A(n_609),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_647),
.B(n_733),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_687),
.B(n_493),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_652),
.A2(n_575),
.B(n_513),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_647),
.B(n_733),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_739),
.B(n_513),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_710),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_711),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_737),
.B(n_513),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_741),
.Y(n_841)
);

NOR3xp33_ASAP7_75t_L g842 ( 
.A(n_728),
.B(n_285),
.C(n_297),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_658),
.B(n_513),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_659),
.A2(n_575),
.B(n_486),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_739),
.B(n_575),
.Y(n_845)
);

NOR3xp33_ASAP7_75t_L g846 ( 
.A(n_728),
.B(n_302),
.C(n_198),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_746),
.B(n_486),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_746),
.B(n_167),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_662),
.A2(n_304),
.B(n_168),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_676),
.B(n_302),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_614),
.A2(n_3),
.B(n_5),
.C(n_8),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_712),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_684),
.A2(n_686),
.B(n_600),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_751),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_676),
.B(n_604),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_595),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_614),
.A2(n_3),
.B(n_9),
.C(n_14),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_654),
.A2(n_289),
.B(n_286),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_654),
.A2(n_277),
.B(n_274),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_657),
.B(n_633),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_714),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_679),
.B(n_672),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_647),
.B(n_194),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_681),
.B(n_20),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_676),
.B(n_267),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_657),
.B(n_266),
.Y(n_866)
);

NOR2x1_ASAP7_75t_L g867 ( 
.A(n_703),
.B(n_717),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_617),
.A2(n_242),
.B(n_232),
.C(n_231),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_633),
.A2(n_229),
.B1(n_227),
.B2(n_222),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_594),
.B(n_220),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_743),
.A2(n_218),
.B1(n_213),
.B2(n_204),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_674),
.B(n_21),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_598),
.A2(n_192),
.B(n_187),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_620),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_594),
.B(n_597),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_667),
.A2(n_184),
.B(n_182),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_605),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_598),
.A2(n_181),
.B(n_180),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_597),
.B(n_177),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_683),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_667),
.A2(n_643),
.B(n_745),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_725),
.A2(n_176),
.B(n_173),
.Y(n_882)
);

NAND3xp33_ASAP7_75t_L g883 ( 
.A(n_736),
.B(n_171),
.C(n_169),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_589),
.B(n_21),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_730),
.A2(n_86),
.B(n_148),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_694),
.B(n_22),
.Y(n_886)
);

AOI21xp33_ASAP7_75t_L g887 ( 
.A1(n_740),
.A2(n_749),
.B(n_690),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_607),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_596),
.B(n_602),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_597),
.A2(n_76),
.B(n_147),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_618),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_683),
.A2(n_663),
.B(n_613),
.C(n_626),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_678),
.A2(n_58),
.B(n_142),
.Y(n_893)
);

CKINVDCx8_ASAP7_75t_R g894 ( 
.A(n_688),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_638),
.A2(n_153),
.B(n_140),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_638),
.A2(n_138),
.B(n_137),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_638),
.A2(n_709),
.B(n_606),
.Y(n_897)
);

INVx11_ASAP7_75t_L g898 ( 
.A(n_620),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_627),
.B(n_23),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_705),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_709),
.A2(n_136),
.B(n_134),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_630),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_709),
.A2(n_121),
.B(n_113),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_648),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_750),
.A2(n_105),
.B(n_104),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_734),
.Y(n_906)
);

AND2x2_ASAP7_75t_SL g907 ( 
.A(n_749),
.B(n_23),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_706),
.A2(n_100),
.B(n_96),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_732),
.B(n_25),
.Y(n_909)
);

INVxp33_ASAP7_75t_SL g910 ( 
.A(n_715),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_734),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_740),
.B(n_28),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_707),
.A2(n_95),
.B(n_87),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_708),
.A2(n_608),
.B(n_655),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_742),
.B(n_32),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_722),
.B(n_34),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_673),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_693),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_604),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_629),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_660),
.A2(n_54),
.B(n_40),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_742),
.B(n_744),
.Y(n_922)
);

AO22x1_ASAP7_75t_L g923 ( 
.A1(n_744),
.A2(n_37),
.B1(n_42),
.B2(n_46),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_726),
.B(n_42),
.Y(n_924)
);

AOI21x1_ASAP7_75t_L g925 ( 
.A1(n_723),
.A2(n_47),
.B(n_53),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_721),
.A2(n_54),
.B(n_729),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_747),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_747),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_603),
.B(n_692),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_603),
.B(n_692),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_748),
.B(n_682),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_756),
.A2(n_724),
.B(n_668),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_761),
.A2(n_668),
.B(n_727),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_765),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_770),
.A2(n_727),
.B(n_729),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_786),
.A2(n_720),
.B(n_649),
.C(n_698),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_847),
.A2(n_701),
.B(n_696),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_763),
.B(n_785),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_792),
.A2(n_701),
.B(n_699),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_887),
.A2(n_603),
.B1(n_673),
.B2(n_700),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_779),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_786),
.B(n_603),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_824),
.B(n_603),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_855),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_797),
.B(n_747),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_R g946 ( 
.A(n_817),
.B(n_747),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_824),
.B(n_747),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_853),
.A2(n_790),
.B(n_784),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_880),
.A2(n_774),
.B1(n_791),
.B2(n_907),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_SL g950 ( 
.A(n_848),
.B(n_793),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_916),
.A2(n_924),
.B(n_846),
.C(n_810),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_855),
.B(n_910),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_907),
.B(n_843),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_916),
.A2(n_924),
.B(n_846),
.C(n_810),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_838),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_757),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_762),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_919),
.B(n_764),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_783),
.B(n_776),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_783),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_SL g961 ( 
.A1(n_884),
.A2(n_899),
.B(n_793),
.C(n_799),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_768),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_781),
.B(n_872),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_864),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_886),
.A2(n_912),
.B(n_842),
.C(n_884),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_860),
.A2(n_904),
.B1(n_902),
.B2(n_861),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_900),
.B(n_839),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_842),
.A2(n_864),
.B1(n_862),
.B2(n_843),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_852),
.B(n_902),
.Y(n_969)
);

AO22x1_ASAP7_75t_L g970 ( 
.A1(n_830),
.A2(n_874),
.B1(n_865),
.B2(n_778),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_904),
.B(n_911),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_755),
.A2(n_819),
.B(n_796),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_801),
.A2(n_758),
.B(n_808),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_767),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_906),
.B(n_850),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_899),
.B(n_850),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_794),
.Y(n_977)
);

NAND3xp33_ASAP7_75t_L g978 ( 
.A(n_851),
.B(n_857),
.C(n_868),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_771),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_922),
.B(n_799),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_SL g981 ( 
.A1(n_760),
.A2(n_873),
.B(n_878),
.C(n_759),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_753),
.A2(n_831),
.B(n_807),
.C(n_892),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_898),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_804),
.B(n_840),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_819),
.A2(n_796),
.B(n_766),
.Y(n_985)
);

INVx5_ASAP7_75t_L g986 ( 
.A(n_927),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_840),
.B(n_889),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_798),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_766),
.A2(n_773),
.B(n_845),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_801),
.A2(n_917),
.B1(n_868),
.B2(n_929),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_828),
.A2(n_918),
.B(n_808),
.C(n_800),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_930),
.A2(n_822),
.B1(n_758),
.B2(n_915),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_837),
.A2(n_772),
.B(n_812),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_768),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_811),
.A2(n_814),
.B(n_836),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_828),
.A2(n_769),
.B1(n_829),
.B2(n_834),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_928),
.B(n_867),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_769),
.A2(n_909),
.B1(n_883),
.B2(n_931),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_894),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_805),
.B(n_832),
.Y(n_1000)
);

BUFx8_ASAP7_75t_L g1001 ( 
.A(n_782),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_909),
.A2(n_866),
.B1(n_777),
.B2(n_771),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_809),
.B(n_871),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_920),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_771),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_757),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_869),
.B(n_870),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_833),
.A2(n_863),
.B(n_823),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_863),
.A2(n_788),
.B(n_775),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_870),
.B(n_879),
.Y(n_1010)
);

AO32x2_ASAP7_75t_L g1011 ( 
.A1(n_815),
.A2(n_800),
.A3(n_914),
.B1(n_925),
.B2(n_923),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_856),
.B(n_891),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_877),
.B(n_888),
.Y(n_1013)
);

CKINVDCx16_ASAP7_75t_R g1014 ( 
.A(n_927),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_879),
.B(n_826),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_893),
.A2(n_881),
.B(n_897),
.C(n_926),
.Y(n_1016)
);

AOI211xp5_ASAP7_75t_L g1017 ( 
.A1(n_921),
.A2(n_876),
.B(n_882),
.C(n_859),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_777),
.B(n_927),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_841),
.B(n_854),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_818),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_875),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_818),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_875),
.B(n_858),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_820),
.A2(n_752),
.B(n_754),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_821),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_816),
.Y(n_1026)
);

BUFx4f_ASAP7_75t_L g1027 ( 
.A(n_813),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_806),
.A2(n_825),
.B(n_802),
.C(n_844),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_787),
.A2(n_780),
.B(n_835),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_795),
.A2(n_827),
.B(n_849),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_789),
.B(n_803),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_913),
.B(n_908),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_905),
.B(n_885),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_890),
.B(n_895),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_896),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_901),
.B(n_903),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_756),
.A2(n_770),
.B(n_761),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_786),
.A2(n_824),
.B(n_616),
.C(n_791),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_907),
.A2(n_797),
.B1(n_761),
.B2(n_770),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_801),
.A2(n_758),
.B(n_808),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_756),
.A2(n_770),
.B(n_761),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_907),
.A2(n_797),
.B1(n_761),
.B2(n_770),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_SL g1043 ( 
.A(n_846),
.B(n_447),
.C(n_442),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_765),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_763),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_786),
.B(n_615),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_763),
.B(n_690),
.Y(n_1047)
);

AOI221xp5_ASAP7_75t_L g1048 ( 
.A1(n_831),
.A2(n_614),
.B1(n_399),
.B2(n_449),
.C(n_446),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_786),
.B(n_615),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_786),
.B(n_615),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_756),
.A2(n_770),
.B(n_761),
.Y(n_1051)
);

OAI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_786),
.A2(n_517),
.B1(n_447),
.B2(n_442),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_907),
.A2(n_797),
.B1(n_761),
.B2(n_770),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_768),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_855),
.B(n_919),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_763),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_765),
.Y(n_1057)
);

AO32x2_ASAP7_75t_L g1058 ( 
.A1(n_791),
.A2(n_917),
.A3(n_815),
.B1(n_585),
.B2(n_911),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_766),
.A2(n_755),
.B(n_773),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_756),
.A2(n_770),
.B(n_761),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_766),
.A2(n_755),
.B(n_773),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_756),
.A2(n_770),
.B(n_761),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_786),
.B(n_308),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_763),
.B(n_690),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_756),
.A2(n_770),
.B(n_761),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_757),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_786),
.A2(n_824),
.B(n_616),
.C(n_791),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_951),
.A2(n_954),
.B(n_964),
.C(n_1052),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_972),
.A2(n_1061),
.B(n_1059),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_983),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_962),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_1056),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_SL g1074 ( 
.A1(n_1038),
.A2(n_1067),
.B1(n_1042),
.B2(n_1053),
.C(n_1039),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_1003),
.Y(n_1075)
);

BUFx10_ASAP7_75t_L g1076 ( 
.A(n_956),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1051),
.A2(n_1062),
.B(n_1060),
.Y(n_1077)
);

AO31x2_ASAP7_75t_L g1078 ( 
.A1(n_1020),
.A2(n_992),
.A3(n_1016),
.B(n_1002),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_1048),
.A2(n_1007),
.B(n_965),
.C(n_982),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_1063),
.B(n_1050),
.Y(n_1080)
);

OA21x2_ASAP7_75t_L g1081 ( 
.A1(n_989),
.A2(n_1040),
.B(n_973),
.Y(n_1081)
);

OA21x2_ASAP7_75t_L g1082 ( 
.A1(n_973),
.A2(n_1040),
.B(n_993),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_934),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1065),
.A2(n_1033),
.B(n_1032),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1039),
.A2(n_1053),
.B(n_1042),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_941),
.Y(n_1086)
);

NAND2x1p5_ASAP7_75t_L g1087 ( 
.A(n_962),
.B(n_994),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_1010),
.A2(n_978),
.B(n_949),
.C(n_998),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_968),
.B(n_966),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1029),
.A2(n_1024),
.B(n_1030),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1009),
.A2(n_1028),
.B(n_995),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_936),
.A2(n_990),
.B(n_933),
.Y(n_1092)
);

OAI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_976),
.A2(n_959),
.B1(n_1064),
.B2(n_1047),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_994),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1027),
.A2(n_984),
.B(n_1008),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1027),
.A2(n_932),
.B(n_1031),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1043),
.A2(n_961),
.B(n_981),
.C(n_990),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1034),
.A2(n_1036),
.B(n_937),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1045),
.B(n_938),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_960),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_998),
.A2(n_991),
.B(n_942),
.C(n_987),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_996),
.A2(n_985),
.B(n_939),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1025),
.A2(n_1035),
.B(n_935),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_957),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1015),
.A2(n_947),
.B(n_967),
.C(n_1017),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_963),
.B(n_952),
.Y(n_1106)
);

BUFx10_ASAP7_75t_L g1107 ( 
.A(n_1066),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_992),
.A2(n_996),
.A3(n_1023),
.B(n_1026),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_950),
.A2(n_1035),
.B(n_943),
.Y(n_1109)
);

BUFx4_ASAP7_75t_SL g1110 ( 
.A(n_1001),
.Y(n_1110)
);

AOI21xp33_ASAP7_75t_L g1111 ( 
.A1(n_945),
.A2(n_971),
.B(n_1019),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1055),
.B(n_1054),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1025),
.A2(n_969),
.B(n_940),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_953),
.A2(n_1044),
.B1(n_1057),
.B2(n_955),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1018),
.A2(n_979),
.B(n_980),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_944),
.B(n_975),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1004),
.A2(n_1013),
.B(n_1012),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_946),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1000),
.A2(n_970),
.B1(n_1006),
.B2(n_1014),
.Y(n_1119)
);

AO32x2_ASAP7_75t_L g1120 ( 
.A1(n_1021),
.A2(n_1058),
.A3(n_1005),
.B1(n_1011),
.B2(n_1022),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_958),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_986),
.A2(n_997),
.B(n_1058),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_974),
.A2(n_977),
.B(n_988),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1054),
.B(n_994),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1011),
.A2(n_986),
.B(n_999),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1054),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_983),
.A2(n_786),
.B1(n_761),
.B2(n_770),
.Y(n_1127)
);

INVx5_ASAP7_75t_L g1128 ( 
.A(n_1001),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_951),
.A2(n_954),
.B(n_982),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_SL g1130 ( 
.A1(n_1038),
.A2(n_1067),
.B1(n_857),
.B2(n_851),
.C(n_1042),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_934),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_SL g1132 ( 
.A1(n_951),
.A2(n_954),
.B(n_786),
.C(n_1046),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_934),
.Y(n_1133)
);

INVx5_ASAP7_75t_L g1134 ( 
.A(n_983),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_948),
.A2(n_1041),
.B(n_1037),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_957),
.Y(n_1137)
);

AOI221xp5_ASAP7_75t_SL g1138 ( 
.A1(n_1038),
.A2(n_1067),
.B1(n_857),
.B2(n_851),
.C(n_1042),
.Y(n_1138)
);

OAI22x1_ASAP7_75t_L g1139 ( 
.A1(n_968),
.A2(n_964),
.B1(n_1063),
.B2(n_442),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_957),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_948),
.A2(n_1041),
.B(n_1037),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1046),
.A2(n_786),
.B1(n_761),
.B2(n_770),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_SL g1143 ( 
.A1(n_1048),
.A2(n_857),
.B(n_851),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_1003),
.Y(n_1144)
);

AO21x1_ASAP7_75t_L g1145 ( 
.A1(n_1039),
.A2(n_1053),
.B(n_1042),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_1045),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_951),
.A2(n_954),
.B(n_1048),
.C(n_1038),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_SL g1148 ( 
.A1(n_951),
.A2(n_954),
.B(n_786),
.C(n_1046),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_951),
.A2(n_954),
.B(n_1048),
.C(n_1038),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_951),
.A2(n_954),
.B(n_1048),
.C(n_1038),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_970),
.B(n_688),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_948),
.A2(n_1041),
.B(n_1037),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_951),
.A2(n_954),
.B(n_1048),
.C(n_1038),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1055),
.B(n_962),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_948),
.A2(n_1041),
.B(n_1037),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1046),
.B(n_786),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1047),
.B(n_1064),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1020),
.A2(n_992),
.A3(n_1016),
.B(n_1002),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_962),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_934),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_948),
.A2(n_1041),
.B(n_1037),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1047),
.B(n_1064),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1056),
.Y(n_1169)
);

AO21x1_ASAP7_75t_L g1170 ( 
.A1(n_1039),
.A2(n_1053),
.B(n_1042),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_962),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_962),
.Y(n_1172)
);

NAND2xp33_ASAP7_75t_L g1173 ( 
.A(n_1046),
.B(n_756),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1055),
.B(n_962),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_951),
.A2(n_954),
.B(n_982),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1063),
.B(n_447),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_934),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_934),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1046),
.A2(n_786),
.B1(n_761),
.B2(n_770),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_934),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_983),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_962),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_948),
.A2(n_1041),
.B(n_1037),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_989),
.A2(n_1040),
.B(n_973),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_963),
.B(n_938),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1055),
.B(n_962),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1056),
.Y(n_1189)
);

INVx3_ASAP7_75t_SL g1190 ( 
.A(n_983),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1020),
.A2(n_992),
.A3(n_1016),
.B(n_1002),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_963),
.B(n_938),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_SL g1193 ( 
.A1(n_951),
.A2(n_954),
.B(n_786),
.C(n_1046),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1083),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1080),
.B(n_1070),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_1121),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1147),
.A2(n_1151),
.B1(n_1149),
.B2(n_1154),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1176),
.A2(n_1143),
.B1(n_1089),
.B2(n_1139),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1086),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1129),
.A2(n_1175),
.B1(n_1085),
.B2(n_1170),
.Y(n_1200)
);

AO22x1_ASAP7_75t_L g1201 ( 
.A1(n_1128),
.A2(n_1175),
.B1(n_1129),
.B2(n_1118),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1085),
.A2(n_1114),
.B1(n_1092),
.B2(n_1142),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1088),
.B(n_1081),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1131),
.Y(n_1204)
);

INVx6_ASAP7_75t_L g1205 ( 
.A(n_1134),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1079),
.A2(n_1068),
.B1(n_1143),
.B2(n_1188),
.Y(n_1206)
);

BUFx2_ASAP7_75t_SL g1207 ( 
.A(n_1134),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1133),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1164),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_1186),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1145),
.A2(n_1093),
.B1(n_1140),
.B2(n_1104),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1108),
.B(n_1161),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1137),
.A2(n_1192),
.B1(n_1114),
.B2(n_1173),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1177),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1166),
.A2(n_1111),
.B1(n_1146),
.B2(n_1179),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1178),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1180),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1071),
.Y(n_1218)
);

OAI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1092),
.A2(n_1101),
.B(n_1136),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1081),
.B(n_1185),
.Y(n_1220)
);

OAI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1106),
.A2(n_1156),
.B1(n_1157),
.B2(n_1150),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1123),
.A2(n_1152),
.B1(n_1183),
.B2(n_1168),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1160),
.B(n_1167),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1073),
.Y(n_1224)
);

INVx6_ASAP7_75t_L g1225 ( 
.A(n_1134),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1123),
.A2(n_1152),
.B1(n_1127),
.B2(n_1159),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1152),
.A2(n_1116),
.B1(n_1119),
.B2(n_1122),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1120),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1119),
.A2(n_1189),
.B1(n_1185),
.B2(n_1169),
.Y(n_1229)
);

OAI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1128),
.A2(n_1100),
.B1(n_1126),
.B2(n_1124),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1082),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1082),
.A2(n_1113),
.B1(n_1144),
.B2(n_1075),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1075),
.A2(n_1144),
.B1(n_1174),
.B2(n_1155),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1112),
.A2(n_1187),
.B1(n_1155),
.B2(n_1174),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_1128),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1120),
.Y(n_1236)
);

CKINVDCx6p67_ASAP7_75t_R g1237 ( 
.A(n_1181),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1105),
.A2(n_1095),
.B1(n_1181),
.B2(n_1097),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1112),
.A2(n_1187),
.B1(n_1163),
.B2(n_1171),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1163),
.A2(n_1182),
.B1(n_1171),
.B2(n_1126),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1181),
.A2(n_1098),
.B1(n_1096),
.B2(n_1102),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1190),
.A2(n_1074),
.B1(n_1077),
.B2(n_1072),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1115),
.Y(n_1243)
);

CKINVDCx6p67_ASAP7_75t_R g1244 ( 
.A(n_1076),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1130),
.A2(n_1138),
.B1(n_1074),
.B2(n_1148),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1132),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1193),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1108),
.B(n_1125),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1108),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1182),
.A2(n_1094),
.B1(n_1172),
.B2(n_1076),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1078),
.B(n_1191),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1107),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1094),
.Y(n_1253)
);

INVx6_ASAP7_75t_L g1254 ( 
.A(n_1087),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1172),
.A2(n_1109),
.B1(n_1138),
.B2(n_1130),
.Y(n_1255)
);

NAND2x1p5_ASAP7_75t_L g1256 ( 
.A(n_1103),
.B(n_1069),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1162),
.Y(n_1257)
);

OAI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1135),
.A2(n_1158),
.B1(n_1184),
.B2(n_1165),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1084),
.A2(n_1153),
.B(n_1141),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1162),
.B(n_1191),
.Y(n_1260)
);

BUFx4_ASAP7_75t_R g1261 ( 
.A(n_1191),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1091),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1090),
.A2(n_694),
.B1(n_1048),
.B2(n_479),
.Y(n_1263)
);

INVx5_ASAP7_75t_L g1264 ( 
.A(n_1152),
.Y(n_1264)
);

BUFx5_ASAP7_75t_L g1265 ( 
.A(n_1083),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1083),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1089),
.A2(n_694),
.B1(n_1048),
.B2(n_479),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1100),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1128),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1118),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1110),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1083),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1089),
.A2(n_694),
.B1(n_1048),
.B2(n_479),
.Y(n_1273)
);

INVx11_ASAP7_75t_L g1274 ( 
.A(n_1110),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1081),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1176),
.A2(n_1048),
.B1(n_1080),
.B2(n_1063),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1128),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1083),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1089),
.A2(n_694),
.B1(n_1048),
.B2(n_479),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1083),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1089),
.A2(n_694),
.B1(n_1048),
.B2(n_479),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1083),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1080),
.A2(n_1147),
.B1(n_1151),
.B2(n_1149),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1083),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1118),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1190),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1117),
.Y(n_1287)
);

BUFx10_ASAP7_75t_L g1288 ( 
.A(n_1176),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1083),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1083),
.Y(n_1290)
);

BUFx12f_ASAP7_75t_L g1291 ( 
.A(n_1128),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1129),
.A2(n_694),
.B1(n_406),
.B2(n_325),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1089),
.A2(n_694),
.B1(n_1048),
.B2(n_479),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1083),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1118),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1083),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1117),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1080),
.B(n_1176),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1190),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1089),
.A2(n_694),
.B1(n_1048),
.B2(n_479),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1129),
.B(n_1175),
.Y(n_1301)
);

BUFx2_ASAP7_75t_SL g1302 ( 
.A(n_1134),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1099),
.Y(n_1303)
);

BUFx12f_ASAP7_75t_L g1304 ( 
.A(n_1128),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1129),
.A2(n_694),
.B1(n_406),
.B2(n_325),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1143),
.A2(n_1048),
.B1(n_831),
.B2(n_550),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1249),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1231),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1275),
.Y(n_1309)
);

NAND2x1_ASAP7_75t_L g1310 ( 
.A(n_1241),
.B(n_1275),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1203),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1268),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1202),
.A2(n_1200),
.B1(n_1283),
.B2(n_1197),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1259),
.A2(n_1258),
.B(n_1257),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1265),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1220),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1276),
.A2(n_1301),
.B1(n_1206),
.B2(n_1306),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1264),
.B(n_1251),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1275),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1231),
.Y(n_1320)
);

AO21x1_ASAP7_75t_L g1321 ( 
.A1(n_1301),
.A2(n_1198),
.B(n_1245),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1262),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1265),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1265),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1231),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1212),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1262),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1212),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1228),
.B(n_1236),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1264),
.B(n_1251),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1196),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1243),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1287),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1287),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1297),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1194),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1260),
.B(n_1248),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1199),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1204),
.B(n_1208),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1256),
.Y(n_1340)
);

AND2x4_ASAP7_75t_SL g1341 ( 
.A(n_1237),
.B(n_1226),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1292),
.A2(n_1305),
.B1(n_1279),
.B2(n_1300),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1209),
.B(n_1214),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1216),
.B(n_1217),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1266),
.Y(n_1345)
);

CKINVDCx6p67_ASAP7_75t_R g1346 ( 
.A(n_1291),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1272),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1278),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1280),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1282),
.B(n_1284),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1294),
.Y(n_1352)
);

OAI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1298),
.A2(n_1195),
.B1(n_1210),
.B2(n_1223),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1261),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1296),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1261),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1238),
.A2(n_1242),
.B(n_1232),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1201),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1246),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1247),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1219),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1221),
.B(n_1288),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1211),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1215),
.B(n_1229),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1303),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1213),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1255),
.A2(n_1222),
.B(n_1227),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1224),
.B(n_1295),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1230),
.A2(n_1263),
.B(n_1293),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1270),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1285),
.Y(n_1371)
);

OR2x6_ASAP7_75t_L g1372 ( 
.A(n_1291),
.B(n_1304),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_SL g1373 ( 
.A(n_1285),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1205),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1271),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1225),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1288),
.B(n_1281),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1370),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1309),
.Y(n_1379)
);

AOI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1313),
.A2(n_1273),
.B1(n_1267),
.B2(n_1250),
.C(n_1233),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1313),
.A2(n_1253),
.B(n_1240),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1311),
.B(n_1316),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1311),
.B(n_1316),
.Y(n_1383)
);

OA21x2_ASAP7_75t_L g1384 ( 
.A1(n_1357),
.A2(n_1239),
.B(n_1234),
.Y(n_1384)
);

NAND3xp33_ASAP7_75t_L g1385 ( 
.A(n_1361),
.B(n_1253),
.C(n_1252),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1372),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1317),
.A2(n_1218),
.B(n_1207),
.C(n_1302),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1361),
.B(n_1252),
.C(n_1299),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_SL g1389 ( 
.A1(n_1317),
.A2(n_1277),
.B(n_1235),
.C(n_1269),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1342),
.A2(n_1277),
.B1(n_1269),
.B2(n_1235),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1321),
.A2(n_1362),
.B1(n_1366),
.B2(n_1364),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1357),
.A2(n_1271),
.B(n_1244),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1336),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1318),
.B(n_1330),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1331),
.B(n_1286),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1336),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1365),
.B(n_1286),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1365),
.B(n_1299),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1338),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1377),
.A2(n_1274),
.B(n_1254),
.Y(n_1400)
);

AO21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1315),
.A2(n_1323),
.B(n_1324),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1337),
.B(n_1339),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1337),
.B(n_1339),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1377),
.A2(n_1367),
.B(n_1358),
.Y(n_1404)
);

AOI211xp5_ASAP7_75t_L g1405 ( 
.A1(n_1321),
.A2(n_1353),
.B(n_1358),
.C(n_1364),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1310),
.A2(n_1309),
.B(n_1340),
.Y(n_1406)
);

AO32x2_ASAP7_75t_L g1407 ( 
.A1(n_1374),
.A2(n_1376),
.A3(n_1329),
.B1(n_1328),
.B2(n_1326),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1365),
.B(n_1322),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1337),
.B(n_1343),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1367),
.A2(n_1359),
.B(n_1360),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1375),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1338),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1366),
.A2(n_1363),
.B1(n_1369),
.B2(n_1341),
.Y(n_1413)
);

AO32x2_ASAP7_75t_L g1414 ( 
.A1(n_1374),
.A2(n_1376),
.A3(n_1328),
.B1(n_1326),
.B2(n_1312),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1333),
.A2(n_1334),
.B(n_1335),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1322),
.B(n_1345),
.Y(n_1416)
);

AOI221xp5_ASAP7_75t_L g1417 ( 
.A1(n_1345),
.A2(n_1355),
.B1(n_1347),
.B2(n_1348),
.C(n_1349),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_R g1418 ( 
.A(n_1372),
.B(n_1327),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1402),
.B(n_1319),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1402),
.B(n_1319),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1393),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1379),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1396),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1403),
.B(n_1409),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1391),
.A2(n_1369),
.B1(n_1367),
.B2(n_1356),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1394),
.B(n_1319),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1417),
.B(n_1344),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1399),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1412),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1401),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1403),
.B(n_1320),
.Y(n_1431)
);

INVxp67_ASAP7_75t_SL g1432 ( 
.A(n_1410),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1406),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1415),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1382),
.B(n_1383),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1408),
.B(n_1352),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1414),
.B(n_1325),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1405),
.A2(n_1369),
.B1(n_1341),
.B2(n_1354),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1414),
.B(n_1308),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1408),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1416),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1380),
.A2(n_1369),
.B1(n_1390),
.B2(n_1413),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1414),
.B(n_1308),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1411),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1414),
.B(n_1314),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1421),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1442),
.A2(n_1404),
.B1(n_1381),
.B2(n_1384),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1437),
.B(n_1414),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1445),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1437),
.B(n_1407),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1421),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1437),
.B(n_1407),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1423),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1433),
.Y(n_1454)
);

AOI221xp5_ASAP7_75t_L g1455 ( 
.A1(n_1442),
.A2(n_1389),
.B1(n_1392),
.B2(n_1387),
.C(n_1388),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1424),
.B(n_1407),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1439),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1432),
.B(n_1350),
.Y(n_1458)
);

OAI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1438),
.A2(n_1389),
.B1(n_1385),
.B2(n_1400),
.C(n_1418),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1439),
.B(n_1378),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1443),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1424),
.B(n_1407),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1443),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1443),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1445),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1435),
.B(n_1407),
.Y(n_1466)
);

AO21x2_ASAP7_75t_L g1467 ( 
.A1(n_1434),
.A2(n_1307),
.B(n_1332),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1425),
.A2(n_1384),
.B1(n_1354),
.B2(n_1356),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1432),
.B(n_1351),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1441),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1430),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1458),
.B(n_1441),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1446),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1470),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1446),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1446),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1449),
.B(n_1426),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1447),
.A2(n_1425),
.B1(n_1438),
.B2(n_1427),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1454),
.B(n_1422),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1450),
.B(n_1452),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1451),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1467),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1450),
.B(n_1452),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1450),
.B(n_1419),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1450),
.B(n_1419),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1452),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1458),
.B(n_1440),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1452),
.B(n_1420),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1451),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1448),
.B(n_1420),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1469),
.B(n_1428),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1448),
.B(n_1420),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1470),
.B(n_1429),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1466),
.B(n_1436),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1467),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1451),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1448),
.B(n_1431),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1448),
.B(n_1456),
.Y(n_1498)
);

CKINVDCx16_ASAP7_75t_R g1499 ( 
.A(n_1471),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1466),
.B(n_1436),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1453),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1456),
.B(n_1431),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1467),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1453),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1449),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1473),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1505),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1480),
.B(n_1456),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1478),
.A2(n_1459),
.B(n_1455),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1478),
.B(n_1466),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1474),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1473),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1486),
.B(n_1470),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1491),
.B(n_1466),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1493),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1486),
.B(n_1460),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1475),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1480),
.B(n_1456),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_1462),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1477),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1475),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1499),
.B(n_1462),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1486),
.B(n_1460),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1499),
.B(n_1462),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1476),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1476),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1472),
.B(n_1462),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1493),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1480),
.B(n_1471),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1505),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1481),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1481),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1489),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1474),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1483),
.B(n_1471),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1489),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1496),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1486),
.A2(n_1455),
.B1(n_1459),
.B2(n_1447),
.Y(n_1538)
);

NAND2x1p5_ASAP7_75t_L g1539 ( 
.A(n_1479),
.B(n_1386),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1486),
.B(n_1483),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1505),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1477),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1472),
.B(n_1427),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1483),
.A2(n_1447),
.B1(n_1455),
.B2(n_1449),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1501),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1505),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1506),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1509),
.B(n_1484),
.Y(n_1549)
);

NOR2x1_ASAP7_75t_L g1550 ( 
.A(n_1538),
.B(n_1444),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1529),
.Y(n_1551)
);

OAI31xp33_ASAP7_75t_L g1552 ( 
.A1(n_1510),
.A2(n_1545),
.A3(n_1465),
.B(n_1449),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1529),
.B(n_1498),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1541),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1535),
.B(n_1498),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1535),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1506),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1544),
.B(n_1484),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1515),
.B(n_1484),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1541),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_1522),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1512),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1528),
.B(n_1485),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1508),
.A2(n_1459),
.B1(n_1468),
.B2(n_1465),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1511),
.B(n_1485),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1542),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1534),
.B(n_1485),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1508),
.B(n_1488),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1512),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1524),
.B(n_1444),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1518),
.B(n_1498),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1518),
.B(n_1488),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1517),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1542),
.B(n_1488),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1525),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1520),
.B(n_1543),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1530),
.A2(n_1465),
.B(n_1471),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1490),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1527),
.A2(n_1468),
.B1(n_1461),
.B2(n_1463),
.Y(n_1579)
);

INVx4_ASAP7_75t_L g1580 ( 
.A(n_1520),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1507),
.B(n_1490),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1520),
.B(n_1490),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1571),
.Y(n_1583)
);

AOI222xp33_ASAP7_75t_L g1584 ( 
.A1(n_1549),
.A2(n_1461),
.B1(n_1463),
.B2(n_1464),
.C1(n_1457),
.C2(n_1519),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1551),
.B(n_1492),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1566),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1564),
.B(n_1539),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_L g1588 ( 
.A1(n_1550),
.A2(n_1523),
.B(n_1516),
.Y(n_1588)
);

AOI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1552),
.A2(n_1464),
.B1(n_1457),
.B2(n_1461),
.C(n_1463),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1575),
.Y(n_1590)
);

AOI32xp33_ASAP7_75t_L g1591 ( 
.A1(n_1550),
.A2(n_1463),
.A3(n_1461),
.B1(n_1457),
.B2(n_1464),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1556),
.B(n_1492),
.Y(n_1592)
);

AOI322xp5_ASAP7_75t_L g1593 ( 
.A1(n_1564),
.A2(n_1514),
.A3(n_1492),
.B1(n_1497),
.B2(n_1502),
.C1(n_1468),
.C2(n_1482),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1566),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1571),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1548),
.Y(n_1596)
);

AOI221xp5_ASAP7_75t_L g1597 ( 
.A1(n_1561),
.A2(n_1482),
.B1(n_1495),
.B2(n_1503),
.C(n_1547),
.Y(n_1597)
);

NOR3xp33_ASAP7_75t_L g1598 ( 
.A(n_1577),
.B(n_1547),
.C(n_1507),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1554),
.B(n_1497),
.Y(n_1599)
);

AOI21xp33_ASAP7_75t_L g1600 ( 
.A1(n_1548),
.A2(n_1521),
.B(n_1517),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1579),
.A2(n_1495),
.B1(n_1482),
.B2(n_1503),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1554),
.B(n_1553),
.Y(n_1602)
);

OAI321xp33_ASAP7_75t_L g1603 ( 
.A1(n_1579),
.A2(n_1523),
.A3(n_1516),
.B1(n_1503),
.B2(n_1495),
.C(n_1513),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1570),
.A2(n_1460),
.B1(n_1513),
.B2(n_1500),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1553),
.B(n_1497),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1558),
.B(n_1411),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1557),
.Y(n_1607)
);

INVxp67_ASAP7_75t_SL g1608 ( 
.A(n_1586),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1603),
.A2(n_1576),
.B(n_1560),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1583),
.B(n_1568),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1594),
.B(n_1555),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1606),
.B(n_1580),
.Y(n_1612)
);

AND2x2_ASAP7_75t_SL g1613 ( 
.A(n_1590),
.B(n_1580),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1595),
.B(n_1555),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1596),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1588),
.A2(n_1567),
.B1(n_1565),
.B2(n_1559),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1602),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1607),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1599),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1587),
.Y(n_1620)
);

AOI21xp33_ASAP7_75t_L g1621 ( 
.A1(n_1603),
.A2(n_1562),
.B(n_1557),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1585),
.Y(n_1622)
);

OAI31xp33_ASAP7_75t_L g1623 ( 
.A1(n_1604),
.A2(n_1581),
.A3(n_1574),
.B(n_1560),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1584),
.A2(n_1572),
.B1(n_1582),
.B2(n_1563),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1592),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1605),
.B(n_1554),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1591),
.A2(n_1578),
.B1(n_1539),
.B2(n_1572),
.Y(n_1627)
);

XNOR2xp5_ASAP7_75t_L g1628 ( 
.A(n_1614),
.B(n_1624),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1608),
.B(n_1582),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1608),
.Y(n_1630)
);

OAI321xp33_ASAP7_75t_L g1631 ( 
.A1(n_1620),
.A2(n_1589),
.A3(n_1601),
.B1(n_1597),
.B2(n_1604),
.C(n_1593),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1610),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1620),
.A2(n_1584),
.B1(n_1598),
.B2(n_1600),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1611),
.Y(n_1634)
);

INVxp33_ASAP7_75t_L g1635 ( 
.A(n_1612),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1621),
.A2(n_1573),
.B1(n_1569),
.B2(n_1562),
.C(n_1536),
.Y(n_1636)
);

OAI21xp33_ASAP7_75t_L g1637 ( 
.A1(n_1626),
.A2(n_1573),
.B(n_1569),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1629),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1630),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1634),
.B(n_1617),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1632),
.B(n_1623),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1636),
.A2(n_1609),
.B1(n_1622),
.B2(n_1625),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1628),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1636),
.B(n_1613),
.C(n_1615),
.Y(n_1644)
);

INVxp67_ASAP7_75t_L g1645 ( 
.A(n_1633),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1637),
.Y(n_1646)
);

OAI211xp5_ASAP7_75t_L g1647 ( 
.A1(n_1642),
.A2(n_1618),
.B(n_1619),
.C(n_1580),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_SL g1648 ( 
.A1(n_1642),
.A2(n_1635),
.B(n_1616),
.Y(n_1648)
);

AND4x1_ASAP7_75t_L g1649 ( 
.A(n_1640),
.B(n_1631),
.C(n_1613),
.D(n_1346),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1645),
.A2(n_1644),
.B1(n_1641),
.B2(n_1646),
.C(n_1643),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1638),
.A2(n_1627),
.B(n_1576),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_SL g1652 ( 
.A(n_1648),
.B(n_1639),
.C(n_1539),
.Y(n_1652)
);

AOI311xp33_ASAP7_75t_L g1653 ( 
.A1(n_1651),
.A2(n_1536),
.A3(n_1546),
.B(n_1521),
.C(n_1537),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1650),
.A2(n_1543),
.B(n_1537),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1647),
.A2(n_1576),
.B1(n_1543),
.B2(n_1546),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1649),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1648),
.B(n_1502),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1652),
.B(n_1346),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1656),
.B(n_1372),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1657),
.B(n_1494),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1654),
.Y(n_1661)
);

NOR2x1_ASAP7_75t_L g1662 ( 
.A(n_1655),
.B(n_1372),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1661),
.A2(n_1653),
.B1(n_1395),
.B2(n_1533),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1660),
.B(n_1526),
.Y(n_1664)
);

AOI21xp33_ASAP7_75t_SL g1665 ( 
.A1(n_1658),
.A2(n_1532),
.B(n_1531),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1664),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1666),
.Y(n_1667)
);

NAND3x1_ASAP7_75t_L g1668 ( 
.A(n_1667),
.B(n_1659),
.C(n_1662),
.Y(n_1668)
);

BUFx2_ASAP7_75t_L g1669 ( 
.A(n_1668),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1669),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1670),
.Y(n_1671)
);

AND3x4_ASAP7_75t_L g1672 ( 
.A(n_1670),
.B(n_1663),
.C(n_1665),
.Y(n_1672)
);

AOI222xp33_ASAP7_75t_L g1673 ( 
.A1(n_1671),
.A2(n_1540),
.B1(n_1398),
.B2(n_1397),
.C1(n_1501),
.C2(n_1504),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1672),
.A2(n_1500),
.B(n_1494),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1674),
.Y(n_1675)
);

XNOR2xp5_ASAP7_75t_L g1676 ( 
.A(n_1673),
.B(n_1373),
.Y(n_1676)
);

OAI221xp5_ASAP7_75t_R g1677 ( 
.A1(n_1676),
.A2(n_1479),
.B1(n_1494),
.B2(n_1500),
.C(n_1487),
.Y(n_1677)
);

AOI211xp5_ASAP7_75t_L g1678 ( 
.A1(n_1677),
.A2(n_1675),
.B(n_1368),
.C(n_1371),
.Y(n_1678)
);


endmodule