module fake_ariane_537_n_1075 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_115, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_262, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_122, n_268, n_257, n_266, n_198, n_148, n_232, n_164, n_52, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_1075);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1075;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_679;
wire n_643;
wire n_924;
wire n_927;
wire n_781;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_958;
wire n_702;
wire n_945;
wire n_905;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_398;
wire n_529;
wire n_502;
wire n_561;
wire n_821;
wire n_928;
wire n_839;
wire n_770;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_998;
wire n_999;
wire n_967;
wire n_472;
wire n_937;
wire n_296;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_394;
wire n_923;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_973;
wire n_523;
wire n_972;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_31),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_224),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_127),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_196),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_2),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_168),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_182),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_89),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_187),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_160),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_27),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_165),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_73),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_162),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_145),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_143),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_57),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_204),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_19),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_250),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_95),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_155),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_18),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_4),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_191),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_181),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_45),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_157),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_3),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_170),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_49),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_62),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_12),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_131),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_217),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_117),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_88),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_218),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_220),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_42),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_83),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_115),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_47),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_25),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_11),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_85),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_133),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_93),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_80),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_24),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_24),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_163),
.Y(n_324)
);

BUFx8_ASAP7_75t_SL g325 ( 
.A(n_112),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_192),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_138),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_75),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_100),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_199),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_180),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_248),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_166),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_142),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_270),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_328),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_287),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_310),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_314),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_280),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_314),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_325),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_302),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_294),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_322),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_274),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_323),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_289),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_283),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_272),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_271),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_273),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_275),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_315),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_287),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_310),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_300),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_276),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_277),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_329),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_305),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_278),
.B(n_0),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_279),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_281),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_287),
.B(n_0),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_288),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_349),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_343),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_344),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_344),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_341),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_346),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_348),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_355),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_338),
.B(n_287),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_350),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_360),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_358),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_359),
.Y(n_395)
);

BUFx12f_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_356),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_362),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_366),
.Y(n_402)
);

NAND2x1_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_287),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_366),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_352),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_340),
.A2(n_284),
.B1(n_285),
.B2(n_282),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_370),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

BUFx8_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_376),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_372),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_376),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_368),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_339),
.B(n_290),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_337),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_379),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_368),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_397),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_379),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_335),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_388),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_397),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_379),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_409),
.B(n_335),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_390),
.A2(n_374),
.B1(n_342),
.B2(n_340),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_426),
.B(n_287),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_423),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_379),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_291),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_399),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_399),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_392),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_SL g446 ( 
.A(n_402),
.B(n_342),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_389),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_426),
.B(n_333),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_399),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_399),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_390),
.A2(n_333),
.B1(n_298),
.B2(n_301),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_295),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_407),
.B(n_304),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_407),
.B(n_306),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_378),
.B(n_307),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_426),
.B(n_333),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_420),
.B(n_308),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_381),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_398),
.B(n_309),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_426),
.B(n_333),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_390),
.A2(n_333),
.B1(n_312),
.B2(n_313),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_386),
.Y(n_471)
);

INVx4_ASAP7_75t_SL g472 ( 
.A(n_390),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_401),
.B(n_311),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

NAND3xp33_ASAP7_75t_L g476 ( 
.A(n_395),
.B(n_318),
.C(n_317),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_408),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_411),
.B(n_320),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_412),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_413),
.B(n_321),
.Y(n_480)
);

INVx4_ASAP7_75t_SL g481 ( 
.A(n_417),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_406),
.B(n_333),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_396),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_387),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_380),
.B(n_324),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_410),
.A2(n_327),
.B1(n_331),
.B2(n_326),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_1),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_418),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_380),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_404),
.B(n_4),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_415),
.Y(n_494)
);

BUFx8_ASAP7_75t_L g495 ( 
.A(n_445),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_475),
.Y(n_496)
);

BUFx12f_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_431),
.B(n_414),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_437),
.B(n_414),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_429),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_485),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_459),
.A2(n_391),
.B1(n_383),
.B2(n_382),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_428),
.B(n_5),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_458),
.B(n_5),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_492),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_473),
.B(n_6),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_461),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

BUFx8_ASAP7_75t_L g509 ( 
.A(n_463),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_468),
.B(n_6),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_473),
.B(n_442),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_475),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_442),
.B(n_7),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_433),
.B(n_7),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_463),
.B(n_8),
.Y(n_515)
);

AND2x6_ASAP7_75t_SL g516 ( 
.A(n_488),
.B(n_8),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_492),
.B(n_9),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_9),
.Y(n_518)
);

BUFx12f_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_486),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_447),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_433),
.B(n_10),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_490),
.B(n_10),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_487),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_456),
.B(n_13),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_479),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_457),
.B(n_479),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_14),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_436),
.B(n_14),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_471),
.B(n_15),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_15),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_464),
.B(n_16),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_477),
.B(n_16),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_464),
.B(n_17),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_484),
.B(n_17),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_483),
.B(n_477),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_483),
.B(n_18),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_441),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_482),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_447),
.B(n_19),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_427),
.B(n_430),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_432),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_427),
.B(n_20),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_487),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_447),
.B(n_21),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_440),
.B(n_22),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_430),
.B(n_23),
.Y(n_549)
);

AND2x6_ASAP7_75t_SL g550 ( 
.A(n_491),
.B(n_23),
.Y(n_550)
);

NOR2x1p5_ASAP7_75t_L g551 ( 
.A(n_484),
.B(n_25),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_440),
.B(n_26),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_443),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_438),
.B(n_26),
.Y(n_554)
);

OR2x6_ASAP7_75t_L g555 ( 
.A(n_448),
.B(n_27),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_443),
.B(n_28),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_444),
.Y(n_558)
);

O2A1O1Ixp33_ASAP7_75t_L g559 ( 
.A1(n_466),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_480),
.B(n_455),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_L g561 ( 
.A(n_448),
.B(n_35),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_480),
.B(n_29),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_450),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_450),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_453),
.A2(n_470),
.B1(n_449),
.B2(n_460),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_511),
.A2(n_449),
.B(n_439),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_560),
.B(n_438),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_494),
.B(n_454),
.Y(n_568)
);

OR2x6_ASAP7_75t_SL g569 ( 
.A(n_525),
.B(n_446),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_529),
.A2(n_543),
.B(n_526),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

O2A1O1Ixp33_ASAP7_75t_L g572 ( 
.A1(n_525),
.A2(n_478),
.B(n_474),
.C(n_460),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_543),
.A2(n_467),
.B(n_439),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_503),
.B(n_454),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_500),
.A2(n_467),
.B(n_452),
.Y(n_575)
);

O2A1O1Ixp33_ASAP7_75t_SL g576 ( 
.A1(n_562),
.A2(n_513),
.B(n_506),
.C(n_504),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_508),
.A2(n_452),
.B(n_451),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_505),
.B(n_544),
.Y(n_578)
);

OAI21xp33_ASAP7_75t_L g579 ( 
.A1(n_510),
.A2(n_489),
.B(n_476),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_554),
.B(n_469),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_L g581 ( 
.A(n_542),
.B(n_446),
.C(n_469),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_507),
.A2(n_452),
.B(n_451),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_520),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_521),
.A2(n_565),
.B1(n_546),
.B2(n_538),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_539),
.A2(n_452),
.B(n_434),
.Y(n_585)
);

AO21x2_ASAP7_75t_L g586 ( 
.A1(n_545),
.A2(n_434),
.B(n_481),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_496),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_539),
.A2(n_434),
.B(n_461),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_501),
.B(n_461),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_512),
.Y(n_590)
);

O2A1O1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_534),
.A2(n_470),
.B(n_453),
.C(n_32),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_553),
.A2(n_434),
.B(n_461),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_558),
.A2(n_472),
.B(n_481),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_522),
.B(n_481),
.Y(n_594)
);

OAI21x1_ASAP7_75t_L g595 ( 
.A1(n_557),
.A2(n_472),
.B(n_37),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_527),
.B(n_472),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_517),
.B(n_30),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_520),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_563),
.A2(n_38),
.B(n_36),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_564),
.A2(n_40),
.B(n_39),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_545),
.A2(n_43),
.B(n_41),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_502),
.B(n_31),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_498),
.B(n_32),
.Y(n_604)
);

BUFx8_ASAP7_75t_SL g605 ( 
.A(n_497),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_515),
.B(n_33),
.Y(n_606)
);

NOR2x1p5_ASAP7_75t_L g607 ( 
.A(n_519),
.B(n_33),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_549),
.A2(n_46),
.B(n_44),
.Y(n_608)
);

CKINVDCx6p67_ASAP7_75t_R g609 ( 
.A(n_537),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_499),
.B(n_551),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_549),
.A2(n_50),
.B(n_48),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_524),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_528),
.Y(n_613)
);

OA22x2_ASAP7_75t_L g614 ( 
.A1(n_537),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_547),
.B(n_34),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_555),
.B(n_53),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_518),
.B(n_54),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_495),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_L g619 ( 
.A(n_533),
.B(n_55),
.C(n_56),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_535),
.B(n_495),
.Y(n_620)
);

O2A1O1Ixp33_ASAP7_75t_L g621 ( 
.A1(n_536),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_509),
.B(n_61),
.Y(n_622)
);

CKINVDCx10_ASAP7_75t_R g623 ( 
.A(n_537),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_556),
.A2(n_63),
.B(n_64),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_556),
.A2(n_65),
.B(n_66),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_555),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_514),
.A2(n_523),
.B(n_532),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_535),
.B(n_67),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_612),
.B(n_555),
.Y(n_629)
);

OA22x2_ASAP7_75t_L g630 ( 
.A1(n_610),
.A2(n_530),
.B1(n_531),
.B2(n_509),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_574),
.A2(n_531),
.B(n_530),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_618),
.Y(n_632)
);

OA22x2_ASAP7_75t_L g633 ( 
.A1(n_610),
.A2(n_552),
.B1(n_548),
.B2(n_516),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_570),
.A2(n_576),
.B(n_627),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_566),
.A2(n_561),
.B(n_559),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_584),
.A2(n_550),
.B1(n_69),
.B2(n_70),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_567),
.B(n_68),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_571),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_572),
.A2(n_71),
.B(n_72),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_595),
.A2(n_74),
.B(n_76),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_580),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_R g642 ( 
.A(n_623),
.B(n_77),
.Y(n_642)
);

A2O1A1Ixp33_ASAP7_75t_L g643 ( 
.A1(n_579),
.A2(n_78),
.B(n_79),
.C(n_81),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_587),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_573),
.A2(n_82),
.B(n_84),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_585),
.A2(n_86),
.B(n_87),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_603),
.B(n_90),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_L g648 ( 
.A1(n_591),
.A2(n_91),
.B(n_92),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_568),
.A2(n_94),
.B(n_96),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_599),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_589),
.B(n_97),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_578),
.B(n_98),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_597),
.A2(n_99),
.B(n_101),
.C(n_102),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_616),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_569),
.B(n_106),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_626),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_590),
.B(n_107),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_581),
.B(n_108),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_626),
.B(n_606),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_626),
.B(n_109),
.Y(n_661)
);

OAI21x1_ASAP7_75t_SL g662 ( 
.A1(n_621),
.A2(n_110),
.B(n_111),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_583),
.B(n_113),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_588),
.A2(n_114),
.B(n_116),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_592),
.A2(n_118),
.B(n_119),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_620),
.B(n_120),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_619),
.B(n_121),
.C(n_122),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_613),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_593),
.A2(n_123),
.B(n_124),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_599),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_616),
.B(n_125),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_583),
.B(n_126),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_598),
.B(n_128),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_599),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_L g675 ( 
.A1(n_617),
.A2(n_129),
.B(n_130),
.C(n_132),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_598),
.B(n_134),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_575),
.A2(n_135),
.B(n_136),
.C(n_137),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_609),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_615),
.B(n_139),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_605),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_622),
.Y(n_681)
);

BUFx2_ASAP7_75t_SL g682 ( 
.A(n_614),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_594),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_577),
.A2(n_140),
.B(n_141),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_607),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_596),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_628),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_602),
.A2(n_148),
.B(n_149),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_658),
.B(n_582),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_681),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_636),
.A2(n_625),
.B1(n_624),
.B2(n_611),
.Y(n_691)
);

BUFx12f_ASAP7_75t_L g692 ( 
.A(n_678),
.Y(n_692)
);

INVx3_ASAP7_75t_SL g693 ( 
.A(n_680),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_631),
.A2(n_608),
.B(n_601),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_656),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_644),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_634),
.A2(n_586),
.B(n_600),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_641),
.B(n_682),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_629),
.B(n_586),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_687),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_700)
);

NAND2x1_ASAP7_75t_L g701 ( 
.A(n_650),
.B(n_153),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_641),
.B(n_269),
.Y(n_702)
);

OAI221xp5_ASAP7_75t_L g703 ( 
.A1(n_636),
.A2(n_648),
.B1(n_655),
.B2(n_633),
.C(n_654),
.Y(n_703)
);

O2A1O1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_648),
.A2(n_154),
.B(n_156),
.C(n_158),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_640),
.A2(n_159),
.B(n_161),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_681),
.B(n_268),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_635),
.A2(n_164),
.B(n_167),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_668),
.Y(n_708)
);

O2A1O1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_671),
.A2(n_169),
.B(n_171),
.C(n_172),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_638),
.B(n_267),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_660),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_647),
.B(n_173),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_657),
.Y(n_713)
);

BUFx12f_ASAP7_75t_L g714 ( 
.A(n_681),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_637),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_670),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_666),
.B(n_266),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_632),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_650),
.B(n_174),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_664),
.A2(n_175),
.B(n_176),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_666),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_674),
.B(n_183),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_630),
.B(n_265),
.Y(n_723)
);

O2A1O1Ixp33_ASAP7_75t_SL g724 ( 
.A1(n_659),
.A2(n_184),
.B(n_185),
.C(n_186),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_639),
.A2(n_651),
.B(n_645),
.Y(n_725)
);

AOI21xp33_ASAP7_75t_L g726 ( 
.A1(n_652),
.A2(n_188),
.B(n_189),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_654),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_683),
.B(n_195),
.Y(n_728)
);

AO22x1_ASAP7_75t_L g729 ( 
.A1(n_685),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_729)
);

INVx5_ASAP7_75t_L g730 ( 
.A(n_683),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_683),
.B(n_201),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_642),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_661),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_679),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_663),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_669),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_672),
.B(n_264),
.Y(n_737)
);

CKINVDCx8_ASAP7_75t_R g738 ( 
.A(n_662),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_673),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_684),
.B(n_202),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_676),
.A2(n_649),
.B(n_684),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_686),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_699),
.B(n_643),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_703),
.A2(n_667),
.B1(n_653),
.B2(n_677),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_718),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_717),
.A2(n_667),
.B1(n_646),
.B2(n_688),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_698),
.B(n_665),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_696),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_730),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_730),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_708),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_711),
.B(n_203),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_695),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_716),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_730),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_689),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_717),
.B(n_715),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_733),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_740),
.A2(n_675),
.B1(n_206),
.B2(n_208),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_715),
.B(n_205),
.Y(n_760)
);

AOI21x1_ASAP7_75t_L g761 ( 
.A1(n_741),
.A2(n_697),
.B(n_725),
.Y(n_761)
);

AO21x1_ASAP7_75t_L g762 ( 
.A1(n_704),
.A2(n_263),
.B(n_210),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_710),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_690),
.B(n_262),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_727),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_714),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_742),
.A2(n_213),
.B(n_214),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_690),
.Y(n_768)
);

OA21x2_ASAP7_75t_L g769 ( 
.A1(n_694),
.A2(n_215),
.B(n_216),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_690),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_732),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_736),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_734),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_702),
.Y(n_774)
);

OAI21x1_ASAP7_75t_L g775 ( 
.A1(n_707),
.A2(n_219),
.B(n_221),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_735),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_719),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_736),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_723),
.A2(n_261),
.B1(n_223),
.B2(n_225),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_736),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_738),
.Y(n_781)
);

INVx6_ASAP7_75t_L g782 ( 
.A(n_692),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_713),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_713),
.A2(n_222),
.B(n_226),
.Y(n_784)
);

OAI21x1_ASAP7_75t_L g785 ( 
.A1(n_720),
.A2(n_227),
.B(n_228),
.Y(n_785)
);

AOI21x1_ASAP7_75t_L g786 ( 
.A1(n_739),
.A2(n_229),
.B(n_230),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_712),
.A2(n_231),
.B(n_232),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_722),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_705),
.A2(n_701),
.B(n_709),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_722),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

CKINVDCx11_ASAP7_75t_R g792 ( 
.A(n_693),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_728),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_737),
.Y(n_794)
);

AOI222xp33_ASAP7_75t_L g795 ( 
.A1(n_700),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.C1(n_236),
.C2(n_237),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_706),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_728),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_737),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_721),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_756),
.B(n_729),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_783),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_776),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_758),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_772),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_772),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_778),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_778),
.Y(n_807)
);

AO21x2_ASAP7_75t_L g808 ( 
.A1(n_761),
.A2(n_744),
.B(n_780),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_780),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_773),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_748),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_751),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_754),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_791),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_769),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_781),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_799),
.A2(n_691),
.B(n_724),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_769),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_757),
.B(n_726),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_777),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_757),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_798),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_743),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_743),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_781),
.Y(n_825)
);

CKINVDCx6p67_ASAP7_75t_R g826 ( 
.A(n_792),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_781),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_769),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_794),
.B(n_238),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_763),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_794),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_794),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_774),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_788),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_753),
.B(n_239),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_747),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_789),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_790),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_799),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_768),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_745),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_799),
.A2(n_240),
.B(n_241),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_760),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_797),
.B(n_242),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_768),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_760),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_786),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_793),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_814),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_821),
.B(n_823),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_821),
.B(n_749),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_817),
.B(n_779),
.C(n_795),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_823),
.B(n_749),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_824),
.B(n_796),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_L g855 ( 
.A(n_836),
.B(n_779),
.C(n_784),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_802),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_810),
.B(n_752),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_814),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_831),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_820),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_839),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_836),
.B(n_752),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_801),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_801),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_830),
.B(n_755),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_839),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_833),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_840),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_833),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_808),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_811),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_822),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_800),
.B(n_768),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_831),
.B(n_746),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_825),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_803),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_803),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_811),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_812),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_830),
.Y(n_880)
);

AOI221xp5_ASAP7_75t_L g881 ( 
.A1(n_800),
.A2(n_762),
.B1(n_759),
.B2(n_746),
.C(n_766),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_812),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_813),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_831),
.B(n_767),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_841),
.B(n_750),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_816),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_831),
.B(n_759),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_832),
.B(n_785),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_813),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_832),
.B(n_785),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_832),
.B(n_792),
.Y(n_891)
);

OR2x2_ASAP7_75t_SL g892 ( 
.A(n_843),
.B(n_782),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_825),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_848),
.Y(n_894)
);

NAND4xp25_ASAP7_75t_L g895 ( 
.A(n_852),
.B(n_835),
.C(n_825),
.D(n_837),
.Y(n_895)
);

OAI221xp5_ASAP7_75t_SL g896 ( 
.A1(n_881),
.A2(n_843),
.B1(n_819),
.B2(n_826),
.C(n_765),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_856),
.B(n_819),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_891),
.B(n_826),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_872),
.B(n_827),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_860),
.B(n_827),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_SL g901 ( 
.A(n_855),
.B(n_842),
.C(n_844),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_850),
.B(n_862),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_850),
.B(n_816),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_891),
.B(n_832),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_887),
.A2(n_838),
.B1(n_846),
.B2(n_848),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_849),
.B(n_846),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_851),
.B(n_853),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_L g908 ( 
.A1(n_870),
.A2(n_838),
.B1(n_818),
.B2(n_815),
.C(n_828),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_849),
.B(n_808),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_SL g910 ( 
.A1(n_887),
.A2(n_844),
.B(n_837),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_866),
.B(n_809),
.C(n_805),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_858),
.B(n_808),
.Y(n_912)
);

NAND4xp25_ASAP7_75t_SL g913 ( 
.A(n_874),
.B(n_782),
.C(n_829),
.D(n_815),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_858),
.B(n_807),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_867),
.B(n_807),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_SL g916 ( 
.A1(n_892),
.A2(n_782),
.B1(n_771),
.B2(n_844),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_867),
.B(n_809),
.Y(n_917)
);

OAI221xp5_ASAP7_75t_SL g918 ( 
.A1(n_857),
.A2(n_828),
.B1(n_818),
.B2(n_847),
.C(n_829),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_851),
.B(n_806),
.Y(n_919)
);

OA21x2_ASAP7_75t_L g920 ( 
.A1(n_870),
.A2(n_847),
.B(n_805),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_892),
.A2(n_885),
.B1(n_851),
.B2(n_886),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_853),
.B(n_806),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_869),
.B(n_806),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_869),
.B(n_806),
.Y(n_924)
);

OA21x2_ASAP7_75t_L g925 ( 
.A1(n_873),
.A2(n_804),
.B(n_834),
.Y(n_925)
);

NOR3xp33_ASAP7_75t_L g926 ( 
.A(n_865),
.B(n_787),
.C(n_837),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_853),
.B(n_845),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_L g928 ( 
.A(n_874),
.B(n_837),
.C(n_775),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_861),
.A2(n_845),
.B1(n_840),
.B2(n_750),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_861),
.A2(n_845),
.B1(n_840),
.B2(n_755),
.Y(n_930)
);

NAND3xp33_ASAP7_75t_L g931 ( 
.A(n_880),
.B(n_804),
.C(n_840),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_897),
.Y(n_932)
);

AND2x2_ASAP7_75t_SL g933 ( 
.A(n_928),
.B(n_868),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_907),
.B(n_893),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_919),
.B(n_922),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_920),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_914),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_899),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_928),
.B(n_875),
.Y(n_939)
);

BUFx2_ASAP7_75t_SL g940 ( 
.A(n_898),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_920),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_927),
.B(n_893),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_904),
.B(n_875),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_915),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_902),
.B(n_859),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_923),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_917),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_924),
.B(n_880),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_903),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_906),
.B(n_900),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_911),
.B(n_859),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_921),
.B(n_859),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_909),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_925),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_931),
.B(n_926),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_910),
.B(n_890),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_952),
.B(n_926),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_954),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_932),
.B(n_937),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_937),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_952),
.B(n_930),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_940),
.B(n_929),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_944),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_939),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_944),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_940),
.B(n_868),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_947),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_947),
.B(n_877),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_938),
.B(n_895),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_948),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_950),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_969),
.B(n_950),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_971),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_964),
.B(n_955),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_970),
.B(n_946),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_961),
.B(n_935),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_958),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_959),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_961),
.B(n_935),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_962),
.B(n_945),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_968),
.Y(n_981)
);

NAND2x1_ASAP7_75t_L g982 ( 
.A(n_964),
.B(n_951),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_957),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_969),
.B(n_949),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_983),
.B(n_957),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_972),
.B(n_960),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_973),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_972),
.B(n_963),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_975),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_978),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_984),
.B(n_965),
.Y(n_991)
);

OAI22xp33_ASAP7_75t_L g992 ( 
.A1(n_991),
.A2(n_974),
.B1(n_984),
.B2(n_901),
.Y(n_992)
);

AOI322xp5_ASAP7_75t_L g993 ( 
.A1(n_985),
.A2(n_990),
.A3(n_988),
.B1(n_986),
.B2(n_989),
.C1(n_987),
.C2(n_936),
.Y(n_993)
);

NOR4xp25_ASAP7_75t_SL g994 ( 
.A(n_989),
.B(n_896),
.C(n_981),
.D(n_982),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_985),
.B(n_976),
.Y(n_995)
);

INVxp67_ASAP7_75t_SL g996 ( 
.A(n_985),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_996),
.B(n_995),
.Y(n_997)
);

AOI222xp33_ASAP7_75t_L g998 ( 
.A1(n_992),
.A2(n_977),
.B1(n_936),
.B2(n_941),
.C1(n_958),
.C2(n_955),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_994),
.Y(n_999)
);

OAI221xp5_ASAP7_75t_SL g1000 ( 
.A1(n_993),
.A2(n_964),
.B1(n_936),
.B2(n_941),
.C(n_980),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_995),
.B(n_979),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_SL g1002 ( 
.A(n_997),
.B(n_771),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_998),
.B(n_1001),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_999),
.B(n_967),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_1000),
.B(n_955),
.Y(n_1005)
);

NAND4xp75_ASAP7_75t_L g1006 ( 
.A(n_999),
.B(n_933),
.C(n_977),
.D(n_956),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_997),
.B(n_933),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_999),
.A2(n_896),
.B(n_901),
.C(n_918),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_L g1009 ( 
.A(n_1004),
.B(n_933),
.C(n_766),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_1003),
.B(n_953),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_1002),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_L g1012 ( 
.A(n_1006),
.B(n_766),
.Y(n_1012)
);

AOI211x1_ASAP7_75t_L g1013 ( 
.A1(n_1005),
.A2(n_966),
.B(n_956),
.C(n_913),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_1007),
.B(n_945),
.Y(n_1014)
);

OAI211xp5_ASAP7_75t_L g1015 ( 
.A1(n_1011),
.A2(n_1008),
.B(n_766),
.C(n_934),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1010),
.B(n_953),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1014),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_SL g1018 ( 
.A(n_1009),
.B(n_764),
.C(n_954),
.Y(n_1018)
);

AOI211xp5_ASAP7_75t_L g1019 ( 
.A1(n_1012),
.A2(n_916),
.B(n_939),
.C(n_918),
.Y(n_1019)
);

NOR3x1_ASAP7_75t_L g1020 ( 
.A(n_1013),
.B(n_770),
.C(n_789),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_1011),
.B(n_951),
.Y(n_1021)
);

OAI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_1012),
.A2(n_912),
.B1(n_908),
.B2(n_905),
.C(n_883),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_1015),
.A2(n_939),
.B1(n_951),
.B2(n_884),
.Y(n_1023)
);

NOR2xp67_ASAP7_75t_L g1024 ( 
.A(n_1017),
.B(n_939),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1016),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1021),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1020),
.Y(n_1027)
);

NOR3xp33_ASAP7_75t_L g1028 ( 
.A(n_1018),
.B(n_770),
.C(n_775),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1022),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1019),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1016),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1016),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1015),
.A2(n_884),
.B1(n_934),
.B2(n_942),
.Y(n_1033)
);

AO22x2_ASAP7_75t_L g1034 ( 
.A1(n_1017),
.A2(n_943),
.B1(n_942),
.B2(n_868),
.Y(n_1034)
);

AOI211xp5_ASAP7_75t_L g1035 ( 
.A1(n_1024),
.A2(n_768),
.B(n_890),
.C(n_888),
.Y(n_1035)
);

OAI211xp5_ASAP7_75t_SL g1036 ( 
.A1(n_1025),
.A2(n_1031),
.B(n_1032),
.C(n_1030),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_1026),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_1034),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1027),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1029),
.B(n_883),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1028),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1033),
.B(n_876),
.Y(n_1042)
);

NAND4xp75_ASAP7_75t_L g1043 ( 
.A(n_1023),
.B(n_943),
.C(n_925),
.D(n_877),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1025),
.B(n_876),
.Y(n_1044)
);

OR2x2_ASAP7_75t_L g1045 ( 
.A(n_1025),
.B(n_894),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1025),
.B(n_894),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1026),
.B(n_889),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1026),
.B(n_889),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1037),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1044),
.Y(n_1050)
);

NAND2xp33_ASAP7_75t_L g1051 ( 
.A(n_1038),
.B(n_840),
.Y(n_1051)
);

NOR2x1_ASAP7_75t_L g1052 ( 
.A(n_1036),
.B(n_888),
.Y(n_1052)
);

NAND3x1_ASAP7_75t_L g1053 ( 
.A(n_1041),
.B(n_864),
.C(n_863),
.Y(n_1053)
);

INVx2_ASAP7_75t_SL g1054 ( 
.A(n_1045),
.Y(n_1054)
);

XOR2x1_ASAP7_75t_SL g1055 ( 
.A(n_1039),
.B(n_882),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_854),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1049),
.Y(n_1057)
);

XOR2xp5_ASAP7_75t_L g1058 ( 
.A(n_1050),
.B(n_1040),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1054),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1053),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_1051),
.A2(n_1052),
.B1(n_1043),
.B2(n_1055),
.Y(n_1061)
);

O2A1O1Ixp5_ASAP7_75t_L g1062 ( 
.A1(n_1059),
.A2(n_1042),
.B(n_1048),
.C(n_1047),
.Y(n_1062)
);

XNOR2xp5_ASAP7_75t_L g1063 ( 
.A(n_1058),
.B(n_1056),
.Y(n_1063)
);

XNOR2xp5_ASAP7_75t_L g1064 ( 
.A(n_1057),
.B(n_1035),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_SL g1065 ( 
.A(n_1061),
.B(n_854),
.C(n_879),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_1060),
.B1(n_879),
.B2(n_882),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1066),
.A2(n_1063),
.B1(n_1062),
.B2(n_1065),
.Y(n_1067)
);

OA21x2_ASAP7_75t_L g1068 ( 
.A1(n_1066),
.A2(n_878),
.B(n_871),
.Y(n_1068)
);

AOI22x1_ASAP7_75t_L g1069 ( 
.A1(n_1067),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_247),
.Y(n_1070)
);

AOI22x1_ASAP7_75t_L g1071 ( 
.A1(n_1069),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1070),
.B(n_253),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1071),
.A2(n_878),
.B1(n_871),
.B2(n_864),
.Y(n_1073)
);

OAI221xp5_ASAP7_75t_R g1074 ( 
.A1(n_1073),
.A2(n_1072),
.B1(n_255),
.B2(n_256),
.C(n_258),
.Y(n_1074)
);

AOI211xp5_ASAP7_75t_L g1075 ( 
.A1(n_1074),
.A2(n_254),
.B(n_259),
.C(n_260),
.Y(n_1075)
);


endmodule