module fake_ibex_1975_n_992 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_992);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_992;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_317;
wire n_340;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_496;
wire n_301;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_980;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_858;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_444;
wire n_200;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_440;
wire n_268;
wire n_955;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_912;
wire n_921;
wire n_890;
wire n_874;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_62),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_72),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_66),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_49),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_174),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_35),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_L g192 ( 
.A(n_48),
.B(n_175),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_13),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_68),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_32),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_109),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_70),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_43),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_74),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_89),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_53),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_78),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_148),
.Y(n_208)
);

BUFx2_ASAP7_75t_SL g209 ( 
.A(n_32),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_5),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_31),
.Y(n_213)
);

NOR2xp67_ASAP7_75t_L g214 ( 
.A(n_28),
.B(n_46),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_28),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_126),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_20),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_130),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_22),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_91),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_86),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_58),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_154),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_16),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_59),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_25),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_116),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_33),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_75),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_23),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_69),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_128),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_167),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_82),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_123),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_83),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_117),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_98),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_14),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_100),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_50),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_131),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_L g251 ( 
.A(n_122),
.B(n_108),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_60),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_87),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_67),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_169),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_97),
.Y(n_256)
);

NOR2xp67_ASAP7_75t_L g257 ( 
.A(n_146),
.B(n_119),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_51),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_25),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_162),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_84),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_56),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_81),
.Y(n_263)
);

HB1xp67_ASAP7_75t_SL g264 ( 
.A(n_1),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_115),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_106),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_101),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_80),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_42),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_141),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_54),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_111),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_158),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_9),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_143),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_163),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_71),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_61),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_33),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_57),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_145),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_135),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_164),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_121),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_4),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_107),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_177),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_124),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_40),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_21),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_19),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_73),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_150),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_36),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_105),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_120),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_1),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_99),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_55),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_103),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_190),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_197),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_241),
.B(n_0),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_193),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_199),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_199),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_193),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_197),
.B(n_0),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_178),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_250),
.B(n_2),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_181),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_213),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_181),
.Y(n_315)
);

BUFx8_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_226),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_202),
.A2(n_242),
.B(n_231),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_202),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_231),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_265),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_250),
.B(n_2),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_269),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_230),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_242),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_179),
.Y(n_331)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_254),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_248),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_270),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_264),
.B(n_3),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_182),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_180),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_186),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_213),
.Y(n_341)
);

OA21x2_ASAP7_75t_L g342 ( 
.A1(n_267),
.A2(n_76),
.B(n_173),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_277),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_187),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_191),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_194),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_213),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_196),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_283),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_201),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_255),
.B(n_280),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_6),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_203),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_280),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_200),
.Y(n_357)
);

CKINVDCx6p67_ASAP7_75t_R g358 ( 
.A(n_183),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_213),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_291),
.B(n_6),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_183),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_205),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_215),
.Y(n_363)
);

AND2x6_ASAP7_75t_L g364 ( 
.A(n_206),
.B(n_44),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_212),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_182),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_218),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_219),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_220),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_292),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_222),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_224),
.Y(n_373)
);

BUFx8_ASAP7_75t_SL g374 ( 
.A(n_230),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_217),
.B(n_7),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_229),
.A2(n_77),
.B(n_171),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_337),
.B(n_184),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_332),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_316),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_375),
.A2(n_228),
.B1(n_235),
.B2(n_290),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_332),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_332),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_185),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_232),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_326),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_339),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_332),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_366),
.B(n_185),
.Y(n_393)
);

CKINVDCx6p67_ASAP7_75t_R g394 ( 
.A(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_SL g396 ( 
.A(n_323),
.B(n_204),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_188),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_SL g399 ( 
.A(n_323),
.B(n_204),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

NAND3xp33_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_233),
.C(n_210),
.Y(n_403)
);

BUFx8_ASAP7_75t_SL g404 ( 
.A(n_374),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_311),
.A2(n_236),
.B(n_234),
.Y(n_405)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_350),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_323),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_375),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_306),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_188),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_306),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_371),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_375),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_305),
.Y(n_416)
);

BUFx10_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_353),
.B(n_189),
.Y(n_418)
);

NAND2xp33_ASAP7_75t_L g419 ( 
.A(n_364),
.B(n_198),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_373),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_306),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_333),
.B(n_309),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_357),
.B(n_316),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_333),
.B(n_292),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_357),
.B(n_271),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_271),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_365),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_365),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_373),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_373),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_307),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_307),
.Y(n_433)
);

NAND2xp33_ASAP7_75t_SL g434 ( 
.A(n_317),
.B(n_223),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_307),
.Y(n_435)
);

OAI22xp33_ASAP7_75t_L g436 ( 
.A1(n_335),
.A2(n_275),
.B1(n_195),
.B2(n_282),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_307),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_307),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_303),
.Y(n_440)
);

AO21x2_ASAP7_75t_L g441 ( 
.A1(n_360),
.A2(n_238),
.B(n_237),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

INVx2_ASAP7_75t_SL g443 ( 
.A(n_325),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_364),
.A2(n_298),
.B1(n_221),
.B2(n_286),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_311),
.B(n_273),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_303),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_308),
.Y(n_448)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

BUFx8_ASAP7_75t_SL g450 ( 
.A(n_302),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_331),
.B(n_338),
.Y(n_451)
);

OA22x2_ASAP7_75t_L g452 ( 
.A1(n_335),
.A2(n_209),
.B1(n_259),
.B2(n_246),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_331),
.B(n_274),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_313),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_318),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_338),
.B(n_281),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

OAI21xp33_ASAP7_75t_SL g458 ( 
.A1(n_340),
.A2(n_214),
.B(n_240),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_340),
.B(n_281),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_344),
.B(n_289),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_317),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_313),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_318),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_327),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_328),
.B(n_370),
.Y(n_465)
);

INVx8_ASAP7_75t_L g466 ( 
.A(n_406),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_406),
.A2(n_364),
.B1(n_372),
.B2(n_369),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_344),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_345),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_345),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_346),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_346),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_454),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_349),
.Y(n_475)
);

AND2x2_ASAP7_75t_SL g476 ( 
.A(n_416),
.B(n_358),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_441),
.B(n_349),
.Y(n_477)
);

INVx4_ASAP7_75t_L g478 ( 
.A(n_406),
.Y(n_478)
);

OAI221xp5_ASAP7_75t_L g479 ( 
.A1(n_383),
.A2(n_304),
.B1(n_372),
.B2(n_369),
.C(n_352),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_465),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_425),
.B(n_358),
.Y(n_481)
);

BUFx5_ASAP7_75t_L g482 ( 
.A(n_377),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_387),
.B(n_352),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_430),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_430),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_430),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_R g487 ( 
.A(n_382),
.B(n_361),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_398),
.B(n_367),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_465),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_431),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_464),
.B(n_394),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_411),
.B(n_367),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_L g495 ( 
.A1(n_452),
.A2(n_361),
.B1(n_275),
.B2(n_282),
.Y(n_495)
);

OA22x2_ASAP7_75t_L g496 ( 
.A1(n_425),
.A2(n_336),
.B1(n_368),
.B2(n_355),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_423),
.B(n_336),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_440),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_423),
.B(n_443),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_441),
.B(n_312),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_443),
.B(n_295),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_449),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_426),
.B(n_362),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_406),
.A2(n_368),
.B1(n_310),
.B2(n_322),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_424),
.B(n_310),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_452),
.A2(n_223),
.B1(n_315),
.B2(n_351),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_427),
.B(n_296),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_400),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_403),
.B(n_378),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_446),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_400),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_393),
.B(n_207),
.Y(n_513)
);

INVx8_ASAP7_75t_L g514 ( 
.A(n_449),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_414),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_397),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_453),
.B(n_456),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_452),
.A2(n_320),
.B1(n_334),
.B2(n_351),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_380),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_382),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_459),
.B(n_208),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_401),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_402),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_420),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_428),
.B(n_211),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_434),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_428),
.B(n_216),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_409),
.B(n_321),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_436),
.B(n_329),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_412),
.A2(n_329),
.B1(n_334),
.B2(n_343),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_429),
.B(n_225),
.Y(n_533)
);

AOI221xp5_ASAP7_75t_L g534 ( 
.A1(n_396),
.A2(n_347),
.B1(n_343),
.B2(n_294),
.C(n_243),
.Y(n_534)
);

NOR3xp33_ASAP7_75t_L g535 ( 
.A(n_399),
.B(n_247),
.C(n_245),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_415),
.B(n_347),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_451),
.B(n_408),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_429),
.B(n_342),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_379),
.B(n_227),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_461),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_384),
.B(n_239),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_414),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_377),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_397),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_449),
.B(n_244),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_386),
.B(n_249),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_399),
.A2(n_322),
.B1(n_324),
.B2(n_342),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_386),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_392),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_405),
.B(n_253),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_466),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_466),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_480),
.A2(n_490),
.B1(n_535),
.B2(n_466),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_472),
.B(n_388),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_538),
.A2(n_419),
.B(n_457),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_L g556 ( 
.A(n_540),
.B(n_458),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_538),
.A2(n_419),
.B(n_457),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_468),
.B(n_417),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_470),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_508),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_543),
.A2(n_457),
.B(n_447),
.Y(n_561)
);

AO21x1_ASAP7_75t_L g562 ( 
.A1(n_500),
.A2(n_438),
.B(n_421),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_478),
.A2(n_537),
.B1(n_499),
.B2(n_477),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_500),
.A2(n_447),
.B(n_444),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_469),
.B(n_417),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_534),
.B(n_417),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_502),
.B(n_447),
.Y(n_567)
);

OAI21xp33_ASAP7_75t_L g568 ( 
.A1(n_501),
.A2(n_461),
.B(n_392),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_496),
.A2(n_278),
.B1(n_279),
.B2(n_284),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_494),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_SL g571 ( 
.A(n_478),
.B(n_252),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_483),
.A2(n_376),
.B(n_381),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_488),
.A2(n_376),
.B(n_381),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_493),
.A2(n_376),
.B(n_395),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_502),
.B(n_256),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_471),
.B(n_260),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_471),
.B(n_262),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_503),
.A2(n_477),
.B(n_475),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_502),
.B(n_266),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_517),
.B(n_297),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_487),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_514),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_492),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_515),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_467),
.A2(n_300),
.B1(n_258),
.B2(n_261),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_479),
.A2(n_288),
.B1(n_293),
.B2(n_287),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_544),
.B(n_299),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_514),
.Y(n_588)
);

NOR2x1_ASAP7_75t_L g589 ( 
.A(n_481),
.B(n_272),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_550),
.A2(n_301),
.B1(n_322),
.B2(n_324),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_521),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_476),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_508),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_550),
.A2(n_520),
.B1(n_524),
.B2(n_523),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_473),
.B(n_322),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_509),
.B(n_322),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_518),
.B(n_324),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_530),
.A2(n_536),
.B(n_512),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_498),
.Y(n_599)
);

A2O1A1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_511),
.A2(n_192),
.B(n_251),
.C(n_257),
.Y(n_600)
);

A2O1A1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_489),
.A2(n_314),
.B(n_341),
.C(n_348),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_527),
.B(n_450),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_496),
.A2(n_314),
.B1(n_341),
.B2(n_348),
.Y(n_603)
);

NOR2xp67_ASAP7_75t_L g604 ( 
.A(n_506),
.B(n_8),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_507),
.B(n_314),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_505),
.B(n_341),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_497),
.B(n_389),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_528),
.A2(n_348),
.B1(n_359),
.B2(n_389),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_547),
.A2(n_390),
.B(n_385),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_505),
.B(n_359),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_531),
.B(n_495),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_519),
.A2(n_359),
.B(n_463),
.C(n_455),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_514),
.A2(n_435),
.B1(n_463),
.B2(n_455),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_505),
.B(n_8),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_522),
.B(n_404),
.Y(n_615)
);

BUFx8_ASAP7_75t_L g616 ( 
.A(n_548),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_506),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_515),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_515),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_516),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_532),
.Y(n_621)
);

AO22x1_ASAP7_75t_L g622 ( 
.A1(n_519),
.A2(n_404),
.B1(n_10),
.B2(n_11),
.Y(n_622)
);

CKINVDCx8_ASAP7_75t_R g623 ( 
.A(n_513),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_532),
.B(n_9),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_549),
.B(n_10),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_504),
.B(n_11),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_474),
.B(n_12),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_526),
.B(n_12),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_529),
.A2(n_407),
.B(n_448),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_482),
.B(n_391),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_533),
.B(n_542),
.Y(n_631)
);

CKINVDCx16_ASAP7_75t_R g632 ( 
.A(n_570),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_552),
.B(n_539),
.Y(n_633)
);

BUFx10_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_599),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_583),
.B(n_541),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_555),
.A2(n_545),
.B(n_525),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_557),
.A2(n_510),
.B(n_546),
.Y(n_638)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_591),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_611),
.B(n_482),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_561),
.A2(n_491),
.B(n_486),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_598),
.A2(n_485),
.B(n_484),
.Y(n_642)
);

AO31x2_ASAP7_75t_L g643 ( 
.A1(n_612),
.A2(n_422),
.A3(n_439),
.B(n_437),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_594),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_625),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_552),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_625),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_582),
.B(n_482),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_616),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_563),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_627),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_572),
.A2(n_433),
.B(n_432),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_569),
.B(n_482),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_617),
.B(n_14),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_573),
.A2(n_574),
.B(n_630),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_609),
.A2(n_413),
.B(n_410),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_554),
.B(n_15),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_621),
.Y(n_658)
);

NOR2xp67_ASAP7_75t_SL g659 ( 
.A(n_582),
.B(n_588),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_604),
.A2(n_391),
.B(n_17),
.C(n_18),
.Y(n_660)
);

A2O1A1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_628),
.A2(n_391),
.B(n_17),
.C(n_18),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_556),
.A2(n_391),
.B(n_19),
.C(n_20),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_558),
.A2(n_565),
.B(n_596),
.Y(n_663)
);

AO31x2_ASAP7_75t_L g664 ( 
.A1(n_600),
.A2(n_15),
.A3(n_21),
.B(n_22),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_582),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_631),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_559),
.B(n_23),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_629),
.A2(n_88),
.B(n_170),
.Y(n_668)
);

AOI21xp33_ASAP7_75t_L g669 ( 
.A1(n_568),
.A2(n_24),
.B(n_26),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_616),
.Y(n_670)
);

AO31x2_ASAP7_75t_L g671 ( 
.A1(n_586),
.A2(n_624),
.A3(n_595),
.B(n_597),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_603),
.B(n_589),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_588),
.Y(n_673)
);

AO22x2_ASAP7_75t_L g674 ( 
.A1(n_614),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_566),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_675)
);

NAND2x1_ASAP7_75t_L g676 ( 
.A(n_567),
.B(n_45),
.Y(n_676)
);

AO31x2_ASAP7_75t_L g677 ( 
.A1(n_590),
.A2(n_30),
.A3(n_34),
.B(n_35),
.Y(n_677)
);

NAND2x1p5_ASAP7_75t_L g678 ( 
.A(n_551),
.B(n_34),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_553),
.B(n_36),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_551),
.B(n_37),
.Y(n_680)
);

INVx3_ASAP7_75t_SL g681 ( 
.A(n_581),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_588),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_576),
.B(n_37),
.Y(n_683)
);

AND3x2_ASAP7_75t_L g684 ( 
.A(n_615),
.B(n_38),
.C(n_39),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_607),
.B(n_38),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_L g686 ( 
.A1(n_585),
.A2(n_92),
.B(n_157),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_618),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_618),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_560),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_577),
.B(n_39),
.Y(n_690)
);

AO31x2_ASAP7_75t_L g691 ( 
.A1(n_601),
.A2(n_40),
.A3(n_41),
.B(n_42),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_592),
.B(n_41),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_623),
.B(n_47),
.Y(n_693)
);

BUFx8_ASAP7_75t_L g694 ( 
.A(n_620),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_606),
.Y(n_695)
);

O2A1O1Ixp5_ASAP7_75t_L g696 ( 
.A1(n_610),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_622),
.B(n_79),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_593),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_602),
.B(n_90),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_605),
.A2(n_93),
.B(n_94),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_571),
.B(n_95),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_608),
.B(n_96),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_619),
.B(n_102),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_L g704 ( 
.A(n_626),
.B(n_104),
.C(n_110),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_613),
.A2(n_112),
.B(n_113),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_618),
.B(n_114),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_580),
.B(n_133),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_587),
.B(n_134),
.Y(n_708)
);

AND2x6_ASAP7_75t_L g709 ( 
.A(n_584),
.B(n_137),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_575),
.A2(n_140),
.B(n_144),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_579),
.B(n_147),
.Y(n_711)
);

OAI22x1_ASAP7_75t_L g712 ( 
.A1(n_567),
.A2(n_176),
.B1(n_155),
.B2(n_156),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_567),
.Y(n_713)
);

AO31x2_ASAP7_75t_L g714 ( 
.A1(n_562),
.A2(n_612),
.A3(n_564),
.B(n_578),
.Y(n_714)
);

OAI22x1_ASAP7_75t_L g715 ( 
.A1(n_625),
.A2(n_361),
.B1(n_540),
.B2(n_336),
.Y(n_715)
);

AO31x2_ASAP7_75t_L g716 ( 
.A1(n_562),
.A2(n_612),
.A3(n_564),
.B(n_578),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_563),
.A2(n_578),
.B1(n_565),
.B2(n_558),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_611),
.B(n_480),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_718),
.A2(n_685),
.B(n_672),
.C(n_662),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_634),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_635),
.B(n_666),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_679),
.A2(n_697),
.B1(n_715),
.B2(n_667),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_666),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_658),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_670),
.B(n_649),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_632),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_639),
.B(n_647),
.Y(n_727)
);

AOI222xp33_ASAP7_75t_L g728 ( 
.A1(n_636),
.A2(n_644),
.B1(n_645),
.B2(n_695),
.C1(n_692),
.C2(n_674),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_697),
.A2(n_650),
.B1(n_717),
.B2(n_702),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_640),
.A2(n_674),
.B1(n_678),
.B2(n_657),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_689),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_634),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_646),
.B(n_665),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_665),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_660),
.B(n_661),
.C(n_669),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_689),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_663),
.A2(n_654),
.B(n_653),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_698),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_675),
.A2(n_651),
.B1(n_690),
.B2(n_683),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_682),
.B(n_673),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_L g741 ( 
.A1(n_638),
.A2(n_637),
.B(n_642),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_SL g742 ( 
.A1(n_676),
.A2(n_686),
.B(n_706),
.C(n_648),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_680),
.A2(n_713),
.B1(n_703),
.B2(n_687),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_696),
.A2(n_641),
.B(n_668),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_694),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_673),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_705),
.A2(n_704),
.B(n_710),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_694),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_643),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_677),
.Y(n_750)
);

CKINVDCx16_ASAP7_75t_R g751 ( 
.A(n_709),
.Y(n_751)
);

AOI22x1_ASAP7_75t_L g752 ( 
.A1(n_712),
.A2(n_700),
.B1(n_699),
.B2(n_711),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_707),
.A2(n_708),
.B(n_701),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_633),
.B(n_681),
.Y(n_754)
);

AOI31xp67_ASAP7_75t_L g755 ( 
.A1(n_714),
.A2(n_716),
.A3(n_643),
.B(n_671),
.Y(n_755)
);

CKINVDCx6p67_ASAP7_75t_R g756 ( 
.A(n_709),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_688),
.Y(n_757)
);

CKINVDCx6p67_ASAP7_75t_R g758 ( 
.A(n_709),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_713),
.B(n_693),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_671),
.B(n_716),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_671),
.B(n_664),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_664),
.B(n_684),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_691),
.A2(n_677),
.B(n_664),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_691),
.A2(n_578),
.B(n_655),
.Y(n_764)
);

OAI21x1_ASAP7_75t_L g765 ( 
.A1(n_691),
.A2(n_652),
.B(n_656),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_718),
.B(n_497),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_639),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_635),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_639),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_639),
.Y(n_770)
);

BUFx8_ASAP7_75t_L g771 ( 
.A(n_670),
.Y(n_771)
);

O2A1O1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_718),
.A2(n_506),
.B(n_495),
.C(n_519),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_635),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_639),
.B(n_480),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_639),
.B(n_480),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_718),
.A2(n_563),
.B1(n_611),
.B2(n_685),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_644),
.A2(n_563),
.B1(n_697),
.B2(n_650),
.Y(n_777)
);

NAND2x1p5_ASAP7_75t_L g778 ( 
.A(n_659),
.B(n_552),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_694),
.Y(n_779)
);

CKINVDCx9p33_ASAP7_75t_R g780 ( 
.A(n_670),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_644),
.A2(n_604),
.B(n_650),
.C(n_563),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_639),
.B(n_480),
.Y(n_782)
);

BUFx2_ASAP7_75t_R g783 ( 
.A(n_649),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_639),
.B(n_480),
.Y(n_784)
);

OA21x2_ASAP7_75t_L g785 ( 
.A1(n_655),
.A2(n_652),
.B(n_656),
.Y(n_785)
);

AO32x2_ASAP7_75t_L g786 ( 
.A1(n_675),
.A2(n_506),
.A3(n_519),
.B1(n_586),
.B2(n_717),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_685),
.A2(n_396),
.B1(n_399),
.B2(n_535),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_L g788 ( 
.A(n_715),
.B(n_540),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_666),
.B(n_552),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_644),
.B(n_666),
.Y(n_790)
);

AOI21xp33_ASAP7_75t_SL g791 ( 
.A1(n_632),
.A2(n_681),
.B(n_476),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_718),
.B(n_611),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_650),
.A2(n_564),
.B(n_578),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_718),
.B(n_497),
.Y(n_794)
);

OA21x2_ASAP7_75t_L g795 ( 
.A1(n_763),
.A2(n_764),
.B(n_765),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_738),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_768),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_767),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_773),
.Y(n_799)
);

CKINVDCx6p67_ASAP7_75t_R g800 ( 
.A(n_780),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_724),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_769),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_731),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_736),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_723),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_779),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_766),
.B(n_794),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_735),
.A2(n_776),
.B(n_719),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_751),
.Y(n_809)
);

CKINVDCx12_ASAP7_75t_R g810 ( 
.A(n_725),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_790),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_785),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_777),
.A2(n_728),
.B1(n_722),
.B2(n_792),
.Y(n_813)
);

AND2x4_ASAP7_75t_SL g814 ( 
.A(n_748),
.B(n_756),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_750),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_758),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_761),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_789),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_755),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_749),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_726),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_721),
.B(n_774),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_770),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_770),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_777),
.A2(n_728),
.B1(n_730),
.B2(n_776),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_775),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_782),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_784),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_733),
.Y(n_829)
);

AO21x2_ASAP7_75t_L g830 ( 
.A1(n_761),
.A2(n_741),
.B(n_760),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_734),
.B(n_739),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_734),
.B(n_739),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_771),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_762),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_730),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_727),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_720),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_786),
.B(n_757),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_786),
.B(n_781),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_793),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_729),
.A2(n_787),
.B1(n_788),
.B2(n_743),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_732),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_793),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_740),
.Y(n_844)
);

BUFx2_ASAP7_75t_L g845 ( 
.A(n_743),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_740),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_791),
.B(n_745),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_778),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_778),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_772),
.B(n_754),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_786),
.B(n_746),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_725),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_725),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_735),
.A2(n_771),
.B1(n_737),
.B2(n_759),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_797),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_822),
.B(n_759),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_799),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_803),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_835),
.B(n_825),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_823),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_804),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_827),
.B(n_752),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_815),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_826),
.B(n_753),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_800),
.A2(n_783),
.B1(n_744),
.B2(n_747),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_828),
.B(n_742),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_813),
.B(n_744),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_806),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_834),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_836),
.B(n_801),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_801),
.B(n_829),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_845),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_838),
.B(n_796),
.Y(n_873)
);

BUFx8_ASAP7_75t_L g874 ( 
.A(n_809),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_824),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_820),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_831),
.B(n_832),
.Y(n_877)
);

NAND2x1p5_ASAP7_75t_L g878 ( 
.A(n_816),
.B(n_818),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_817),
.B(n_805),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_800),
.A2(n_809),
.B1(n_814),
.B2(n_854),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_817),
.B(n_811),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_811),
.B(n_851),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_807),
.B(n_798),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_851),
.B(n_839),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_839),
.B(n_808),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_802),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_831),
.B(n_832),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_819),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_819),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_810),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_884),
.B(n_843),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_884),
.B(n_843),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_885),
.B(n_840),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_873),
.B(n_830),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_865),
.B(n_880),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_869),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_863),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_885),
.B(n_830),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_888),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_882),
.B(n_812),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_876),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_881),
.B(n_841),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_868),
.B(n_816),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_868),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_877),
.B(n_795),
.Y(n_905)
);

NOR2x1_ASAP7_75t_L g906 ( 
.A(n_866),
.B(n_816),
.Y(n_906)
);

NOR2x1p5_ASAP7_75t_L g907 ( 
.A(n_867),
.B(n_833),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_877),
.B(n_887),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_859),
.B(n_850),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_887),
.B(n_795),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_901),
.Y(n_911)
);

AND2x4_ASAP7_75t_SL g912 ( 
.A(n_900),
.B(n_879),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_891),
.B(n_886),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_905),
.B(n_887),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_905),
.B(n_889),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_901),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_904),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_891),
.B(n_860),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_899),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_898),
.B(n_893),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_892),
.B(n_875),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_898),
.B(n_872),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_897),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_892),
.B(n_859),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_897),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_910),
.B(n_894),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_909),
.B(n_855),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_912),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_920),
.B(n_894),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_923),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_917),
.B(n_895),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_911),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_923),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_925),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_919),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_918),
.A2(n_895),
.B1(n_909),
.B2(n_907),
.Y(n_936)
);

NOR2x1p5_ASAP7_75t_SL g937 ( 
.A(n_922),
.B(n_899),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_912),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_912),
.A2(n_908),
.B(n_883),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_936),
.A2(n_907),
.B1(n_924),
.B2(n_908),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_930),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_928),
.A2(n_917),
.B1(n_921),
.B2(n_904),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_931),
.A2(n_906),
.B(n_896),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_932),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_935),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_938),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_933),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_939),
.A2(n_902),
.B1(n_906),
.B2(n_915),
.Y(n_948)
);

AOI32xp33_ASAP7_75t_L g949 ( 
.A1(n_928),
.A2(n_914),
.A3(n_926),
.B1(n_904),
.B2(n_814),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_934),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_935),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_946),
.A2(n_938),
.B1(n_928),
.B2(n_931),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_946),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_944),
.B(n_926),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_948),
.B(n_920),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_953),
.B(n_833),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_954),
.Y(n_957)
);

OAI21xp33_ASAP7_75t_L g958 ( 
.A1(n_952),
.A2(n_940),
.B(n_949),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_957),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_956),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_959),
.B(n_958),
.Y(n_961)
);

NAND4xp75_ASAP7_75t_L g962 ( 
.A(n_960),
.B(n_847),
.C(n_943),
.D(n_955),
.Y(n_962)
);

NOR3xp33_ASAP7_75t_L g963 ( 
.A(n_961),
.B(n_962),
.C(n_960),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_L g964 ( 
.A1(n_961),
.A2(n_806),
.B(n_942),
.Y(n_964)
);

NAND4xp75_ASAP7_75t_L g965 ( 
.A(n_963),
.B(n_821),
.C(n_903),
.D(n_937),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_964),
.A2(n_890),
.B(n_852),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_966),
.A2(n_878),
.B1(n_853),
.B2(n_864),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_965),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_966),
.Y(n_969)
);

NOR2x1_ASAP7_75t_L g970 ( 
.A(n_968),
.B(n_821),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_969),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_967),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_968),
.Y(n_973)
);

OAI211xp5_ASAP7_75t_L g974 ( 
.A1(n_968),
.A2(n_821),
.B(n_842),
.C(n_837),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_970),
.Y(n_975)
);

OAI22xp33_ASAP7_75t_L g976 ( 
.A1(n_973),
.A2(n_878),
.B1(n_927),
.B2(n_947),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_972),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_971),
.Y(n_978)
);

OAI22xp33_ASAP7_75t_L g979 ( 
.A1(n_974),
.A2(n_878),
.B1(n_950),
.B2(n_941),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_973),
.A2(n_913),
.B1(n_862),
.B2(n_945),
.Y(n_980)
);

NAND2x1_ASAP7_75t_SL g981 ( 
.A(n_970),
.B(n_810),
.Y(n_981)
);

AOI221x1_ASAP7_75t_L g982 ( 
.A1(n_978),
.A2(n_951),
.B1(n_857),
.B2(n_870),
.C(n_861),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_975),
.A2(n_916),
.B(n_951),
.Y(n_983)
);

XNOR2xp5_ASAP7_75t_L g984 ( 
.A(n_977),
.B(n_874),
.Y(n_984)
);

OAI22xp33_ASAP7_75t_L g985 ( 
.A1(n_980),
.A2(n_945),
.B1(n_929),
.B2(n_896),
.Y(n_985)
);

AOI22x1_ASAP7_75t_L g986 ( 
.A1(n_984),
.A2(n_981),
.B1(n_976),
.B2(n_979),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_983),
.A2(n_848),
.B(n_849),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_985),
.A2(n_874),
.B1(n_846),
.B2(n_844),
.Y(n_988)
);

OA21x2_ASAP7_75t_L g989 ( 
.A1(n_986),
.A2(n_982),
.B(n_858),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_988),
.A2(n_871),
.B(n_856),
.Y(n_990)
);

XOR2xp5_ASAP7_75t_L g991 ( 
.A(n_989),
.B(n_987),
.Y(n_991)
);

AOI21xp33_ASAP7_75t_L g992 ( 
.A1(n_991),
.A2(n_990),
.B(n_874),
.Y(n_992)
);


endmodule